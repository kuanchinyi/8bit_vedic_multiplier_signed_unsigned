// This is the unpowered netlist.
module vmsu_8bit_top (clk,
    control,
    rst,
    a,
    b,
    p);
 input clk;
 input control;
 input rst;
 input [7:0] a;
 input [7:0] b;
 output [15:0] p;

 wire \FA0.q ;
 wire \FA1.q ;
 wire \FA2.q ;
 wire \FA3.q ;
 wire \FA4.q ;
 wire \FA5.q ;
 wire \FA6.q ;
 wire \FA7.q ;
 wire \FB0.q ;
 wire \FB1.q ;
 wire \FB2.q ;
 wire \FB3.q ;
 wire \FB4.q ;
 wire \FB5.q ;
 wire \FB6.q ;
 wire \FB7.q ;
 wire \FC.q ;
 wire \FP0.d ;
 wire \FP1.d ;
 wire \FP10.d ;
 wire \FP11.d ;
 wire \FP12.d ;
 wire \FP13.d ;
 wire \FP14.d ;
 wire \FP15.d ;
 wire \FP2.d ;
 wire \FP3.d ;
 wire \FP4.d ;
 wire \FP5.d ;
 wire \FP6.d ;
 wire \FP7.d ;
 wire \FP8.d ;
 wire \FP9.d ;
 wire \M0.FAM0.d ;
 wire \M0.FAM0.q ;
 wire \M0.FAM1.d ;
 wire \M0.FAM1.q ;
 wire \M0.FAM2.d ;
 wire \M0.FAM2.q ;
 wire \M0.FAM3.d ;
 wire \M0.FAM3.q ;
 wire \M0.FAM4.d ;
 wire \M0.FAM4.q ;
 wire \M0.FAM5.d ;
 wire \M0.FAM5.q ;
 wire \M0.FAM6.d ;
 wire \M0.FAM6.q ;
 wire \M0.FAM7.d ;
 wire \M0.FAM7.q ;
 wire \M0.FBM0.d ;
 wire \M0.FBM0.q ;
 wire \M0.FBM1.d ;
 wire \M0.FBM1.q ;
 wire \M0.FBM2.d ;
 wire \M0.FBM2.q ;
 wire \M0.FBM3.d ;
 wire \M0.FBM3.q ;
 wire \M0.FBM4.d ;
 wire \M0.FBM4.q ;
 wire \M0.FBM5.d ;
 wire \M0.FBM5.q ;
 wire \M0.FBM6.d ;
 wire \M0.FBM6.q ;
 wire \M0.FBM7.d ;
 wire \M0.FBM7.q ;
 wire \M0.FPM0.d ;
 wire \M0.FPM0.q ;
 wire \M0.FPM1.d ;
 wire \M0.FPM1.q ;
 wire \M0.FPM10.d ;
 wire \M0.FPM10.q ;
 wire \M0.FPM11.d ;
 wire \M0.FPM11.q ;
 wire \M0.FPM12.d ;
 wire \M0.FPM12.q ;
 wire \M0.FPM13.d ;
 wire \M0.FPM13.q ;
 wire \M0.FPM14.d ;
 wire \M0.FPM14.q ;
 wire \M0.FPM15.d ;
 wire \M0.FPM15.q ;
 wire \M0.FPM2.d ;
 wire \M0.FPM2.q ;
 wire \M0.FPM3.d ;
 wire \M0.FPM3.q ;
 wire \M0.FPM4.d ;
 wire \M0.FPM4.q ;
 wire \M0.FPM5.d ;
 wire \M0.FPM5.q ;
 wire \M0.FPM6.d ;
 wire \M0.FPM6.q ;
 wire \M0.FPM7.d ;
 wire \M0.FPM7.q ;
 wire \M0.FPM8.d ;
 wire \M0.FPM8.q ;
 wire \M0.FPM9.d ;
 wire \M0.FPM9.q ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__0545__B1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0548__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0550__B1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0552__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0554__C1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0556__B1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0558__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0564__B1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0567__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0569__B1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0571__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0573__C1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0575__B1 (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0577__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0589__A (.DIODE(\FC.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0590__A (.DIODE(_0095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0591__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0593__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0595__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0597__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0599__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0601__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0603__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0605__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0607__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0609__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0611__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0613__A (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0615__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0617__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0619__B (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0626__B (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__C (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0631__D (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__B (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__C (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0632__D (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__C (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0633__D (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0635__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0636__B (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0638__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0639__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0641__B (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0642__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0646__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0647__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0648__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0649__B (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0653__B2 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__B1 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0661__C1 (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0685__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0687__B (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__A1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0688__A2 (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0689__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__A (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0690__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__B (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__B (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__C (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0696__D (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__C (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0697__D (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0699__B (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0704__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0705__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0708__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0710__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__A1 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__A2 (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__B1 (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0711__B2 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__C (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0712__D (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__C (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__D (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0722__B (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0723__A1 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__A (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__A (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0748__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__B1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__C1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__B1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0754__C1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__A1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__B1 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0758__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0759__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0760__A1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0760__B1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0761__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0762__C_N (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0763__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0764__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0768__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0769__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0770__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0771__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A2 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__C (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__D (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__A1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__A2 (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0785__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__A (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0790__B (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0793__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0794__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0797__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0798__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__A_N (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0799__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0800__B1 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0801__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0802__A1 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0804__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__A (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0805__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__A_N (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0807__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__A1 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__A2 (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0808__B1_N (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__A_N (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__B (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0809__C (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__A1 (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__C1 (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0841__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0842__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0843__B1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0845__A1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0846__A (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__C (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0847__D (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__C (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__D (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__C (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0858__D (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0861__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0862__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__C1 (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__D1 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A1 (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A2 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__C (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0866__D (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0867__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0870__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0874__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0875__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0876__A (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__A1 (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__A3 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0879__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0882__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0886__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0887__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0895__A1 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__B (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__C (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0902__D (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0903__A1 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0908__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0926__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0954__B (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A2 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A3 (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0955__A4 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__A (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0956__B (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__B1 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0964__C1 (.DIODE(_0247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0984__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0985__B (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0986__B2 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0987__A (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__A1_N (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0988__A2_N (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0990__A1 (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0991__B (.DIODE(_0120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0992__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A1 (.DIODE(_0113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1010__A2 (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__A (.DIODE(_0176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1048__B (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__A (.DIODE(_0174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1049__B (.DIODE(_0236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__A (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1052__C (.DIODE(_0237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1053__A1 (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1055__A1 (.DIODE(_0234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1066__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1067__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1068__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1069__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1070__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1071__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1072__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1073__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1074__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1075__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1076__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1077__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1078__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1079__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1080__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1081__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1082__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1083__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1084__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1085__A (.DIODE(_0540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1086__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1087__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1088__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1089__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1090__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1091__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1092__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1093__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1094__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1095__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1096__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1097__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1098__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1099__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1100__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1101__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1102__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1103__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1104__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1105__A (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1106__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1110__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1112__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1115__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1116__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1118__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1123__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1124__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1125__A (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1126__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1127__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1128__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1129__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1130__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1131__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1132__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1133__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__CLK (.DIODE(net17));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__or4_1 _0543_ (.A(\FB0.q ),
    .B(\FB1.q ),
    .C(\FB2.q ),
    .D(\FB3.q ),
    .X(_0065_));
 sky130_fd_sc_hd__or3_1 _0544_ (.A(\FB4.q ),
    .B(\FB5.q ),
    .C(_0065_),
    .X(_0066_));
 sky130_fd_sc_hd__o21ai_1 _0545_ (.A1(\FB6.q ),
    .A2(_0066_),
    .B1(\FC.q ),
    .Y(_0067_));
 sky130_fd_sc_hd__and2_1 _0546_ (.A(\FB7.q ),
    .B(_0067_),
    .X(_0068_));
 sky130_fd_sc_hd__clkbuf_1 _0547_ (.A(_0068_),
    .X(\M0.FBM7.d ));
 sky130_fd_sc_hd__and3_1 _0548_ (.A(\FC.q ),
    .B(\FB7.q ),
    .C(_0066_),
    .X(_0069_));
 sky130_fd_sc_hd__xor2_1 _0549_ (.A(\FB6.q ),
    .B(_0069_),
    .X(\M0.FBM6.d ));
 sky130_fd_sc_hd__o211a_1 _0550_ (.A1(\FB4.q ),
    .A2(_0065_),
    .B1(\FC.q ),
    .C1(\FB7.q ),
    .X(_0070_));
 sky130_fd_sc_hd__xor2_1 _0551_ (.A(\FB5.q ),
    .B(_0070_),
    .X(\M0.FBM5.d ));
 sky130_fd_sc_hd__and3_1 _0552_ (.A(\FC.q ),
    .B(\FB7.q ),
    .C(_0065_),
    .X(_0071_));
 sky130_fd_sc_hd__xor2_1 _0553_ (.A(\FB4.q ),
    .B(_0071_),
    .X(\M0.FBM4.d ));
 sky130_fd_sc_hd__o311a_1 _0554_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .A3(\FB2.q ),
    .B1(\FB7.q ),
    .C1(\FC.q ),
    .X(_0072_));
 sky130_fd_sc_hd__xor2_1 _0555_ (.A(\FB3.q ),
    .B(_0072_),
    .X(\M0.FBM3.d ));
 sky130_fd_sc_hd__o211a_1 _0556_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .B1(\FC.q ),
    .C1(\FB7.q ),
    .X(_0073_));
 sky130_fd_sc_hd__xor2_1 _0557_ (.A(\FB2.q ),
    .B(_0073_),
    .X(\M0.FBM2.d ));
 sky130_fd_sc_hd__and3_1 _0558_ (.A(\FC.q ),
    .B(\FB7.q ),
    .C(\FB0.q ),
    .X(_0074_));
 sky130_fd_sc_hd__xor2_1 _0559_ (.A(\FB1.q ),
    .B(_0074_),
    .X(\M0.FBM1.d ));
 sky130_fd_sc_hd__clkbuf_1 _0560_ (.A(\FB0.q ),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_1 _0561_ (.A(_0075_),
    .X(\M0.FBM0.d ));
 sky130_fd_sc_hd__or4_2 _0562_ (.A(\FA0.q ),
    .B(\FA1.q ),
    .C(\FA2.q ),
    .D(\FA3.q ),
    .X(_0076_));
 sky130_fd_sc_hd__or3_1 _0563_ (.A(\FA4.q ),
    .B(\FA5.q ),
    .C(_0076_),
    .X(_0077_));
 sky130_fd_sc_hd__o21ai_1 _0564_ (.A1(\FA6.q ),
    .A2(_0077_),
    .B1(\FC.q ),
    .Y(_0078_));
 sky130_fd_sc_hd__and2_1 _0565_ (.A(\FA7.q ),
    .B(_0078_),
    .X(_0079_));
 sky130_fd_sc_hd__clkbuf_1 _0566_ (.A(_0079_),
    .X(\M0.FAM7.d ));
 sky130_fd_sc_hd__and3_1 _0567_ (.A(\FC.q ),
    .B(\FA7.q ),
    .C(_0077_),
    .X(_0080_));
 sky130_fd_sc_hd__xor2_1 _0568_ (.A(\FA6.q ),
    .B(_0080_),
    .X(\M0.FAM6.d ));
 sky130_fd_sc_hd__o211a_1 _0569_ (.A1(\FA4.q ),
    .A2(_0076_),
    .B1(\FC.q ),
    .C1(\FA7.q ),
    .X(_0081_));
 sky130_fd_sc_hd__xor2_1 _0570_ (.A(\FA5.q ),
    .B(_0081_),
    .X(\M0.FAM5.d ));
 sky130_fd_sc_hd__and3_1 _0571_ (.A(\FC.q ),
    .B(\FA7.q ),
    .C(_0076_),
    .X(_0082_));
 sky130_fd_sc_hd__xor2_1 _0572_ (.A(\FA4.q ),
    .B(_0082_),
    .X(\M0.FAM4.d ));
 sky130_fd_sc_hd__o311a_1 _0573_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .A3(\FA2.q ),
    .B1(\FA7.q ),
    .C1(\FC.q ),
    .X(_0083_));
 sky130_fd_sc_hd__xor2_1 _0574_ (.A(\FA3.q ),
    .B(_0083_),
    .X(\M0.FAM3.d ));
 sky130_fd_sc_hd__o211a_1 _0575_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .B1(\FC.q ),
    .C1(\FA7.q ),
    .X(_0084_));
 sky130_fd_sc_hd__xor2_1 _0576_ (.A(\FA2.q ),
    .B(_0084_),
    .X(\M0.FAM2.d ));
 sky130_fd_sc_hd__and3_1 _0577_ (.A(\FC.q ),
    .B(\FA7.q ),
    .C(\FA0.q ),
    .X(_0085_));
 sky130_fd_sc_hd__xor2_1 _0578_ (.A(\FA1.q ),
    .B(_0085_),
    .X(\M0.FAM1.d ));
 sky130_fd_sc_hd__clkbuf_1 _0579_ (.A(\FA0.q ),
    .X(_0086_));
 sky130_fd_sc_hd__clkbuf_1 _0580_ (.A(_0086_),
    .X(\M0.FAM0.d ));
 sky130_fd_sc_hd__or4_1 _0581_ (.A(\M0.FPM0.q ),
    .B(\M0.FPM1.q ),
    .C(\M0.FPM2.q ),
    .D(\M0.FPM3.q ),
    .X(_0087_));
 sky130_fd_sc_hd__or3_1 _0582_ (.A(\M0.FPM4.q ),
    .B(\M0.FPM5.q ),
    .C(_0087_),
    .X(_0088_));
 sky130_fd_sc_hd__or2_1 _0583_ (.A(\M0.FPM6.q ),
    .B(_0088_),
    .X(_0089_));
 sky130_fd_sc_hd__or3_1 _0584_ (.A(\M0.FPM7.q ),
    .B(\M0.FPM8.q ),
    .C(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__or2_1 _0585_ (.A(\M0.FPM9.q ),
    .B(_0090_),
    .X(_0091_));
 sky130_fd_sc_hd__or3_1 _0586_ (.A(\M0.FPM10.q ),
    .B(\M0.FPM11.q ),
    .C(_0091_),
    .X(_0092_));
 sky130_fd_sc_hd__or2_1 _0587_ (.A(\M0.FPM12.q ),
    .B(_0092_),
    .X(_0093_));
 sky130_fd_sc_hd__xor2_1 _0588_ (.A(\FB7.q ),
    .B(\FA7.q ),
    .X(_0094_));
 sky130_fd_sc_hd__and2_1 _0589_ (.A(\FC.q ),
    .B(_0094_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_4 _0590_ (.A(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__o31a_1 _0591_ (.A1(\M0.FPM14.q ),
    .A2(\M0.FPM13.q ),
    .A3(_0093_),
    .B1(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__xor2_1 _0592_ (.A(\M0.FPM15.q ),
    .B(_0097_),
    .X(\FP15.d ));
 sky130_fd_sc_hd__o21ai_1 _0593_ (.A1(\M0.FPM13.q ),
    .A2(_0093_),
    .B1(_0096_),
    .Y(_0098_));
 sky130_fd_sc_hd__xnor2_1 _0594_ (.A(\M0.FPM14.q ),
    .B(_0098_),
    .Y(\FP14.d ));
 sky130_fd_sc_hd__nand2_1 _0595_ (.A(_0096_),
    .B(_0093_),
    .Y(_0099_));
 sky130_fd_sc_hd__xnor2_1 _0596_ (.A(\M0.FPM13.q ),
    .B(_0099_),
    .Y(\FP13.d ));
 sky130_fd_sc_hd__nand2_1 _0597_ (.A(_0096_),
    .B(_0092_),
    .Y(_0100_));
 sky130_fd_sc_hd__xnor2_1 _0598_ (.A(\M0.FPM12.q ),
    .B(_0100_),
    .Y(\FP12.d ));
 sky130_fd_sc_hd__o21ai_1 _0599_ (.A1(\M0.FPM10.q ),
    .A2(_0091_),
    .B1(_0096_),
    .Y(_0101_));
 sky130_fd_sc_hd__xnor2_1 _0600_ (.A(\M0.FPM11.q ),
    .B(_0101_),
    .Y(\FP11.d ));
 sky130_fd_sc_hd__nand2_1 _0601_ (.A(_0096_),
    .B(_0091_),
    .Y(_0102_));
 sky130_fd_sc_hd__xnor2_1 _0602_ (.A(\M0.FPM10.q ),
    .B(_0102_),
    .Y(\FP10.d ));
 sky130_fd_sc_hd__nand2_1 _0603_ (.A(_0096_),
    .B(_0090_),
    .Y(_0103_));
 sky130_fd_sc_hd__xnor2_1 _0604_ (.A(\M0.FPM9.q ),
    .B(_0103_),
    .Y(\FP9.d ));
 sky130_fd_sc_hd__o21ai_1 _0605_ (.A1(\M0.FPM7.q ),
    .A2(_0089_),
    .B1(_0096_),
    .Y(_0104_));
 sky130_fd_sc_hd__xnor2_1 _0606_ (.A(\M0.FPM8.q ),
    .B(_0104_),
    .Y(\FP8.d ));
 sky130_fd_sc_hd__nand2_1 _0607_ (.A(_0096_),
    .B(_0089_),
    .Y(_0105_));
 sky130_fd_sc_hd__xnor2_1 _0608_ (.A(\M0.FPM7.q ),
    .B(_0105_),
    .Y(\FP7.d ));
 sky130_fd_sc_hd__nand2_1 _0609_ (.A(_0096_),
    .B(_0088_),
    .Y(_0106_));
 sky130_fd_sc_hd__xnor2_1 _0610_ (.A(\M0.FPM6.q ),
    .B(_0106_),
    .Y(\FP6.d ));
 sky130_fd_sc_hd__o21ai_1 _0611_ (.A1(\M0.FPM4.q ),
    .A2(_0087_),
    .B1(_0096_),
    .Y(_0107_));
 sky130_fd_sc_hd__xnor2_1 _0612_ (.A(\M0.FPM5.q ),
    .B(_0107_),
    .Y(\FP5.d ));
 sky130_fd_sc_hd__nand2_1 _0613_ (.A(_0096_),
    .B(_0087_),
    .Y(_0108_));
 sky130_fd_sc_hd__xnor2_1 _0614_ (.A(\M0.FPM4.q ),
    .B(_0108_),
    .Y(\FP4.d ));
 sky130_fd_sc_hd__o31a_1 _0615_ (.A1(\M0.FPM0.q ),
    .A2(\M0.FPM1.q ),
    .A3(\M0.FPM2.q ),
    .B1(_0096_),
    .X(_0109_));
 sky130_fd_sc_hd__xor2_1 _0616_ (.A(\M0.FPM3.q ),
    .B(_0109_),
    .X(\FP3.d ));
 sky130_fd_sc_hd__o21ai_1 _0617_ (.A1(\M0.FPM0.q ),
    .A2(\M0.FPM1.q ),
    .B1(_0096_),
    .Y(_0110_));
 sky130_fd_sc_hd__xnor2_1 _0618_ (.A(\M0.FPM2.q ),
    .B(_0110_),
    .Y(\FP2.d ));
 sky130_fd_sc_hd__nand2_1 _0619_ (.A(\M0.FPM0.q ),
    .B(_0096_),
    .Y(_0111_));
 sky130_fd_sc_hd__xnor2_1 _0620_ (.A(\M0.FPM1.q ),
    .B(_0111_),
    .Y(\FP1.d ));
 sky130_fd_sc_hd__clkbuf_1 _0621_ (.A(\M0.FPM0.q ),
    .X(_0112_));
 sky130_fd_sc_hd__clkbuf_1 _0622_ (.A(_0112_),
    .X(\FP0.d ));
 sky130_fd_sc_hd__buf_4 _0623_ (.A(\M0.FAM7.q ),
    .X(_0113_));
 sky130_fd_sc_hd__buf_6 _0624_ (.A(\M0.FAM6.q ),
    .X(_0114_));
 sky130_fd_sc_hd__buf_6 _0625_ (.A(\M0.FBM6.q ),
    .X(_0115_));
 sky130_fd_sc_hd__and2_1 _0626_ (.A(_0114_),
    .B(_0115_),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_8 _0627_ (.A(\M0.FAM5.q ),
    .X(_0117_));
 sky130_fd_sc_hd__buf_8 _0628_ (.A(\M0.FAM4.q ),
    .X(_0118_));
 sky130_fd_sc_hd__clkbuf_8 _0629_ (.A(\M0.FBM5.q ),
    .X(_0119_));
 sky130_fd_sc_hd__buf_8 _0630_ (.A(\M0.FBM4.q ),
    .X(_0120_));
 sky130_fd_sc_hd__and4_1 _0631_ (.A(_0117_),
    .B(_0118_),
    .C(_0119_),
    .D(_0120_),
    .X(_0121_));
 sky130_fd_sc_hd__and4_1 _0632_ (.A(\M0.FBM7.q ),
    .B(_0115_),
    .C(_0117_),
    .D(_0118_),
    .X(_0122_));
 sky130_fd_sc_hd__and4_1 _0633_ (.A(_0113_),
    .B(_0114_),
    .C(_0119_),
    .D(_0120_),
    .X(_0123_));
 sky130_fd_sc_hd__xnor2_1 _0634_ (.A(_0122_),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__nand2_1 _0635_ (.A(\M0.FBM7.q ),
    .B(_0118_),
    .Y(_0125_));
 sky130_fd_sc_hd__nand2_1 _0636_ (.A(_0115_),
    .B(_0117_),
    .Y(_0126_));
 sky130_fd_sc_hd__xor2_2 _0637_ (.A(_0125_),
    .B(_0126_),
    .X(_0127_));
 sky130_fd_sc_hd__nand2_1 _0638_ (.A(_0113_),
    .B(_0120_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _0639_ (.A(_0114_),
    .B(_0119_),
    .Y(_0129_));
 sky130_fd_sc_hd__xor2_2 _0640_ (.A(_0128_),
    .B(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__nand2_1 _0641_ (.A(_0114_),
    .B(_0115_),
    .Y(_0131_));
 sky130_fd_sc_hd__nand2_2 _0642_ (.A(_0118_),
    .B(_0120_),
    .Y(_0132_));
 sky130_fd_sc_hd__nor2_1 _0643_ (.A(_0131_),
    .B(_0132_),
    .Y(_0133_));
 sky130_fd_sc_hd__a21o_1 _0644_ (.A1(_0127_),
    .A2(_0130_),
    .B1(_0133_),
    .X(_0134_));
 sky130_fd_sc_hd__o21a_1 _0645_ (.A1(_0127_),
    .A2(_0130_),
    .B1(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__nand2_1 _0646_ (.A(_0114_),
    .B(_0120_),
    .Y(_0136_));
 sky130_fd_sc_hd__and3_1 _0647_ (.A(_0113_),
    .B(_0119_),
    .C(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__nand2_1 _0648_ (.A(_0115_),
    .B(_0118_),
    .Y(_0138_));
 sky130_fd_sc_hd__and3_1 _0649_ (.A(\M0.FBM7.q ),
    .B(_0117_),
    .C(_0138_),
    .X(_0139_));
 sky130_fd_sc_hd__xnor2_1 _0650_ (.A(_0137_),
    .B(_0139_),
    .Y(_0140_));
 sky130_fd_sc_hd__xnor2_1 _0651_ (.A(_0135_),
    .B(_0140_),
    .Y(_0141_));
 sky130_fd_sc_hd__nand2_1 _0652_ (.A(_0117_),
    .B(_0119_),
    .Y(_0142_));
 sky130_fd_sc_hd__o22a_1 _0653_ (.A1(_0118_),
    .A2(_0136_),
    .B1(_0138_),
    .B2(_0120_),
    .X(_0143_));
 sky130_fd_sc_hd__nor2_1 _0654_ (.A(_0142_),
    .B(_0143_),
    .Y(_0144_));
 sky130_fd_sc_hd__xnor2_1 _0655_ (.A(_0127_),
    .B(_0130_),
    .Y(_0145_));
 sky130_fd_sc_hd__xnor2_1 _0656_ (.A(_0133_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__o21a_1 _0657_ (.A1(_0121_),
    .A2(_0144_),
    .B1(_0146_),
    .X(_0147_));
 sky130_fd_sc_hd__nand2_1 _0658_ (.A(_0141_),
    .B(_0147_),
    .Y(_0148_));
 sky130_fd_sc_hd__nor2_1 _0659_ (.A(_0124_),
    .B(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__and2_1 _0660_ (.A(_0121_),
    .B(_0149_),
    .X(_0150_));
 sky130_fd_sc_hd__o211ai_1 _0661_ (.A1(_0121_),
    .A2(_0131_),
    .B1(_0113_),
    .C1(\M0.FBM7.q ),
    .Y(_0151_));
 sky130_fd_sc_hd__o2bb2a_1 _0662_ (.A1_N(_0144_),
    .A2_N(_0149_),
    .B1(_0150_),
    .B2(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__or2_1 _0663_ (.A(_0135_),
    .B(_0147_),
    .X(_0153_));
 sky130_fd_sc_hd__a21o_1 _0664_ (.A1(_0135_),
    .A2(_0147_),
    .B1(_0137_),
    .X(_0154_));
 sky130_fd_sc_hd__a21o_1 _0665_ (.A1(_0153_),
    .A2(_0154_),
    .B1(_0139_),
    .X(_0155_));
 sky130_fd_sc_hd__o21ai_1 _0666_ (.A1(_0137_),
    .A2(_0153_),
    .B1(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__a21oi_2 _0667_ (.A1(_0124_),
    .A2(_0156_),
    .B1(_0149_),
    .Y(_0157_));
 sky130_fd_sc_hd__nand2_2 _0668_ (.A(_0113_),
    .B(_0115_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand2_2 _0669_ (.A(\M0.FBM7.q ),
    .B(_0114_),
    .Y(_0159_));
 sky130_fd_sc_hd__xor2_4 _0670_ (.A(_0158_),
    .B(_0159_),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_1 _0671_ (.A(_0157_),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__or2_1 _0672_ (.A(_0141_),
    .B(_0147_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_2 _0673_ (.A(_0148_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__or2_1 _0674_ (.A(_0131_),
    .B(_0163_),
    .X(_0164_));
 sky130_fd_sc_hd__or2_1 _0675_ (.A(_0157_),
    .B(_0160_),
    .X(_0165_));
 sky130_fd_sc_hd__o21a_1 _0676_ (.A1(_0152_),
    .A2(_0165_),
    .B1(_0161_),
    .X(_0166_));
 sky130_fd_sc_hd__or2b_1 _0677_ (.A(_0152_),
    .B_N(_0165_),
    .X(_0167_));
 sky130_fd_sc_hd__o21ai_1 _0678_ (.A1(_0164_),
    .A2(_0166_),
    .B1(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__nand2_1 _0679_ (.A(_0131_),
    .B(_0163_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_1 _0680_ (.A(_0164_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__buf_6 _0681_ (.A(\M0.FAM3.q ),
    .X(_0171_));
 sky130_fd_sc_hd__buf_6 _0682_ (.A(\M0.FAM2.q ),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_2 _0683_ (.A(_0120_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__buf_6 _0684_ (.A(\M0.FAM0.q ),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_2 _0685_ (.A(_0115_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__buf_6 _0686_ (.A(\M0.FAM1.q ),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _0687_ (.A(\M0.FBM7.q ),
    .B(_0176_),
    .X(_0177_));
 sky130_fd_sc_hd__a32oi_4 _0688_ (.A1(_0119_),
    .A2(_0171_),
    .A3(_0173_),
    .B1(_0175_),
    .B2(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_4 _0689_ (.A(_0119_),
    .B(_0172_),
    .Y(_0179_));
 sky130_fd_sc_hd__nand2_2 _0690_ (.A(_0120_),
    .B(_0171_),
    .Y(_0180_));
 sky130_fd_sc_hd__xor2_4 _0691_ (.A(_0179_),
    .B(_0180_),
    .X(_0181_));
 sky130_fd_sc_hd__nand2_2 _0692_ (.A(\M0.FBM7.q ),
    .B(_0174_),
    .Y(_0182_));
 sky130_fd_sc_hd__nand2_2 _0693_ (.A(_0115_),
    .B(_0176_),
    .Y(_0183_));
 sky130_fd_sc_hd__xor2_4 _0694_ (.A(_0182_),
    .B(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_1 _0695_ (.A(_0181_),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__and4_1 _0696_ (.A(\M0.FBM7.q ),
    .B(_0115_),
    .C(_0176_),
    .D(_0174_),
    .X(_0186_));
 sky130_fd_sc_hd__and4_1 _0697_ (.A(_0119_),
    .B(_0120_),
    .C(_0171_),
    .D(_0172_),
    .X(_0187_));
 sky130_fd_sc_hd__xnor2_1 _0698_ (.A(_0186_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand2_1 _0699_ (.A(_0119_),
    .B(_0176_),
    .Y(_0189_));
 sky130_fd_sc_hd__nand2_1 _0700_ (.A(\M0.FBM7.q ),
    .B(_0171_),
    .Y(_0190_));
 sky130_fd_sc_hd__and4bb_2 _0701_ (.A_N(_0189_),
    .B_N(_0190_),
    .C(_0175_),
    .D(_0173_),
    .X(_0191_));
 sky130_fd_sc_hd__inv_2 _0702_ (.A(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__o211a_1 _0703_ (.A1(_0178_),
    .A2(_0185_),
    .B1(_0188_),
    .C1(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__nand2_1 _0704_ (.A(\M0.FBM7.q ),
    .B(_0172_),
    .Y(_0194_));
 sky130_fd_sc_hd__nand2_1 _0705_ (.A(_0115_),
    .B(_0171_),
    .Y(_0195_));
 sky130_fd_sc_hd__xnor2_2 _0706_ (.A(_0194_),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__nor2_1 _0707_ (.A(_0193_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__and2_1 _0708_ (.A(_0115_),
    .B(_0172_),
    .X(_0198_));
 sky130_fd_sc_hd__xnor2_2 _0709_ (.A(_0182_),
    .B(_0183_),
    .Y(_0199_));
 sky130_fd_sc_hd__and2_1 _0710_ (.A(_0115_),
    .B(_0174_),
    .X(_0200_));
 sky130_fd_sc_hd__a22o_1 _0711_ (.A1(_0120_),
    .A2(_0172_),
    .B1(_0176_),
    .B2(_0119_),
    .X(_0201_));
 sky130_fd_sc_hd__and4_1 _0712_ (.A(_0119_),
    .B(_0120_),
    .C(_0172_),
    .D(_0176_),
    .X(_0202_));
 sky130_fd_sc_hd__and4_1 _0713_ (.A(_0119_),
    .B(_0120_),
    .C(_0176_),
    .D(_0174_),
    .X(_0203_));
 sky130_fd_sc_hd__a211o_1 _0714_ (.A1(_0200_),
    .A2(_0201_),
    .B1(_0202_),
    .C1(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__nor2_1 _0715_ (.A(_0181_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__xnor2_2 _0716_ (.A(_0179_),
    .B(_0180_),
    .Y(_0206_));
 sky130_fd_sc_hd__nor3_1 _0717_ (.A(_0206_),
    .B(_0191_),
    .C(_0178_),
    .Y(_0207_));
 sky130_fd_sc_hd__or3_1 _0718_ (.A(_0184_),
    .B(_0191_),
    .C(_0178_),
    .X(_0208_));
 sky130_fd_sc_hd__o31ai_1 _0719_ (.A1(_0199_),
    .A2(_0205_),
    .A3(_0207_),
    .B1(_0208_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _0720_ (.A(_0191_),
    .B(_0178_),
    .Y(_0210_));
 sky130_fd_sc_hd__or2_1 _0721_ (.A(_0172_),
    .B(_0174_),
    .X(_0211_));
 sky130_fd_sc_hd__and2_1 _0722_ (.A(_0119_),
    .B(_0176_),
    .X(_0212_));
 sky130_fd_sc_hd__o211a_1 _0723_ (.A1(_0120_),
    .A2(_0200_),
    .B1(_0211_),
    .C1(_0212_),
    .X(_0213_));
 sky130_fd_sc_hd__a21o_1 _0724_ (.A1(_0213_),
    .A2(_0184_),
    .B1(_0198_),
    .X(_0214_));
 sky130_fd_sc_hd__nor2_2 _0725_ (.A(_0173_),
    .B(_0175_),
    .Y(_0215_));
 sky130_fd_sc_hd__a31o_1 _0726_ (.A1(_0181_),
    .A2(_0199_),
    .A3(_0198_),
    .B1(_0215_),
    .X(_0216_));
 sky130_fd_sc_hd__a32o_1 _0727_ (.A1(_0206_),
    .A2(_0210_),
    .A3(_0214_),
    .B1(_0216_),
    .B2(_0213_),
    .X(_0217_));
 sky130_fd_sc_hd__inv_2 _0728_ (.A(_0215_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_2 _0729_ (.A(_0120_),
    .B(_0174_),
    .Y(_0219_));
 sky130_fd_sc_hd__a31o_1 _0730_ (.A1(_0173_),
    .A2(_0175_),
    .A3(_0219_),
    .B1(_0189_),
    .X(_0220_));
 sky130_fd_sc_hd__or4_1 _0731_ (.A(_0220_),
    .B(_0184_),
    .C(_0191_),
    .D(_0178_),
    .X(_0221_));
 sky130_fd_sc_hd__a21oi_1 _0732_ (.A1(_0218_),
    .A2(_0221_),
    .B1(_0206_),
    .Y(_0222_));
 sky130_fd_sc_hd__a211o_1 _0733_ (.A1(_0198_),
    .A2(_0209_),
    .B1(_0217_),
    .C1(_0222_),
    .X(_0223_));
 sky130_fd_sc_hd__nand2_1 _0734_ (.A(_0193_),
    .B(_0196_),
    .Y(_0224_));
 sky130_fd_sc_hd__o21a_1 _0735_ (.A1(_0197_),
    .A2(_0223_),
    .B1(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__nand2_1 _0736_ (.A(_0184_),
    .B(_0215_),
    .Y(_0226_));
 sky130_fd_sc_hd__a21oi_1 _0737_ (.A1(_0208_),
    .A2(_0226_),
    .B1(_0206_),
    .Y(_0227_));
 sky130_fd_sc_hd__a31oi_1 _0738_ (.A1(_0206_),
    .A2(_0184_),
    .A3(_0210_),
    .B1(_0227_),
    .Y(_0228_));
 sky130_fd_sc_hd__o21ba_1 _0739_ (.A1(_0220_),
    .A2(_0228_),
    .B1_N(_0197_),
    .X(_0229_));
 sky130_fd_sc_hd__nand2_1 _0740_ (.A(_0115_),
    .B(_0172_),
    .Y(_0230_));
 sky130_fd_sc_hd__o21ba_1 _0741_ (.A1(_0230_),
    .A2(_0203_),
    .B1_N(_0190_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_2 _0742_ (.A0(_0225_),
    .A1(_0229_),
    .S(_0231_),
    .X(_0232_));
 sky130_fd_sc_hd__inv_2 _0743_ (.A(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__buf_8 _0744_ (.A(\M0.FBM0.q ),
    .X(_0234_));
 sky130_fd_sc_hd__and2_2 _0745_ (.A(_0114_),
    .B(_0234_),
    .X(_0235_));
 sky130_fd_sc_hd__clkbuf_8 _0746_ (.A(\M0.FBM1.q ),
    .X(_0236_));
 sky130_fd_sc_hd__buf_8 _0747_ (.A(\M0.FBM2.q ),
    .X(_0237_));
 sky130_fd_sc_hd__or2_1 _0748_ (.A(_0237_),
    .B(_0234_),
    .X(_0238_));
 sky130_fd_sc_hd__o2111ai_2 _0749_ (.A1(_0118_),
    .A2(_0235_),
    .B1(_0236_),
    .C1(_0117_),
    .D1(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand2_2 _0750_ (.A(_0113_),
    .B(_0234_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_2 _0751_ (.A(_0114_),
    .B(_0236_),
    .Y(_0241_));
 sky130_fd_sc_hd__xor2_4 _0752_ (.A(_0240_),
    .B(_0241_),
    .X(_0242_));
 sky130_fd_sc_hd__or2_1 _0753_ (.A(_0239_),
    .B(_0242_),
    .X(_0243_));
 sky130_fd_sc_hd__o2111a_1 _0754_ (.A1(_0118_),
    .A2(_0235_),
    .B1(_0236_),
    .C1(_0117_),
    .D1(_0238_),
    .X(_0244_));
 sky130_fd_sc_hd__nand2_1 _0755_ (.A(_0244_),
    .B(_0242_),
    .Y(_0245_));
 sky130_fd_sc_hd__o21a_1 _0756_ (.A1(_0117_),
    .A2(_0235_),
    .B1(_0237_),
    .X(_0246_));
 sky130_fd_sc_hd__clkbuf_8 _0757_ (.A(\M0.FBM3.q ),
    .X(_0247_));
 sky130_fd_sc_hd__nand2_1 _0758_ (.A(_0118_),
    .B(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__nand2_1 _0759_ (.A(_0117_),
    .B(_0237_),
    .Y(_0249_));
 sky130_fd_sc_hd__o21a_1 _0760_ (.A1(_0247_),
    .A2(_0235_),
    .B1(_0118_),
    .X(_0250_));
 sky130_fd_sc_hd__nand2_1 _0761_ (.A(_0117_),
    .B(_0247_),
    .Y(_0251_));
 sky130_fd_sc_hd__or3b_1 _0762_ (.A(_0117_),
    .B(_0247_),
    .C_N(_0237_),
    .X(_0252_));
 sky130_fd_sc_hd__clkinvlp_2 _0763_ (.A(_0118_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand2_2 _0764_ (.A(_0114_),
    .B(_0234_),
    .Y(_0254_));
 sky130_fd_sc_hd__a211o_1 _0765_ (.A1(_0251_),
    .A2(_0252_),
    .B1(_0253_),
    .C1(_0254_),
    .X(_0255_));
 sky130_fd_sc_hd__o221a_1 _0766_ (.A1(_0246_),
    .A2(_0248_),
    .B1(_0249_),
    .B2(_0250_),
    .C1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_2 _0767_ (.A0(_0243_),
    .A1(_0245_),
    .S(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__and2_1 _0768_ (.A(_0114_),
    .B(_0237_),
    .X(_0258_));
 sky130_fd_sc_hd__nand2_2 _0769_ (.A(_0118_),
    .B(_0237_),
    .Y(_0259_));
 sky130_fd_sc_hd__xnor2_1 _0770_ (.A(_0117_),
    .B(_0247_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _0771_ (.A(_0113_),
    .B(_0236_),
    .Y(_0261_));
 sky130_fd_sc_hd__a311o_1 _0772_ (.A1(_0117_),
    .A2(_0247_),
    .A3(_0259_),
    .B1(_0235_),
    .C1(_0261_),
    .X(_0262_));
 sky130_fd_sc_hd__and2_1 _0773_ (.A(_0113_),
    .B(_0236_),
    .X(_0263_));
 sky130_fd_sc_hd__a221o_1 _0774_ (.A1(_0118_),
    .A2(_0237_),
    .B1(_0254_),
    .B2(_0263_),
    .C1(_0251_),
    .X(_0264_));
 sky130_fd_sc_hd__o311a_1 _0775_ (.A1(_0259_),
    .A2(_0254_),
    .A3(_0260_),
    .B1(_0262_),
    .C1(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__nand2_1 _0776_ (.A(_0264_),
    .B(_0262_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _0777_ (.A(_0253_),
    .B(_0249_),
    .Y(_0267_));
 sky130_fd_sc_hd__nor2_1 _0778_ (.A(_0117_),
    .B(_0247_),
    .Y(_0268_));
 sky130_fd_sc_hd__and4_1 _0779_ (.A(_0117_),
    .B(_0118_),
    .C(_0247_),
    .D(_0237_),
    .X(_0269_));
 sky130_fd_sc_hd__o21ai_1 _0780_ (.A1(_0268_),
    .A2(_0269_),
    .B1(_0254_),
    .Y(_0270_));
 sky130_fd_sc_hd__o2111a_1 _0781_ (.A1(_0247_),
    .A2(_0237_),
    .B1(_0242_),
    .C1(_0267_),
    .D1(_0270_),
    .X(_0271_));
 sky130_fd_sc_hd__mux2_1 _0782_ (.A0(_0265_),
    .A1(_0266_),
    .S(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__xnor2_1 _0783_ (.A(_0258_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__xnor2_2 _0784_ (.A(_0257_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__and2_1 _0785_ (.A(_0118_),
    .B(_0120_),
    .X(_0275_));
 sky130_fd_sc_hd__and2_1 _0786_ (.A(_0174_),
    .B(_0234_),
    .X(_0276_));
 sky130_fd_sc_hd__buf_1 _0787_ (.A(_0276_),
    .X(\M0.FPM0.d ));
 sky130_fd_sc_hd__and2_1 _0788_ (.A(_0275_),
    .B(\M0.FPM0.d ),
    .X(_0277_));
 sky130_fd_sc_hd__nand2_1 _0789_ (.A(_0119_),
    .B(_0174_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _0790_ (.A(_0120_),
    .B(_0176_),
    .Y(_0279_));
 sky130_fd_sc_hd__xor2_1 _0791_ (.A(_0278_),
    .B(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__nor2_1 _0792_ (.A(_0277_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _0793_ (.A(_0117_),
    .B(_0234_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _0794_ (.A(_0118_),
    .B(_0236_),
    .Y(_0283_));
 sky130_fd_sc_hd__xor2_2 _0795_ (.A(_0282_),
    .B(_0283_),
    .X(_0284_));
 sky130_fd_sc_hd__a21oi_1 _0796_ (.A1(_0277_),
    .A2(_0280_),
    .B1(_0284_),
    .Y(_0285_));
 sky130_fd_sc_hd__nand2_1 _0797_ (.A(_0117_),
    .B(_0236_),
    .Y(_0286_));
 sky130_fd_sc_hd__o211a_1 _0798_ (.A1(_0118_),
    .A2(_0286_),
    .B1(_0259_),
    .C1(_0114_),
    .X(_0287_));
 sky130_fd_sc_hd__and2b_1 _0799_ (.A_N(_0237_),
    .B(_0118_),
    .X(_0288_));
 sky130_fd_sc_hd__o21ai_1 _0800_ (.A1(_0114_),
    .A2(_0288_),
    .B1(_0234_),
    .Y(_0289_));
 sky130_fd_sc_hd__o211a_1 _0801_ (.A1(_0118_),
    .A2(_0235_),
    .B1(_0286_),
    .C1(_0238_),
    .X(_0290_));
 sky130_fd_sc_hd__o21ba_1 _0802_ (.A1(_0234_),
    .A2(_0259_),
    .B1_N(_0286_),
    .X(_0291_));
 sky130_fd_sc_hd__o22a_1 _0803_ (.A1(_0287_),
    .A2(_0289_),
    .B1(_0290_),
    .B2(_0291_),
    .X(_0292_));
 sky130_fd_sc_hd__inv_2 _0804_ (.A(_0174_),
    .Y(_0293_));
 sky130_fd_sc_hd__and4_1 _0805_ (.A(_0120_),
    .B(_0172_),
    .C(_0293_),
    .D(_0212_),
    .X(_0294_));
 sky130_fd_sc_hd__and3b_1 _0806_ (.A_N(_0201_),
    .B(_0219_),
    .C(_0175_),
    .X(_0295_));
 sky130_fd_sc_hd__and2b_1 _0807_ (.A_N(_0172_),
    .B(_0120_),
    .X(_0296_));
 sky130_fd_sc_hd__a21bo_1 _0808_ (.A1(_0120_),
    .A2(_0172_),
    .B1_N(_0115_),
    .X(_0297_));
 sky130_fd_sc_hd__and3b_1 _0809_ (.A_N(_0120_),
    .B(_0176_),
    .C(_0119_),
    .X(_0298_));
 sky130_fd_sc_hd__o221a_1 _0810_ (.A1(_0115_),
    .A2(_0296_),
    .B1(_0297_),
    .B2(_0298_),
    .C1(_0174_),
    .X(_0299_));
 sky130_fd_sc_hd__nor3_1 _0811_ (.A(_0294_),
    .B(_0295_),
    .C(_0299_),
    .Y(_0300_));
 sky130_fd_sc_hd__a2bb2o_1 _0812_ (.A1_N(_0281_),
    .A2_N(_0285_),
    .B1(_0292_),
    .B2(_0300_),
    .X(_0301_));
 sky130_fd_sc_hd__or2_1 _0813_ (.A(_0292_),
    .B(_0300_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _0814_ (.A(_0239_),
    .B(_0242_),
    .Y(_0303_));
 sky130_fd_sc_hd__or2_1 _0815_ (.A(_0244_),
    .B(_0242_),
    .X(_0304_));
 sky130_fd_sc_hd__mux2_1 _0816_ (.A0(_0303_),
    .A1(_0304_),
    .S(_0256_),
    .X(_0305_));
 sky130_fd_sc_hd__a22o_1 _0817_ (.A1(_0301_),
    .A2(_0302_),
    .B1(_0257_),
    .B2(_0305_),
    .X(_0306_));
 sky130_fd_sc_hd__xnor2_1 _0818_ (.A(_0181_),
    .B(_0215_),
    .Y(_0307_));
 sky130_fd_sc_hd__xnor2_1 _0819_ (.A(_0213_),
    .B(_0199_),
    .Y(_0308_));
 sky130_fd_sc_hd__xnor2_2 _0820_ (.A(_0307_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__a41o_1 _0821_ (.A1(_0301_),
    .A2(_0302_),
    .A3(_0257_),
    .A4(_0305_),
    .B1(_0309_),
    .X(_0310_));
 sky130_fd_sc_hd__and2_1 _0822_ (.A(_0306_),
    .B(_0310_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _0823_ (.A(_0274_),
    .B(_0311_),
    .X(_0312_));
 sky130_fd_sc_hd__a211oi_1 _0824_ (.A1(_0208_),
    .A2(_0185_),
    .B1(_0218_),
    .C1(_0189_),
    .Y(_0313_));
 sky130_fd_sc_hd__a21o_1 _0825_ (.A1(_0181_),
    .A2(_0184_),
    .B1(_0204_),
    .X(_0314_));
 sky130_fd_sc_hd__a211o_1 _0826_ (.A1(_0212_),
    .A2(_0215_),
    .B1(_0184_),
    .C1(_0181_),
    .X(_0315_));
 sky130_fd_sc_hd__a21oi_1 _0827_ (.A1(_0314_),
    .A2(_0315_),
    .B1(_0210_),
    .Y(_0316_));
 sky130_fd_sc_hd__or2_1 _0828_ (.A(_0184_),
    .B(_0204_),
    .X(_0317_));
 sky130_fd_sc_hd__a32o_1 _0829_ (.A1(_0213_),
    .A2(_0184_),
    .A3(_0210_),
    .B1(_0207_),
    .B2(_0317_),
    .X(_0318_));
 sky130_fd_sc_hd__o31ai_1 _0830_ (.A1(_0313_),
    .A2(_0316_),
    .A3(_0318_),
    .B1(_0198_),
    .Y(_0319_));
 sky130_fd_sc_hd__or4_1 _0831_ (.A(_0198_),
    .B(_0313_),
    .C(_0316_),
    .D(_0318_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_1 _0832_ (.A(_0319_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__a21o_1 _0833_ (.A1(_0274_),
    .A2(_0311_),
    .B1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__nand2_2 _0834_ (.A(_0312_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor2_1 _0835_ (.A(_0257_),
    .B(_0272_),
    .Y(_0324_));
 sky130_fd_sc_hd__nand2_1 _0836_ (.A(_0257_),
    .B(_0272_),
    .Y(_0325_));
 sky130_fd_sc_hd__o21a_1 _0837_ (.A1(_0258_),
    .A2(_0324_),
    .B1(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0838_ (.A(_0113_),
    .B(_0237_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _0839_ (.A(_0114_),
    .B(_0247_),
    .Y(_0328_));
 sky130_fd_sc_hd__xor2_2 _0840_ (.A(_0327_),
    .B(_0328_),
    .X(_0329_));
 sky130_fd_sc_hd__inv_2 _0841_ (.A(_0117_),
    .Y(_0330_));
 sky130_fd_sc_hd__and2_1 _0842_ (.A(_0253_),
    .B(_0237_),
    .X(_0331_));
 sky130_fd_sc_hd__a31o_1 _0843_ (.A1(_0118_),
    .A2(_0254_),
    .A3(_0263_),
    .B1(_0117_),
    .X(_0332_));
 sky130_fd_sc_hd__o311a_1 _0844_ (.A1(_0330_),
    .A2(_0288_),
    .A3(_0331_),
    .B1(_0332_),
    .C1(_0242_),
    .X(_0333_));
 sky130_fd_sc_hd__a41o_1 _0845_ (.A1(_0117_),
    .A2(_0259_),
    .A3(_0254_),
    .A4(_0263_),
    .B1(_0333_),
    .X(_0334_));
 sky130_fd_sc_hd__nor2_1 _0846_ (.A(_0247_),
    .B(_0249_),
    .Y(_0335_));
 sky130_fd_sc_hd__and4_1 _0847_ (.A(_0113_),
    .B(_0114_),
    .C(_0236_),
    .D(_0234_),
    .X(_0336_));
 sky130_fd_sc_hd__xor2_1 _0848_ (.A(_0269_),
    .B(_0336_),
    .X(_0337_));
 sky130_fd_sc_hd__a41o_1 _0849_ (.A1(_0254_),
    .A2(_0242_),
    .A3(_0263_),
    .A4(_0335_),
    .B1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__a21o_1 _0850_ (.A1(_0247_),
    .A2(_0334_),
    .B1(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__xnor2_1 _0851_ (.A(_0329_),
    .B(_0339_),
    .Y(_0340_));
 sky130_fd_sc_hd__xnor2_2 _0852_ (.A(_0326_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__xnor2_1 _0853_ (.A(_0193_),
    .B(_0196_),
    .Y(_0342_));
 sky130_fd_sc_hd__xnor2_2 _0854_ (.A(_0223_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__xor2_2 _0855_ (.A(_0341_),
    .B(_0343_),
    .X(_0344_));
 sky130_fd_sc_hd__xnor2_4 _0856_ (.A(_0323_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__and4_1 _0857_ (.A(_0171_),
    .B(_0172_),
    .C(_0236_),
    .D(_0234_),
    .X(_0346_));
 sky130_fd_sc_hd__and4_1 _0858_ (.A(_0176_),
    .B(_0174_),
    .C(_0247_),
    .D(_0237_),
    .X(_0347_));
 sky130_fd_sc_hd__xnor2_2 _0859_ (.A(_0346_),
    .B(_0347_),
    .Y(_0348_));
 sky130_fd_sc_hd__and2_2 _0860_ (.A(_0174_),
    .B(_0237_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_2 _0861_ (.A(_0176_),
    .B(_0247_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_2 _0862_ (.A(_0172_),
    .B(_0234_),
    .Y(_0351_));
 sky130_fd_sc_hd__o2111a_1 _0863_ (.A1(_0349_),
    .A2(_0350_),
    .B1(_0351_),
    .C1(_0171_),
    .D1(_0236_),
    .X(_0352_));
 sky130_fd_sc_hd__a311oi_4 _0864_ (.A1(_0171_),
    .A2(_0236_),
    .A3(_0351_),
    .B1(_0350_),
    .C1(_0349_),
    .Y(_0353_));
 sky130_fd_sc_hd__or2_2 _0865_ (.A(_0352_),
    .B(_0353_),
    .X(_0354_));
 sky130_fd_sc_hd__and4_2 _0866_ (.A(_0172_),
    .B(_0174_),
    .C(_0237_),
    .D(_0234_),
    .X(_0355_));
 sky130_fd_sc_hd__nand2_2 _0867_ (.A(_0176_),
    .B(_0237_),
    .Y(_0356_));
 sky130_fd_sc_hd__nand2_2 _0868_ (.A(_0174_),
    .B(_0247_),
    .Y(_0357_));
 sky130_fd_sc_hd__xor2_4 _0869_ (.A(_0356_),
    .B(_0357_),
    .X(_0358_));
 sky130_fd_sc_hd__nand2_2 _0870_ (.A(_0171_),
    .B(_0234_),
    .Y(_0359_));
 sky130_fd_sc_hd__nand2_2 _0871_ (.A(_0172_),
    .B(_0236_),
    .Y(_0360_));
 sky130_fd_sc_hd__xor2_4 _0872_ (.A(_0359_),
    .B(_0360_),
    .X(_0361_));
 sky130_fd_sc_hd__xor2_4 _0873_ (.A(_0358_),
    .B(_0361_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_2 _0874_ (.A(_0176_),
    .B(_0236_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _0875_ (.A(_0174_),
    .B(_0237_),
    .Y(_0364_));
 sky130_fd_sc_hd__nor2_1 _0876_ (.A(_0234_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__a31o_1 _0877_ (.A1(_0172_),
    .A2(_0293_),
    .A3(_0234_),
    .B1(_0365_),
    .X(_0366_));
 sky130_fd_sc_hd__o2111ai_4 _0878_ (.A1(_0354_),
    .A2(_0355_),
    .B1(_0362_),
    .C1(_0363_),
    .D1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__and3_1 _0879_ (.A(_0171_),
    .B(_0236_),
    .C(_0351_),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_1 _0880_ (.A(_0349_),
    .B(_0350_),
    .Y(_0369_));
 sky130_fd_sc_hd__a22o_1 _0881_ (.A1(_0358_),
    .A2(_0361_),
    .B1(_0368_),
    .B2(_0369_),
    .X(_0370_));
 sky130_fd_sc_hd__nand2_1 _0882_ (.A(_0176_),
    .B(_0236_),
    .Y(_0371_));
 sky130_fd_sc_hd__or3_1 _0883_ (.A(_0371_),
    .B(_0364_),
    .C(_0351_),
    .X(_0372_));
 sky130_fd_sc_hd__or3b_1 _0884_ (.A(_0368_),
    .B(_0369_),
    .C_N(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_2 _0885_ (.A(_0370_),
    .B(_0373_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_1 _0886_ (.A(_0171_),
    .B(_0237_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _0887_ (.A(_0172_),
    .B(_0247_),
    .Y(_0376_));
 sky130_fd_sc_hd__xor2_2 _0888_ (.A(_0375_),
    .B(_0376_),
    .X(_0377_));
 sky130_fd_sc_hd__and3b_1 _0889_ (.A_N(_0348_),
    .B(_0362_),
    .C(_0354_),
    .X(_0378_));
 sky130_fd_sc_hd__a311o_1 _0890_ (.A1(_0348_),
    .A2(_0367_),
    .A3(_0374_),
    .B1(_0377_),
    .C1(_0378_),
    .X(_0379_));
 sky130_fd_sc_hd__and2_1 _0891_ (.A(_0363_),
    .B(\M0.FPM0.d ),
    .X(_0380_));
 sky130_fd_sc_hd__and3_1 _0892_ (.A(_0362_),
    .B(_0354_),
    .C(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__a41oi_4 _0893_ (.A1(_0348_),
    .A2(_0367_),
    .A3(_0374_),
    .A4(_0377_),
    .B1(_0381_),
    .Y(_0382_));
 sky130_fd_sc_hd__and2_1 _0894_ (.A(_0379_),
    .B(_0382_),
    .X(_0383_));
 sky130_fd_sc_hd__a21oi_1 _0895_ (.A1(_0234_),
    .A2(_0211_),
    .B1(_0349_),
    .Y(_0384_));
 sky130_fd_sc_hd__nor2_1 _0896_ (.A(_0371_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a211o_1 _0897_ (.A1(_0361_),
    .A2(_0355_),
    .B1(_0353_),
    .C1(_0352_),
    .X(_0386_));
 sky130_fd_sc_hd__xor2_1 _0898_ (.A(_0361_),
    .B(_0355_),
    .X(_0387_));
 sky130_fd_sc_hd__a22o_1 _0899_ (.A1(_0358_),
    .A2(_0386_),
    .B1(_0387_),
    .B2(_0354_),
    .X(_0388_));
 sky130_fd_sc_hd__nor2_1 _0900_ (.A(_0352_),
    .B(_0353_),
    .Y(_0389_));
 sky130_fd_sc_hd__nor3b_1 _0901_ (.A(_0358_),
    .B(_0361_),
    .C_N(_0372_),
    .Y(_0390_));
 sky130_fd_sc_hd__and4_1 _0902_ (.A(_0176_),
    .B(_0174_),
    .C(_0237_),
    .D(_0236_),
    .X(_0391_));
 sky130_fd_sc_hd__a311o_1 _0903_ (.A1(_0234_),
    .A2(_0211_),
    .A3(_0363_),
    .B1(_0355_),
    .C1(_0391_),
    .X(_0392_));
 sky130_fd_sc_hd__inv_2 _0904_ (.A(_0392_),
    .Y(_0393_));
 sky130_fd_sc_hd__a211oi_1 _0905_ (.A1(_0358_),
    .A2(_0361_),
    .B1(_0352_),
    .C1(_0353_),
    .Y(_0394_));
 sky130_fd_sc_hd__o211a_1 _0906_ (.A1(_0352_),
    .A2(_0353_),
    .B1(_0358_),
    .C1(_0361_),
    .X(_0395_));
 sky130_fd_sc_hd__a221o_1 _0907_ (.A1(_0389_),
    .A2(_0390_),
    .B1(_0393_),
    .B2(_0394_),
    .C1(_0395_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_2 _0908_ (.A(_0172_),
    .B(_0237_),
    .Y(_0397_));
 sky130_fd_sc_hd__a211o_1 _0909_ (.A1(_0385_),
    .A2(_0388_),
    .B1(_0396_),
    .C1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _0910_ (.A(_0118_),
    .B(_0234_),
    .Y(_0399_));
 sky130_fd_sc_hd__xnor2_2 _0911_ (.A(_0219_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__a22o_1 _0912_ (.A1(_0389_),
    .A2(_0390_),
    .B1(_0393_),
    .B2(_0394_),
    .X(_0401_));
 sky130_fd_sc_hd__and3_1 _0913_ (.A(_0358_),
    .B(_0385_),
    .C(_0386_),
    .X(_0402_));
 sky130_fd_sc_hd__a31o_1 _0914_ (.A1(_0354_),
    .A2(_0385_),
    .A3(_0387_),
    .B1(_0395_),
    .X(_0403_));
 sky130_fd_sc_hd__o31a_1 _0915_ (.A1(_0401_),
    .A2(_0402_),
    .A3(_0403_),
    .B1(_0397_),
    .X(_0404_));
 sky130_fd_sc_hd__a21o_1 _0916_ (.A1(_0398_),
    .A2(_0400_),
    .B1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__and2_1 _0917_ (.A(_0277_),
    .B(_0280_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_1 _0918_ (.A(_0281_),
    .B(_0406_),
    .Y(_0407_));
 sky130_fd_sc_hd__xnor2_2 _0919_ (.A(_0284_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__a211o_1 _0920_ (.A1(_0379_),
    .A2(_0382_),
    .B1(_0400_),
    .C1(_0404_),
    .X(_0409_));
 sky130_fd_sc_hd__a21oi_1 _0921_ (.A1(_0379_),
    .A2(_0382_),
    .B1(_0398_),
    .Y(_0410_));
 sky130_fd_sc_hd__a221oi_4 _0922_ (.A1(_0383_),
    .A2(_0405_),
    .B1(_0408_),
    .B2(_0409_),
    .C1(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__a21o_1 _0923_ (.A1(_0379_),
    .A2(_0382_),
    .B1(_0398_),
    .X(_0412_));
 sky130_fd_sc_hd__inv_2 _0924_ (.A(_0377_),
    .Y(_0413_));
 sky130_fd_sc_hd__a311o_1 _0925_ (.A1(_0348_),
    .A2(_0367_),
    .A3(_0374_),
    .B1(_0413_),
    .C1(_0381_),
    .X(_0414_));
 sky130_fd_sc_hd__nand2_1 _0926_ (.A(_0171_),
    .B(_0247_),
    .Y(_0415_));
 sky130_fd_sc_hd__o21ba_1 _0927_ (.A1(_0397_),
    .A2(_0380_),
    .B1_N(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__or2b_1 _0928_ (.A(_0415_),
    .B_N(_0397_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(_0416_),
    .A1(_0417_),
    .S(_0378_),
    .X(_0418_));
 sky130_fd_sc_hd__xor2_1 _0930_ (.A(_0414_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__or2_1 _0931_ (.A(_0281_),
    .B(_0285_),
    .X(_0420_));
 sky130_fd_sc_hd__xnor2_1 _0932_ (.A(_0292_),
    .B(net36),
    .Y(_0421_));
 sky130_fd_sc_hd__xnor2_2 _0933_ (.A(_0420_),
    .B(_0421_),
    .Y(_0422_));
 sky130_fd_sc_hd__nand3_1 _0934_ (.A(_0412_),
    .B(_0419_),
    .C(_0422_),
    .Y(_0423_));
 sky130_fd_sc_hd__a21oi_1 _0935_ (.A1(_0412_),
    .A2(_0419_),
    .B1(_0422_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand2_1 _0936_ (.A(_0257_),
    .B(_0305_),
    .Y(_0425_));
 sky130_fd_sc_hd__nand3_1 _0937_ (.A(_0301_),
    .B(_0302_),
    .C(_0309_),
    .Y(_0426_));
 sky130_fd_sc_hd__a21o_1 _0938_ (.A1(_0301_),
    .A2(_0302_),
    .B1(_0309_),
    .X(_0427_));
 sky130_fd_sc_hd__nand3_1 _0939_ (.A(_0425_),
    .B(_0426_),
    .C(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21o_1 _0940_ (.A1(_0426_),
    .A2(_0427_),
    .B1(_0425_),
    .X(_0429_));
 sky130_fd_sc_hd__clkinvlp_2 _0941_ (.A(_0378_),
    .Y(_0430_));
 sky130_fd_sc_hd__a31o_1 _0942_ (.A1(_0397_),
    .A2(_0430_),
    .A3(_0414_),
    .B1(_0415_),
    .X(_0431_));
 sky130_fd_sc_hd__a21oi_1 _0943_ (.A1(_0428_),
    .A2(_0429_),
    .B1(_0431_),
    .Y(_0432_));
 sky130_fd_sc_hd__a211o_1 _0944_ (.A1(_0411_),
    .A2(_0423_),
    .B1(_0424_),
    .C1(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__nand3_2 _0945_ (.A(_0431_),
    .B(_0428_),
    .C(_0429_),
    .Y(_0434_));
 sky130_fd_sc_hd__xnor2_1 _0946_ (.A(_0274_),
    .B(_0321_),
    .Y(_0435_));
 sky130_fd_sc_hd__xnor2_2 _0947_ (.A(_0311_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__and3_2 _0948_ (.A(_0433_),
    .B(_0434_),
    .C(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__nand2_4 _0949_ (.A(_0345_),
    .B(_0437_),
    .Y(_0438_));
 sky130_fd_sc_hd__nor2_1 _0950_ (.A(_0233_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a21o_1 _0951_ (.A1(_0230_),
    .A2(_0229_),
    .B1(_0190_),
    .X(_0440_));
 sky130_fd_sc_hd__a31o_1 _0952_ (.A1(_0312_),
    .A2(_0322_),
    .A3(_0343_),
    .B1(_0341_),
    .X(_0441_));
 sky130_fd_sc_hd__a21o_1 _0953_ (.A1(_0312_),
    .A2(_0322_),
    .B1(_0343_),
    .X(_0442_));
 sky130_fd_sc_hd__nand2_1 _0954_ (.A(_0114_),
    .B(_0237_),
    .Y(_0443_));
 sky130_fd_sc_hd__a41o_1 _0955_ (.A1(_0117_),
    .A2(_0118_),
    .A3(_0236_),
    .A4(_0234_),
    .B1(_0443_),
    .X(_0444_));
 sky130_fd_sc_hd__and3_1 _0956_ (.A(_0113_),
    .B(_0247_),
    .C(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__or2_1 _0957_ (.A(_0329_),
    .B(_0445_),
    .X(_0446_));
 sky130_fd_sc_hd__a21o_1 _0958_ (.A1(_0258_),
    .A2(_0325_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__nand2_1 _0959_ (.A(_0329_),
    .B(_0445_),
    .Y(_0448_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(_0446_),
    .A1(_0448_),
    .S(_0339_),
    .X(_0449_));
 sky130_fd_sc_hd__o311a_2 _0961_ (.A1(_0326_),
    .A2(_0339_),
    .A3(_0445_),
    .B1(_0447_),
    .C1(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__a21oi_1 _0962_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__o21a_1 _0963_ (.A1(_0324_),
    .A2(_0339_),
    .B1(_0329_),
    .X(_0452_));
 sky130_fd_sc_hd__o211ai_2 _0964_ (.A1(_0258_),
    .A2(_0452_),
    .B1(_0113_),
    .C1(_0247_),
    .Y(_0453_));
 sky130_fd_sc_hd__o21a_1 _0965_ (.A1(_0440_),
    .A2(_0451_),
    .B1(_0453_),
    .X(_0454_));
 sky130_fd_sc_hd__a21oi_1 _0966_ (.A1(_0440_),
    .A2(_0451_),
    .B1(_0454_),
    .Y(_0455_));
 sky130_fd_sc_hd__and3_1 _0967_ (.A(_0441_),
    .B(_0442_),
    .C(_0450_),
    .X(_0456_));
 sky130_fd_sc_hd__a21o_1 _0968_ (.A1(_0233_),
    .A2(_0438_),
    .B1(_0440_),
    .X(_0457_));
 sky130_fd_sc_hd__and3_1 _0969_ (.A(_0233_),
    .B(_0438_),
    .C(_0440_),
    .X(_0458_));
 sky130_fd_sc_hd__a21oi_1 _0970_ (.A1(_0453_),
    .A2(_0457_),
    .B1(_0458_),
    .Y(_0459_));
 sky130_fd_sc_hd__o22a_2 _0971_ (.A1(_0439_),
    .A2(_0455_),
    .B1(_0456_),
    .B2(_0459_),
    .X(_0460_));
 sky130_fd_sc_hd__or2_1 _0972_ (.A(_0232_),
    .B(_0450_),
    .X(_0461_));
 sky130_fd_sc_hd__a22o_1 _0973_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0450_),
    .B2(_0232_),
    .X(_0462_));
 sky130_fd_sc_hd__a22oi_2 _0974_ (.A1(_0345_),
    .A2(_0437_),
    .B1(_0461_),
    .B2(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__and2_1 _0975_ (.A(_0233_),
    .B(_0451_),
    .X(_0464_));
 sky130_fd_sc_hd__and4_1 _0976_ (.A(_0232_),
    .B(_0345_),
    .C(_0437_),
    .D(_0456_),
    .X(_0465_));
 sky130_fd_sc_hd__xor2_1 _0977_ (.A(_0453_),
    .B(_0440_),
    .X(_0466_));
 sky130_fd_sc_hd__o31ai_2 _0978_ (.A1(_0463_),
    .A2(_0464_),
    .A3(_0465_),
    .B1(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__or4_1 _0979_ (.A(_0463_),
    .B(_0464_),
    .C(_0465_),
    .D(_0466_),
    .X(_0468_));
 sky130_fd_sc_hd__xor2_1 _0980_ (.A(_0232_),
    .B(_0450_),
    .X(_0469_));
 sky130_fd_sc_hd__a21oi_1 _0981_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0469_),
    .Y(_0470_));
 sky130_fd_sc_hd__and3_1 _0982_ (.A(_0441_),
    .B(_0442_),
    .C(_0469_),
    .X(_0471_));
 sky130_fd_sc_hd__nor2_2 _0983_ (.A(_0470_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__o21ai_1 _0984_ (.A1(_0118_),
    .A2(_0142_),
    .B1(_0138_),
    .Y(_0473_));
 sky130_fd_sc_hd__nor2_1 _0985_ (.A(_0114_),
    .B(_0115_),
    .Y(_0474_));
 sky130_fd_sc_hd__a22o_1 _0986_ (.A1(_0114_),
    .A2(_0473_),
    .B1(_0474_),
    .B2(_0118_),
    .X(_0475_));
 sky130_fd_sc_hd__nor2_1 _0987_ (.A(_0120_),
    .B(_0138_),
    .Y(_0476_));
 sky130_fd_sc_hd__a2bb2o_1 _0988_ (.A1_N(_0115_),
    .A2_N(_0120_),
    .B1(_0136_),
    .B2(_0253_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_1 _0989_ (.A0(_0476_),
    .A1(_0477_),
    .S(_0142_),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_4 _0990_ (.A1(_0120_),
    .A2(_0475_),
    .B1(_0478_),
    .Y(_0479_));
 sky130_fd_sc_hd__nand2_1 _0991_ (.A(_0117_),
    .B(_0120_),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_1 _0992_ (.A(_0118_),
    .B(_0119_),
    .Y(_0481_));
 sky130_fd_sc_hd__xor2_2 _0993_ (.A(_0480_),
    .B(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__o2111a_1 _0994_ (.A1(_0275_),
    .A2(_0436_),
    .B1(_0482_),
    .C1(_0433_),
    .D1(_0434_),
    .X(_0483_));
 sky130_fd_sc_hd__a311o_1 _0995_ (.A1(_0275_),
    .A2(_0436_),
    .A3(_0482_),
    .B1(_0483_),
    .C1(_0345_),
    .X(_0484_));
 sky130_fd_sc_hd__a21oi_1 _0996_ (.A1(_0433_),
    .A2(_0434_),
    .B1(_0436_),
    .Y(_0485_));
 sky130_fd_sc_hd__o21bai_2 _0997_ (.A1(_0132_),
    .A2(_0485_),
    .B1_N(_0482_),
    .Y(_0486_));
 sky130_fd_sc_hd__o2111ai_4 _0998_ (.A1(_0472_),
    .A2(_0479_),
    .B1(_0438_),
    .C1(_0484_),
    .D1(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__o2111a_1 _0999_ (.A1(_0470_),
    .A2(_0471_),
    .B1(_0479_),
    .C1(_0437_),
    .D1(_0345_),
    .X(_0488_));
 sky130_fd_sc_hd__a31oi_2 _1000_ (.A1(_0438_),
    .A2(_0472_),
    .A3(_0479_),
    .B1(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__a22o_1 _1001_ (.A1(_0467_),
    .A2(_0468_),
    .B1(_0487_),
    .B2(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__nor3_1 _1002_ (.A(_0121_),
    .B(_0146_),
    .C(_0144_),
    .Y(_0491_));
 sky130_fd_sc_hd__or2_1 _1003_ (.A(_0147_),
    .B(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__a41o_1 _1004_ (.A1(_0467_),
    .A2(_0468_),
    .A3(_0487_),
    .A4(_0489_),
    .B1(_0492_),
    .X(_0493_));
 sky130_fd_sc_hd__and2_1 _1005_ (.A(_0490_),
    .B(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__and2b_1 _1006_ (.A_N(_0460_),
    .B(_0494_),
    .X(_0495_));
 sky130_fd_sc_hd__nand2b_1 _1007_ (.A_N(_0494_),
    .B(_0460_),
    .Y(_0496_));
 sky130_fd_sc_hd__o21ai_1 _1008_ (.A1(_0170_),
    .A2(_0495_),
    .B1(_0496_),
    .Y(_0497_));
 sky130_fd_sc_hd__a2bb2o_1 _1009_ (.A1_N(_0152_),
    .A2_N(_0161_),
    .B1(_0168_),
    .B2(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__a311o_1 _1010_ (.A1(_0113_),
    .A2(\M0.FBM7.q ),
    .A3(_0116_),
    .B1(_0150_),
    .C1(_0498_),
    .X(\M0.FPM15.d ));
 sky130_fd_sc_hd__a21o_1 _1011_ (.A1(_0490_),
    .A2(_0493_),
    .B1(_0163_),
    .X(_0499_));
 sky130_fd_sc_hd__nand3_2 _1012_ (.A(_0163_),
    .B(_0490_),
    .C(_0493_),
    .Y(_0500_));
 sky130_fd_sc_hd__a21bo_1 _1013_ (.A1(_0131_),
    .A2(_0499_),
    .B1_N(_0500_),
    .X(_0501_));
 sky130_fd_sc_hd__a21boi_1 _1014_ (.A1(_0161_),
    .A2(_0501_),
    .B1_N(_0165_),
    .Y(_0502_));
 sky130_fd_sc_hd__nor2_1 _1015_ (.A(_0163_),
    .B(_0494_),
    .Y(_0503_));
 sky130_fd_sc_hd__a21o_1 _1016_ (.A1(_0160_),
    .A2(_0500_),
    .B1(_0116_),
    .X(_0504_));
 sky130_fd_sc_hd__o21a_1 _1017_ (.A1(_0160_),
    .A2(_0503_),
    .B1(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__or3_1 _1018_ (.A(_0116_),
    .B(_0160_),
    .C(_0500_),
    .X(_0506_));
 sky130_fd_sc_hd__o221ai_1 _1019_ (.A1(_0460_),
    .A2(_0502_),
    .B1(_0505_),
    .B2(_0157_),
    .C1(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__a21oi_1 _1020_ (.A1(_0152_),
    .A2(_0507_),
    .B1(_0498_),
    .Y(\M0.FPM14.d ));
 sky130_fd_sc_hd__o21a_1 _1021_ (.A1(_0460_),
    .A2(_0503_),
    .B1(_0500_),
    .X(_0508_));
 sky130_fd_sc_hd__or3b_1 _1022_ (.A(_0164_),
    .B(_0494_),
    .C_N(_0460_),
    .X(_0509_));
 sky130_fd_sc_hd__o221a_1 _1023_ (.A1(_0460_),
    .A2(_0500_),
    .B1(_0508_),
    .B2(_0116_),
    .C1(_0509_),
    .X(_0510_));
 sky130_fd_sc_hd__xnor2_1 _1024_ (.A(_0157_),
    .B(_0160_),
    .Y(_0511_));
 sky130_fd_sc_hd__xnor2_1 _1025_ (.A(_0510_),
    .B(_0511_),
    .Y(\M0.FPM13.d ));
 sky130_fd_sc_hd__xnor2_1 _1026_ (.A(_0170_),
    .B(_0460_),
    .Y(_0512_));
 sky130_fd_sc_hd__xnor2_1 _1027_ (.A(_0494_),
    .B(_0512_),
    .Y(\M0.FPM12.d ));
 sky130_fd_sc_hd__nand2_1 _1028_ (.A(_0487_),
    .B(_0489_),
    .Y(_0513_));
 sky130_fd_sc_hd__nand2_1 _1029_ (.A(_0467_),
    .B(_0468_),
    .Y(_0514_));
 sky130_fd_sc_hd__xnor2_1 _1030_ (.A(_0514_),
    .B(_0492_),
    .Y(_0515_));
 sky130_fd_sc_hd__xor2_1 _1031_ (.A(_0513_),
    .B(_0515_),
    .X(\M0.FPM11.d ));
 sky130_fd_sc_hd__nand3_1 _1032_ (.A(_0438_),
    .B(_0484_),
    .C(_0486_),
    .Y(_0516_));
 sky130_fd_sc_hd__xnor2_1 _1033_ (.A(_0438_),
    .B(_0472_),
    .Y(_0517_));
 sky130_fd_sc_hd__nor2_1 _1034_ (.A(_0517_),
    .B(_0479_),
    .Y(_0518_));
 sky130_fd_sc_hd__and2b_1 _1035_ (.A_N(_0518_),
    .B(_0489_),
    .X(_0519_));
 sky130_fd_sc_hd__xnor2_1 _1036_ (.A(_0516_),
    .B(_0519_),
    .Y(\M0.FPM10.d ));
 sky130_fd_sc_hd__o21ba_1 _1037_ (.A1(_0275_),
    .A2(_0437_),
    .B1_N(_0485_),
    .X(_0520_));
 sky130_fd_sc_hd__xnor2_1 _1038_ (.A(_0345_),
    .B(_0482_),
    .Y(_0521_));
 sky130_fd_sc_hd__xnor2_1 _1039_ (.A(_0520_),
    .B(_0521_),
    .Y(\M0.FPM9.d ));
 sky130_fd_sc_hd__or3_1 _1040_ (.A(_0401_),
    .B(_0402_),
    .C(_0403_),
    .X(_0522_));
 sky130_fd_sc_hd__xor2_1 _1041_ (.A(_0397_),
    .B(_0400_),
    .X(_0523_));
 sky130_fd_sc_hd__xnor2_1 _1042_ (.A(_0522_),
    .B(_0523_),
    .Y(\M0.FPM4.d ));
 sky130_fd_sc_hd__nand2_1 _1043_ (.A(_0433_),
    .B(_0434_),
    .Y(_0524_));
 sky130_fd_sc_hd__xnor2_1 _1044_ (.A(_0132_),
    .B(_0436_),
    .Y(_0525_));
 sky130_fd_sc_hd__xnor2_1 _1045_ (.A(_0524_),
    .B(_0525_),
    .Y(\M0.FPM8.d ));
 sky130_fd_sc_hd__nand2_1 _1046_ (.A(_0372_),
    .B(_0392_),
    .Y(_0526_));
 sky130_fd_sc_hd__xnor2_1 _1047_ (.A(_0362_),
    .B(_0526_),
    .Y(\M0.FPM3.d ));
 sky130_fd_sc_hd__nand2_1 _1048_ (.A(_0176_),
    .B(_0234_),
    .Y(_0527_));
 sky130_fd_sc_hd__nand2_1 _1049_ (.A(_0174_),
    .B(_0236_),
    .Y(_0528_));
 sky130_fd_sc_hd__xor2_1 _1050_ (.A(_0527_),
    .B(_0528_),
    .X(\M0.FPM1.d ));
 sky130_fd_sc_hd__a21o_1 _1051_ (.A1(_0293_),
    .A2(_0363_),
    .B1(_0349_),
    .X(_0529_));
 sky130_fd_sc_hd__or3_1 _1052_ (.A(_0172_),
    .B(_0293_),
    .C(_0237_),
    .X(_0530_));
 sky130_fd_sc_hd__a21bo_1 _1053_ (.A1(_0172_),
    .A2(_0529_),
    .B1_N(_0530_),
    .X(_0531_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(_0365_),
    .A1(_0384_),
    .S(_0371_),
    .X(_0532_));
 sky130_fd_sc_hd__a21oi_1 _1055_ (.A1(_0234_),
    .A2(_0531_),
    .B1(_0532_),
    .Y(\M0.FPM2.d ));
 sky130_fd_sc_hd__a21oi_1 _1056_ (.A1(_0411_),
    .A2(_0423_),
    .B1(_0424_),
    .Y(_0533_));
 sky130_fd_sc_hd__and2b_1 _1057_ (.A_N(_0432_),
    .B(_0434_),
    .X(_0534_));
 sky130_fd_sc_hd__xnor2_1 _1058_ (.A(_0533_),
    .B(_0534_),
    .Y(\M0.FPM7.d ));
 sky130_fd_sc_hd__a21o_1 _1059_ (.A1(_0412_),
    .A2(_0419_),
    .B1(_0422_),
    .X(_0535_));
 sky130_fd_sc_hd__a21oi_1 _1060_ (.A1(_0423_),
    .A2(_0535_),
    .B1(_0411_),
    .Y(_0536_));
 sky130_fd_sc_hd__and3_1 _1061_ (.A(_0411_),
    .B(_0423_),
    .C(_0535_),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_1 _1062_ (.A(_0536_),
    .B(_0537_),
    .Y(\M0.FPM6.d ));
 sky130_fd_sc_hd__xor2_1 _1063_ (.A(_0383_),
    .B(_0408_),
    .X(_0538_));
 sky130_fd_sc_hd__xnor2_1 _1064_ (.A(_0405_),
    .B(_0538_),
    .Y(\M0.FPM5.d ));
 sky130_fd_sc_hd__buf_8 _1065_ (.A(net19),
    .X(_0539_));
 sky130_fd_sc_hd__clkbuf_16 _1066_ (.A(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__inv_2 _1067_ (.A(_0540_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _1068_ (.A(_0540_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1069_ (.A(_0540_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1070_ (.A(_0540_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1071_ (.A(_0540_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1072_ (.A(_0540_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1073_ (.A(_0540_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1074_ (.A(_0540_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1075_ (.A(_0540_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1076_ (.A(_0540_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1077_ (.A(_0540_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1078_ (.A(_0540_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1079_ (.A(_0540_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1080_ (.A(_0540_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1081_ (.A(_0540_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1082_ (.A(_0540_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1083_ (.A(_0540_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1084_ (.A(_0540_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1085_ (.A(_0540_),
    .Y(_0018_));
 sky130_fd_sc_hd__clkbuf_16 _1086_ (.A(_0539_),
    .X(_0541_));
 sky130_fd_sc_hd__inv_2 _1087_ (.A(_0541_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1088_ (.A(_0541_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1089_ (.A(_0541_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1090_ (.A(_0541_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1091_ (.A(_0541_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1092_ (.A(_0541_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1093_ (.A(_0541_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1094_ (.A(_0541_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1095_ (.A(_0541_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1096_ (.A(_0541_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1097_ (.A(_0541_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1098_ (.A(_0541_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1099_ (.A(_0541_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1100_ (.A(_0541_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1101_ (.A(_0541_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1102_ (.A(_0541_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1103_ (.A(_0541_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1104_ (.A(_0541_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1105_ (.A(_0541_),
    .Y(_0037_));
 sky130_fd_sc_hd__clkbuf_16 _1106_ (.A(_0539_),
    .X(_0542_));
 sky130_fd_sc_hd__inv_2 _1107_ (.A(_0542_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1108_ (.A(_0542_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1109_ (.A(_0542_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1110_ (.A(_0542_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1111_ (.A(_0542_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1112_ (.A(_0542_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1113_ (.A(_0542_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1114_ (.A(_0542_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1115_ (.A(_0542_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1116_ (.A(_0542_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1117_ (.A(_0542_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1118_ (.A(_0542_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1119_ (.A(_0542_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1120_ (.A(_0542_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1121_ (.A(_0542_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1122_ (.A(_0542_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1123_ (.A(_0542_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1124_ (.A(_0542_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1125_ (.A(_0542_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1126_ (.A(_0539_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1127_ (.A(_0539_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1128_ (.A(_0539_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1129_ (.A(_0539_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1130_ (.A(_0539_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1131_ (.A(_0539_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1132_ (.A(_0539_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1133_ (.A(_0539_),
    .Y(_0064_));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(net17),
    .D(\M0.FPM15.d ),
    .RESET_B(_0000_),
    .Q(\M0.FPM15.q ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(net17),
    .D(\M0.FPM14.d ),
    .RESET_B(_0001_),
    .Q(\M0.FPM14.q ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(net17),
    .D(\M0.FPM13.d ),
    .RESET_B(_0002_),
    .Q(\M0.FPM13.q ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(net17),
    .D(\M0.FPM12.d ),
    .RESET_B(_0003_),
    .Q(\M0.FPM12.q ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(net17),
    .D(\M0.FPM11.d ),
    .RESET_B(_0004_),
    .Q(\M0.FPM11.q ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(net17),
    .D(\M0.FPM10.d ),
    .RESET_B(_0005_),
    .Q(\M0.FPM10.q ));
 sky130_fd_sc_hd__dfrtp_1 _1140_ (.CLK(net17),
    .D(\M0.FPM9.d ),
    .RESET_B(_0006_),
    .Q(\M0.FPM9.q ));
 sky130_fd_sc_hd__dfrtp_1 _1141_ (.CLK(net17),
    .D(\M0.FPM8.d ),
    .RESET_B(_0007_),
    .Q(\M0.FPM8.q ));
 sky130_fd_sc_hd__dfrtp_1 _1142_ (.CLK(net17),
    .D(\M0.FPM7.d ),
    .RESET_B(_0008_),
    .Q(\M0.FPM7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(net17),
    .D(\M0.FPM6.d ),
    .RESET_B(_0009_),
    .Q(\M0.FPM6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(net17),
    .D(\M0.FPM5.d ),
    .RESET_B(_0010_),
    .Q(\M0.FPM5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(net17),
    .D(\M0.FPM4.d ),
    .RESET_B(_0011_),
    .Q(\M0.FPM4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1146_ (.CLK(net17),
    .D(\M0.FPM3.d ),
    .RESET_B(_0012_),
    .Q(\M0.FPM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1147_ (.CLK(net17),
    .D(\M0.FPM2.d ),
    .RESET_B(_0013_),
    .Q(\M0.FPM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1148_ (.CLK(net17),
    .D(\M0.FPM1.d ),
    .RESET_B(_0014_),
    .Q(\M0.FPM1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1149_ (.CLK(net17),
    .D(\M0.FPM0.d ),
    .RESET_B(_0015_),
    .Q(\M0.FPM0.q ));
 sky130_fd_sc_hd__dfrtp_4 _1150_ (.CLK(net17),
    .D(\M0.FBM7.d ),
    .RESET_B(_0016_),
    .Q(\M0.FBM7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1151_ (.CLK(net17),
    .D(\M0.FBM6.d ),
    .RESET_B(_0017_),
    .Q(\M0.FBM6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1152_ (.CLK(net17),
    .D(\M0.FBM5.d ),
    .RESET_B(_0018_),
    .Q(\M0.FBM5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1153_ (.CLK(net17),
    .D(\M0.FBM4.d ),
    .RESET_B(_0019_),
    .Q(\M0.FBM4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1154_ (.CLK(net17),
    .D(\M0.FBM3.d ),
    .RESET_B(_0020_),
    .Q(\M0.FBM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1155_ (.CLK(net17),
    .D(\M0.FBM2.d ),
    .RESET_B(_0021_),
    .Q(\M0.FBM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1156_ (.CLK(net17),
    .D(\M0.FBM1.d ),
    .RESET_B(_0022_),
    .Q(\M0.FBM1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1157_ (.CLK(net17),
    .D(\M0.FBM0.d ),
    .RESET_B(_0023_),
    .Q(\M0.FBM0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1158_ (.CLK(net17),
    .D(\M0.FAM7.d ),
    .RESET_B(_0024_),
    .Q(\M0.FAM7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1159_ (.CLK(net17),
    .D(\M0.FAM6.d ),
    .RESET_B(_0025_),
    .Q(\M0.FAM6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1160_ (.CLK(net17),
    .D(\M0.FAM5.d ),
    .RESET_B(_0026_),
    .Q(\M0.FAM5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1161_ (.CLK(net17),
    .D(\M0.FAM4.d ),
    .RESET_B(_0027_),
    .Q(\M0.FAM4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1162_ (.CLK(net17),
    .D(\M0.FAM3.d ),
    .RESET_B(_0028_),
    .Q(\M0.FAM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1163_ (.CLK(net17),
    .D(\M0.FAM2.d ),
    .RESET_B(_0029_),
    .Q(\M0.FAM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1164_ (.CLK(net17),
    .D(\M0.FAM1.d ),
    .RESET_B(_0030_),
    .Q(\M0.FAM1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1165_ (.CLK(net17),
    .D(\M0.FAM0.d ),
    .RESET_B(_0031_),
    .Q(\M0.FAM0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1166_ (.CLK(net17),
    .D(\FP0.d ),
    .RESET_B(_0032_),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _1167_ (.CLK(net17),
    .D(\FP1.d ),
    .RESET_B(_0033_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _1168_ (.CLK(net17),
    .D(\FP2.d ),
    .RESET_B(_0034_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _1169_ (.CLK(net17),
    .D(\FP3.d ),
    .RESET_B(_0035_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _1170_ (.CLK(net17),
    .D(\FP4.d ),
    .RESET_B(_0036_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _1171_ (.CLK(net17),
    .D(\FP5.d ),
    .RESET_B(_0037_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _1172_ (.CLK(net17),
    .D(\FP6.d ),
    .RESET_B(_0038_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _1173_ (.CLK(net17),
    .D(\FP7.d ),
    .RESET_B(_0039_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _1174_ (.CLK(net17),
    .D(\FP8.d ),
    .RESET_B(_0040_),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _1175_ (.CLK(net17),
    .D(\FP9.d ),
    .RESET_B(_0041_),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _1176_ (.CLK(net17),
    .D(\FP10.d ),
    .RESET_B(_0042_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _1177_ (.CLK(net17),
    .D(\FP11.d ),
    .RESET_B(_0043_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _1178_ (.CLK(net17),
    .D(\FP12.d ),
    .RESET_B(_0044_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _1179_ (.CLK(net17),
    .D(\FP13.d ),
    .RESET_B(_0045_),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _1180_ (.CLK(net17),
    .D(\FP14.d ),
    .RESET_B(_0046_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _1181_ (.CLK(net17),
    .D(\FP15.d ),
    .RESET_B(_0047_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _1182_ (.CLK(net17),
    .D(net1),
    .RESET_B(_0048_),
    .Q(\FA0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1183_ (.CLK(net17),
    .D(net2),
    .RESET_B(_0049_),
    .Q(\FA1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1184_ (.CLK(net17),
    .D(net3),
    .RESET_B(_0050_),
    .Q(\FA2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1185_ (.CLK(net17),
    .D(net4),
    .RESET_B(_0051_),
    .Q(\FA3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1186_ (.CLK(net17),
    .D(net5),
    .RESET_B(_0052_),
    .Q(\FA4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1187_ (.CLK(net17),
    .D(net6),
    .RESET_B(_0053_),
    .Q(\FA5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1188_ (.CLK(net17),
    .D(net7),
    .RESET_B(_0054_),
    .Q(\FA6.q ));
 sky130_fd_sc_hd__dfrtp_4 _1189_ (.CLK(net17),
    .D(net8),
    .RESET_B(_0055_),
    .Q(\FA7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1190_ (.CLK(net17),
    .D(net9),
    .RESET_B(_0056_),
    .Q(\FB0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1191_ (.CLK(net17),
    .D(net10),
    .RESET_B(_0057_),
    .Q(\FB1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1192_ (.CLK(net17),
    .D(net11),
    .RESET_B(_0058_),
    .Q(\FB2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1193_ (.CLK(net17),
    .D(net12),
    .RESET_B(_0059_),
    .Q(\FB3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1194_ (.CLK(net17),
    .D(net13),
    .RESET_B(_0060_),
    .Q(\FB4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1195_ (.CLK(net17),
    .D(net14),
    .RESET_B(_0061_),
    .Q(\FB5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1196_ (.CLK(net17),
    .D(net15),
    .RESET_B(_0062_),
    .Q(\FB6.q ));
 sky130_fd_sc_hd__dfrtp_4 _1197_ (.CLK(net17),
    .D(net16),
    .RESET_B(_0063_),
    .Q(\FB7.q ));
 sky130_fd_sc_hd__dfrtp_4 _1198_ (.CLK(net17),
    .D(net18),
    .RESET_B(_0064_),
    .Q(\FC.q ));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(clk),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(control),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(rst),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap36 (.A(_0300_),
    .X(net36));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(p[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(p[10]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(p[11]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(p[12]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(p[13]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(p[14]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(p[15]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(p[1]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(p[2]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(p[3]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(p[4]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(p[5]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(p[6]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(p[7]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(p[8]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(p[9]));
endmodule

