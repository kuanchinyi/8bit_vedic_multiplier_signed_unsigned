magic
tech sky130A
magscale 1 2
timestamp 1729948589
<< obsli1 >>
rect 1104 2159 35236 36465
<< obsm1 >>
rect 934 2128 35296 36496
<< metal2 >>
rect 9034 0 9090 800
rect 27250 0 27306 800
<< obsm2 >>
rect 938 856 35242 36825
rect 938 800 8978 856
rect 9146 800 27194 856
rect 27362 800 35242 856
<< metal3 >>
rect 0 36728 800 36848
rect 35600 35640 36400 35760
rect 0 34552 800 34672
rect 35600 33464 36400 33584
rect 0 32376 800 32496
rect 35600 31288 36400 31408
rect 0 30200 800 30320
rect 35600 29112 36400 29232
rect 0 28024 800 28144
rect 35600 26936 36400 27056
rect 0 25848 800 25968
rect 35600 24760 36400 24880
rect 0 23672 800 23792
rect 35600 22584 36400 22704
rect 0 21496 800 21616
rect 35600 20408 36400 20528
rect 0 19320 800 19440
rect 35600 18232 36400 18352
rect 0 17144 800 17264
rect 35600 16056 36400 16176
rect 0 14968 800 15088
rect 35600 13880 36400 14000
rect 0 12792 800 12912
rect 35600 11704 36400 11824
rect 0 10616 800 10736
rect 35600 9528 36400 9648
rect 0 8440 800 8560
rect 35600 7352 36400 7472
rect 0 6264 800 6384
rect 35600 5176 36400 5296
rect 0 4088 800 4208
rect 35600 3000 36400 3120
rect 0 1912 800 2032
<< obsm3 >>
rect 880 36648 35600 36821
rect 798 35840 35600 36648
rect 798 35560 35520 35840
rect 798 34752 35600 35560
rect 880 34472 35600 34752
rect 798 33664 35600 34472
rect 798 33384 35520 33664
rect 798 32576 35600 33384
rect 880 32296 35600 32576
rect 798 31488 35600 32296
rect 798 31208 35520 31488
rect 798 30400 35600 31208
rect 880 30120 35600 30400
rect 798 29312 35600 30120
rect 798 29032 35520 29312
rect 798 28224 35600 29032
rect 880 27944 35600 28224
rect 798 27136 35600 27944
rect 798 26856 35520 27136
rect 798 26048 35600 26856
rect 880 25768 35600 26048
rect 798 24960 35600 25768
rect 798 24680 35520 24960
rect 798 23872 35600 24680
rect 880 23592 35600 23872
rect 798 22784 35600 23592
rect 798 22504 35520 22784
rect 798 21696 35600 22504
rect 880 21416 35600 21696
rect 798 20608 35600 21416
rect 798 20328 35520 20608
rect 798 19520 35600 20328
rect 880 19240 35600 19520
rect 798 18432 35600 19240
rect 798 18152 35520 18432
rect 798 17344 35600 18152
rect 880 17064 35600 17344
rect 798 16256 35600 17064
rect 798 15976 35520 16256
rect 798 15168 35600 15976
rect 880 14888 35600 15168
rect 798 14080 35600 14888
rect 798 13800 35520 14080
rect 798 12992 35600 13800
rect 880 12712 35600 12992
rect 798 11904 35600 12712
rect 798 11624 35520 11904
rect 798 10816 35600 11624
rect 880 10536 35600 10816
rect 798 9728 35600 10536
rect 798 9448 35520 9728
rect 798 8640 35600 9448
rect 880 8360 35600 8640
rect 798 7552 35600 8360
rect 798 7272 35520 7552
rect 798 6464 35600 7272
rect 880 6184 35600 6464
rect 798 5376 35600 6184
rect 798 5096 35520 5376
rect 798 4288 35600 5096
rect 880 4008 35600 4288
rect 798 3200 35600 4008
rect 798 2920 35520 3200
rect 798 2112 35600 2920
rect 880 1939 35600 2112
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< obsm4 >>
rect 5395 15131 5461 20773
<< labels >>
rlabel metal3 s 0 4088 800 4208 6 a[0]
port 1 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 a[1]
port 2 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 a[2]
port 3 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 a[3]
port 4 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 a[4]
port 5 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 a[5]
port 6 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 a[6]
port 7 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 a[7]
port 8 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 b[0]
port 9 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 b[1]
port 10 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 b[2]
port 11 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 b[3]
port 12 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 b[4]
port 13 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 b[5]
port 14 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 b[6]
port 15 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 b[7]
port 16 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 clk
port 17 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 control
port 18 nsew signal input
rlabel metal3 s 35600 3000 36400 3120 6 p[0]
port 19 nsew signal output
rlabel metal3 s 35600 24760 36400 24880 6 p[10]
port 20 nsew signal output
rlabel metal3 s 35600 26936 36400 27056 6 p[11]
port 21 nsew signal output
rlabel metal3 s 35600 29112 36400 29232 6 p[12]
port 22 nsew signal output
rlabel metal3 s 35600 31288 36400 31408 6 p[13]
port 23 nsew signal output
rlabel metal3 s 35600 33464 36400 33584 6 p[14]
port 24 nsew signal output
rlabel metal3 s 35600 35640 36400 35760 6 p[15]
port 25 nsew signal output
rlabel metal3 s 35600 5176 36400 5296 6 p[1]
port 26 nsew signal output
rlabel metal3 s 35600 7352 36400 7472 6 p[2]
port 27 nsew signal output
rlabel metal3 s 35600 9528 36400 9648 6 p[3]
port 28 nsew signal output
rlabel metal3 s 35600 11704 36400 11824 6 p[4]
port 29 nsew signal output
rlabel metal3 s 35600 13880 36400 14000 6 p[5]
port 30 nsew signal output
rlabel metal3 s 35600 16056 36400 16176 6 p[6]
port 31 nsew signal output
rlabel metal3 s 35600 18232 36400 18352 6 p[7]
port 32 nsew signal output
rlabel metal3 s 35600 20408 36400 20528 6 p[8]
port 33 nsew signal output
rlabel metal3 s 35600 22584 36400 22704 6 p[9]
port 34 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 rst
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 37 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36400 38800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2806810
string GDS_FILE /home/cykuan/chinyi2/8bit_vedic_multiplier_signed_unsigned/openlane/vmsu_8bit_top/runs/24_10_26_21_14/results/signoff/vmsu_8bit_top.magic.gds
string GDS_START 780886
<< end >>

