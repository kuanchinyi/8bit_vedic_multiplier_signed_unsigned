// This is the unpowered netlist.
module vmsu_8bit_top (clk,
    control,
    rst,
    a,
    b,
    p);
 input clk;
 input control;
 input rst;
 input [7:0] a;
 input [7:0] b;
 output [15:0] p;

 wire \FA0.q ;
 wire \FA1.q ;
 wire \FA2.q ;
 wire \FA3.q ;
 wire \FA4.q ;
 wire \FA5.q ;
 wire \FA6.q ;
 wire \FA7.q ;
 wire \FB0.q ;
 wire \FB1.q ;
 wire \FB2.q ;
 wire \FB3.q ;
 wire \FB4.q ;
 wire \FB5.q ;
 wire \FB6.q ;
 wire \FB7.q ;
 wire \FC.q ;
 wire \FP0.d ;
 wire \FP1.d ;
 wire \FP10.d ;
 wire \FP11.d ;
 wire \FP12.d ;
 wire \FP13.d ;
 wire \FP14.d ;
 wire \FP15.d ;
 wire \FP2.d ;
 wire \FP3.d ;
 wire \FP4.d ;
 wire \FP5.d ;
 wire \FP6.d ;
 wire \FP7.d ;
 wire \FP8.d ;
 wire \FP9.d ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__415__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__429__B1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__439__B1 (.DIODE(\FP0.d ));
 sky130_fd_sc_hd__diode_2 ANTENNA__442__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__465__A1 (.DIODE(_395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__492__A1 (.DIODE(_395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__528__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__549__B (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__562__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__585__C (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__585__D_N (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__586__A2_N (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__586__B1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__606__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__620__B (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__622__A2 (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__622__B1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__A3 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__640__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__658__A2_N (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__658__B1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__659__A2 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__679__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__687__A2 (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__687__B1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__699__B (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__710__A1 (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__714__C1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__726__C (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__726__D_N (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__727__A2_N (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__727__B1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__741__A (.DIODE(_396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__742__B (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__744__C_N (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__760__A1 (.DIODE(_395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__761__B (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__762__B (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__763__A1 (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__782__A2 (.DIODE(_136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__782__C1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__787__B1 (.DIODE(_172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__789__A1 (.DIODE(_395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__791__A1 (.DIODE(_395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__807__A (.DIODE(\FP0.d ));
 sky130_fd_sc_hd__diode_2 ANTENNA__807__B (.DIODE(_395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__810__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__811__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__812__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__813__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__814__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__815__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__816__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__817__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__818__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__819__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__820__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__821__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__822__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__823__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__824__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__825__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__826__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__827__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__828__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__829__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__830__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__831__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__832__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__833__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__834__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__835__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__836__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__837__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__838__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__839__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__840__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__841__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__842__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__842__D (.DIODE(\FP0.d ));
 sky130_fd_sc_hd__diode_2 ANTENNA__843__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__844__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__845__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__846__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__847__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__848__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__849__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__850__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__851__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__852__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__853__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__854__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__855__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__856__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__857__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__858__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__859__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__860__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__861__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__862__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__863__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__864__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__865__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__866__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__867__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__868__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__869__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__870__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__871__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__872__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__873__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__874__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_367 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__inv_2 _413_ (.A(\FA0.q ),
    .Y(_383_));
 sky130_fd_sc_hd__inv_2 _414_ (.A(\FB0.q ),
    .Y(_384_));
 sky130_fd_sc_hd__inv_2 _415_ (.A(net19),
    .Y(_000_));
 sky130_fd_sc_hd__nand2_1 _416_ (.A(\FA0.q ),
    .B(\FB0.q ),
    .Y(_385_));
 sky130_fd_sc_hd__inv_2 _417_ (.A(_385_),
    .Y(\FP0.d ));
 sky130_fd_sc_hd__and2_4 _418_ (.A(\FC.q ),
    .B(\FB7.q ),
    .X(_386_));
 sky130_fd_sc_hd__and3_4 _419_ (.A(\FC.q ),
    .B(\FB7.q ),
    .C(\FB0.q ),
    .X(_387_));
 sky130_fd_sc_hd__xor2_4 _420_ (.A(\FB1.q ),
    .B(_387_),
    .X(_388_));
 sky130_fd_sc_hd__xnor2_4 _421_ (.A(\FB1.q ),
    .B(_387_),
    .Y(_389_));
 sky130_fd_sc_hd__and2_4 _422_ (.A(\FA7.q ),
    .B(\FC.q ),
    .X(_390_));
 sky130_fd_sc_hd__and3_2 _423_ (.A(\FA7.q ),
    .B(\FC.q ),
    .C(\FA0.q ),
    .X(_391_));
 sky130_fd_sc_hd__xor2_2 _424_ (.A(\FA1.q ),
    .B(_391_),
    .X(_392_));
 sky130_fd_sc_hd__xnor2_4 _425_ (.A(\FA1.q ),
    .B(_391_),
    .Y(_393_));
 sky130_fd_sc_hd__o22a_1 _426_ (.A1(_383_),
    .A2(_389_),
    .B1(_393_),
    .B2(_384_),
    .X(_394_));
 sky130_fd_sc_hd__xor2_4 _427_ (.A(_386_),
    .B(_390_),
    .X(_395_));
 sky130_fd_sc_hd__xnor2_4 _428_ (.A(_386_),
    .B(_390_),
    .Y(_396_));
 sky130_fd_sc_hd__a21o_1 _429_ (.A1(_385_),
    .A2(_394_),
    .B1(_396_),
    .X(_397_));
 sky130_fd_sc_hd__o211a_2 _430_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .B1(\FC.q ),
    .C1(\FB7.q ),
    .X(_398_));
 sky130_fd_sc_hd__xor2_2 _431_ (.A(\FB2.q ),
    .B(_398_),
    .X(_399_));
 sky130_fd_sc_hd__xnor2_4 _432_ (.A(\FB2.q ),
    .B(_398_),
    .Y(_400_));
 sky130_fd_sc_hd__nand2_1 _433_ (.A(\FA0.q ),
    .B(_399_),
    .Y(_401_));
 sky130_fd_sc_hd__o211a_4 _434_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .B1(\FA7.q ),
    .C1(\FC.q ),
    .X(_402_));
 sky130_fd_sc_hd__xor2_4 _435_ (.A(\FA2.q ),
    .B(_402_),
    .X(_403_));
 sky130_fd_sc_hd__xnor2_4 _436_ (.A(\FA2.q ),
    .B(_402_),
    .Y(_404_));
 sky130_fd_sc_hd__nand2_1 _437_ (.A(\FB0.q ),
    .B(_403_),
    .Y(_405_));
 sky130_fd_sc_hd__nand2_1 _438_ (.A(_401_),
    .B(_405_),
    .Y(_406_));
 sky130_fd_sc_hd__a2111o_1 _439_ (.A1(_401_),
    .A2(_405_),
    .B1(\FP0.d ),
    .C1(_389_),
    .D1(_393_),
    .X(_407_));
 sky130_fd_sc_hd__a31o_1 _440_ (.A1(_385_),
    .A2(_388_),
    .A3(_392_),
    .B1(_406_),
    .X(_408_));
 sky130_fd_sc_hd__nand2_1 _441_ (.A(_407_),
    .B(_408_),
    .Y(_409_));
 sky130_fd_sc_hd__o21a_1 _442_ (.A1(_396_),
    .A2(_409_),
    .B1(_397_),
    .X(_410_));
 sky130_fd_sc_hd__o311a_4 _443_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .A3(\FB2.q ),
    .B1(\FB7.q ),
    .C1(\FC.q ),
    .X(_411_));
 sky130_fd_sc_hd__xor2_4 _444_ (.A(\FB3.q ),
    .B(_411_),
    .X(_412_));
 sky130_fd_sc_hd__xnor2_4 _445_ (.A(\FB3.q ),
    .B(_411_),
    .Y(_033_));
 sky130_fd_sc_hd__or4_2 _446_ (.A(_383_),
    .B(_393_),
    .C(_400_),
    .D(_033_),
    .X(_034_));
 sky130_fd_sc_hd__a22o_1 _447_ (.A1(_392_),
    .A2(_399_),
    .B1(_412_),
    .B2(\FA0.q ),
    .X(_035_));
 sky130_fd_sc_hd__o311a_4 _448_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .A3(\FA2.q ),
    .B1(\FC.q ),
    .C1(\FA7.q ),
    .X(_036_));
 sky130_fd_sc_hd__xor2_4 _449_ (.A(\FA3.q ),
    .B(_036_),
    .X(_037_));
 sky130_fd_sc_hd__xnor2_4 _450_ (.A(\FA3.q ),
    .B(_036_),
    .Y(_038_));
 sky130_fd_sc_hd__or4_2 _451_ (.A(_384_),
    .B(_389_),
    .C(_404_),
    .D(_038_),
    .X(_039_));
 sky130_fd_sc_hd__a22o_1 _452_ (.A1(_388_),
    .A2(_403_),
    .B1(_037_),
    .B2(\FB0.q ),
    .X(_040_));
 sky130_fd_sc_hd__nand4_2 _453_ (.A(_034_),
    .B(_035_),
    .C(_039_),
    .D(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__a22o_1 _454_ (.A1(_034_),
    .A2(_035_),
    .B1(_039_),
    .B2(_040_),
    .X(_042_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(_401_),
    .B(_405_),
    .Y(_043_));
 sky130_fd_sc_hd__and3_1 _456_ (.A(_041_),
    .B(_042_),
    .C(_043_),
    .X(_044_));
 sky130_fd_sc_hd__a21o_1 _457_ (.A1(_041_),
    .A2(_042_),
    .B1(_043_),
    .X(_045_));
 sky130_fd_sc_hd__and2b_1 _458_ (.A_N(_044_),
    .B(_045_),
    .X(_046_));
 sky130_fd_sc_hd__and4_1 _459_ (.A(\FA0.q ),
    .B(\FB0.q ),
    .C(_388_),
    .D(_392_),
    .X(_047_));
 sky130_fd_sc_hd__inv_2 _460_ (.A(_047_),
    .Y(_048_));
 sky130_fd_sc_hd__nand2_1 _461_ (.A(_407_),
    .B(_048_),
    .Y(_049_));
 sky130_fd_sc_hd__and3b_1 _462_ (.A_N(_044_),
    .B(_045_),
    .C(_049_),
    .X(_050_));
 sky130_fd_sc_hd__nor2_1 _463_ (.A(_046_),
    .B(_049_),
    .Y(_051_));
 sky130_fd_sc_hd__nor2_1 _464_ (.A(_050_),
    .B(_051_),
    .Y(_052_));
 sky130_fd_sc_hd__a21bo_1 _465_ (.A1(_395_),
    .A2(_052_),
    .B1_N(_410_),
    .X(_053_));
 sky130_fd_sc_hd__or4_4 _466_ (.A(\FB0.q ),
    .B(\FB1.q ),
    .C(\FB2.q ),
    .D(\FB3.q ),
    .X(_054_));
 sky130_fd_sc_hd__nand2_2 _467_ (.A(_386_),
    .B(_054_),
    .Y(_055_));
 sky130_fd_sc_hd__xor2_4 _468_ (.A(\FB4.q ),
    .B(_055_),
    .X(_056_));
 sky130_fd_sc_hd__inv_2 _469_ (.A(_056_),
    .Y(_057_));
 sky130_fd_sc_hd__nor2_2 _470_ (.A(_383_),
    .B(_056_),
    .Y(_058_));
 sky130_fd_sc_hd__or4_4 _471_ (.A(\FA0.q ),
    .B(\FA1.q ),
    .C(\FA2.q ),
    .D(\FA3.q ),
    .X(_059_));
 sky130_fd_sc_hd__nand2_2 _472_ (.A(_390_),
    .B(_059_),
    .Y(_060_));
 sky130_fd_sc_hd__xor2_4 _473_ (.A(\FA4.q ),
    .B(_060_),
    .X(_061_));
 sky130_fd_sc_hd__nor2_1 _474_ (.A(_384_),
    .B(_061_),
    .Y(_062_));
 sky130_fd_sc_hd__nand2_2 _475_ (.A(_058_),
    .B(_062_),
    .Y(_063_));
 sky130_fd_sc_hd__or2_1 _476_ (.A(_058_),
    .B(_062_),
    .X(_064_));
 sky130_fd_sc_hd__nand2_1 _477_ (.A(_063_),
    .B(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__nor2_1 _478_ (.A(_400_),
    .B(_404_),
    .Y(_066_));
 sky130_fd_sc_hd__or3b_1 _479_ (.A(_393_),
    .B(_033_),
    .C_N(_401_),
    .X(_067_));
 sky130_fd_sc_hd__or3b_1 _480_ (.A(_389_),
    .B(_038_),
    .C_N(_405_),
    .X(_068_));
 sky130_fd_sc_hd__and2_1 _481_ (.A(_067_),
    .B(_068_),
    .X(_069_));
 sky130_fd_sc_hd__xor2_1 _482_ (.A(_067_),
    .B(_068_),
    .X(_070_));
 sky130_fd_sc_hd__a21boi_1 _483_ (.A1(_042_),
    .A2(_043_),
    .B1_N(_041_),
    .Y(_071_));
 sky130_fd_sc_hd__xnor2_2 _484_ (.A(_070_),
    .B(_071_),
    .Y(_072_));
 sky130_fd_sc_hd__xor2_1 _485_ (.A(_050_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__and2_1 _486_ (.A(_066_),
    .B(_073_),
    .X(_074_));
 sky130_fd_sc_hd__nor2_1 _487_ (.A(_066_),
    .B(_073_),
    .Y(_075_));
 sky130_fd_sc_hd__or2_1 _488_ (.A(_074_),
    .B(_075_),
    .X(_076_));
 sky130_fd_sc_hd__nor2_1 _489_ (.A(_065_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__and2_1 _490_ (.A(_065_),
    .B(_076_),
    .X(_078_));
 sky130_fd_sc_hd__nor2_1 _491_ (.A(_077_),
    .B(_078_),
    .Y(_079_));
 sky130_fd_sc_hd__a21oi_1 _492_ (.A1(_395_),
    .A2(_079_),
    .B1(_053_),
    .Y(_080_));
 sky130_fd_sc_hd__or4_1 _493_ (.A(_400_),
    .B(_404_),
    .C(_033_),
    .D(_038_),
    .X(_081_));
 sky130_fd_sc_hd__a22o_1 _494_ (.A1(_403_),
    .A2(_412_),
    .B1(_037_),
    .B2(_399_),
    .X(_082_));
 sky130_fd_sc_hd__nand2_1 _495_ (.A(_081_),
    .B(_082_),
    .Y(_083_));
 sky130_fd_sc_hd__xnor2_1 _496_ (.A(_034_),
    .B(_039_),
    .Y(_084_));
 sky130_fd_sc_hd__o21a_1 _497_ (.A1(_067_),
    .A2(_068_),
    .B1(_041_),
    .X(_085_));
 sky130_fd_sc_hd__o21ai_2 _498_ (.A1(_069_),
    .A2(_085_),
    .B1(_084_),
    .Y(_086_));
 sky130_fd_sc_hd__nand3_1 _499_ (.A(_050_),
    .B(_072_),
    .C(_086_),
    .Y(_087_));
 sky130_fd_sc_hd__a21o_1 _500_ (.A1(_050_),
    .A2(_072_),
    .B1(_086_),
    .X(_088_));
 sky130_fd_sc_hd__nand3b_2 _501_ (.A_N(_083_),
    .B(_087_),
    .C(_088_),
    .Y(_089_));
 sky130_fd_sc_hd__a21bo_1 _502_ (.A1(_087_),
    .A2(_088_),
    .B1_N(_083_),
    .X(_090_));
 sky130_fd_sc_hd__nand2_1 _503_ (.A(_089_),
    .B(_090_),
    .Y(_091_));
 sky130_fd_sc_hd__nand3_1 _504_ (.A(_074_),
    .B(_089_),
    .C(_090_),
    .Y(_092_));
 sky130_fd_sc_hd__a21o_1 _505_ (.A1(_089_),
    .A2(_090_),
    .B1(_074_),
    .X(_093_));
 sky130_fd_sc_hd__o21ai_4 _506_ (.A1(\FB4.q ),
    .A2(_054_),
    .B1(_386_),
    .Y(_094_));
 sky130_fd_sc_hd__xnor2_1 _507_ (.A(\FB5.q ),
    .B(_094_),
    .Y(_095_));
 sky130_fd_sc_hd__xor2_4 _508_ (.A(\FB5.q ),
    .B(_094_),
    .X(_096_));
 sky130_fd_sc_hd__or4_1 _509_ (.A(_383_),
    .B(_393_),
    .C(_056_),
    .D(_096_),
    .X(_097_));
 sky130_fd_sc_hd__a2bb2o_1 _510_ (.A1_N(_393_),
    .A2_N(_056_),
    .B1(_095_),
    .B2(\FA0.q ),
    .X(_098_));
 sky130_fd_sc_hd__and2_1 _511_ (.A(_097_),
    .B(_098_),
    .X(_099_));
 sky130_fd_sc_hd__o21ai_4 _512_ (.A1(\FA4.q ),
    .A2(_059_),
    .B1(_390_),
    .Y(_100_));
 sky130_fd_sc_hd__xnor2_1 _513_ (.A(\FA5.q ),
    .B(_100_),
    .Y(_101_));
 sky130_fd_sc_hd__xor2_4 _514_ (.A(\FA5.q ),
    .B(_100_),
    .X(_102_));
 sky130_fd_sc_hd__or4_1 _515_ (.A(_384_),
    .B(_389_),
    .C(_061_),
    .D(_102_),
    .X(_103_));
 sky130_fd_sc_hd__a2bb2o_1 _516_ (.A1_N(_389_),
    .A2_N(_061_),
    .B1(_101_),
    .B2(\FB0.q ),
    .X(_104_));
 sky130_fd_sc_hd__and2_1 _517_ (.A(_103_),
    .B(_104_),
    .X(_105_));
 sky130_fd_sc_hd__nand2_1 _518_ (.A(_099_),
    .B(_105_),
    .Y(_106_));
 sky130_fd_sc_hd__nor2_1 _519_ (.A(_099_),
    .B(_105_),
    .Y(_107_));
 sky130_fd_sc_hd__inv_2 _520_ (.A(_107_),
    .Y(_108_));
 sky130_fd_sc_hd__nand2_1 _521_ (.A(_106_),
    .B(_108_),
    .Y(_109_));
 sky130_fd_sc_hd__xnor2_1 _522_ (.A(_063_),
    .B(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__xor2_1 _523_ (.A(_063_),
    .B(_109_),
    .X(_111_));
 sky130_fd_sc_hd__a21o_1 _524_ (.A1(_092_),
    .A2(_093_),
    .B1(_111_),
    .X(_112_));
 sky130_fd_sc_hd__nand3_1 _525_ (.A(_092_),
    .B(_093_),
    .C(_111_),
    .Y(_113_));
 sky130_fd_sc_hd__nand2_1 _526_ (.A(_112_),
    .B(_113_),
    .Y(_114_));
 sky130_fd_sc_hd__xor2_1 _527_ (.A(_077_),
    .B(_114_),
    .X(_115_));
 sky130_fd_sc_hd__o21ai_1 _528_ (.A1(_396_),
    .A2(_115_),
    .B1(_080_),
    .Y(_116_));
 sky130_fd_sc_hd__a2111o_1 _529_ (.A1(_091_),
    .A2(_110_),
    .B1(_065_),
    .C1(_074_),
    .D1(_075_),
    .X(_117_));
 sky130_fd_sc_hd__nand2_1 _530_ (.A(_113_),
    .B(_117_),
    .Y(_118_));
 sky130_fd_sc_hd__nand3_1 _531_ (.A(_046_),
    .B(_047_),
    .C(_086_),
    .Y(_119_));
 sky130_fd_sc_hd__a211oi_1 _532_ (.A1(_407_),
    .A2(_066_),
    .B1(_038_),
    .C1(_033_),
    .Y(_120_));
 sky130_fd_sc_hd__o2bb2a_1 _533_ (.A1_N(_119_),
    .A2_N(_120_),
    .B1(_034_),
    .B2(_039_),
    .X(_121_));
 sky130_fd_sc_hd__a21bo_1 _534_ (.A1(_074_),
    .A2(_090_),
    .B1_N(_089_),
    .X(_122_));
 sky130_fd_sc_hd__xor2_1 _535_ (.A(_121_),
    .B(_122_),
    .X(_123_));
 sky130_fd_sc_hd__a21oi_1 _536_ (.A1(_063_),
    .A2(_106_),
    .B1(_107_),
    .Y(_124_));
 sky130_fd_sc_hd__o31a_2 _537_ (.A1(\FB5.q ),
    .A2(\FB4.q ),
    .A3(_054_),
    .B1(_386_),
    .X(_125_));
 sky130_fd_sc_hd__xnor2_4 _538_ (.A(\FB6.q ),
    .B(_125_),
    .Y(_126_));
 sky130_fd_sc_hd__or2_1 _539_ (.A(_383_),
    .B(_126_),
    .X(_127_));
 sky130_fd_sc_hd__or2_1 _540_ (.A(_404_),
    .B(_056_),
    .X(_128_));
 sky130_fd_sc_hd__o311a_1 _541_ (.A1(_393_),
    .A2(_058_),
    .A3(_096_),
    .B1(_127_),
    .C1(_128_),
    .X(_129_));
 sky130_fd_sc_hd__nor2_1 _542_ (.A(_127_),
    .B(_128_),
    .Y(_130_));
 sky130_fd_sc_hd__a2111o_1 _543_ (.A1(_127_),
    .A2(_128_),
    .B1(_393_),
    .C1(_058_),
    .D1(_096_),
    .X(_131_));
 sky130_fd_sc_hd__and2b_1 _544_ (.A_N(_129_),
    .B(_131_),
    .X(_132_));
 sky130_fd_sc_hd__inv_2 _545_ (.A(_132_),
    .Y(_133_));
 sky130_fd_sc_hd__or2_2 _546_ (.A(_400_),
    .B(_061_),
    .X(_134_));
 sky130_fd_sc_hd__o31a_2 _547_ (.A1(\FA5.q ),
    .A2(\FA4.q ),
    .A3(_059_),
    .B1(_390_),
    .X(_135_));
 sky130_fd_sc_hd__xnor2_4 _548_ (.A(\FA6.q ),
    .B(_135_),
    .Y(_136_));
 sky130_fd_sc_hd__or2_2 _549_ (.A(_384_),
    .B(_136_),
    .X(_137_));
 sky130_fd_sc_hd__o311a_1 _550_ (.A1(_389_),
    .A2(_062_),
    .A3(_102_),
    .B1(_134_),
    .C1(_137_),
    .X(_138_));
 sky130_fd_sc_hd__nor2_1 _551_ (.A(_134_),
    .B(_137_),
    .Y(_139_));
 sky130_fd_sc_hd__a2111o_1 _552_ (.A1(_134_),
    .A2(_137_),
    .B1(_389_),
    .C1(_062_),
    .D1(_102_),
    .X(_140_));
 sky130_fd_sc_hd__or3b_1 _553_ (.A(_138_),
    .B(_139_),
    .C_N(_140_),
    .X(_141_));
 sky130_fd_sc_hd__nor3_1 _554_ (.A(_130_),
    .B(_133_),
    .C(_141_),
    .Y(_142_));
 sky130_fd_sc_hd__o21ai_1 _555_ (.A1(_130_),
    .A2(_133_),
    .B1(_141_),
    .Y(_143_));
 sky130_fd_sc_hd__and2b_1 _556_ (.A_N(_142_),
    .B(_143_),
    .X(_144_));
 sky130_fd_sc_hd__xnor2_1 _557_ (.A(_124_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(_123_),
    .B(_145_),
    .Y(_146_));
 sky130_fd_sc_hd__or2_1 _559_ (.A(_123_),
    .B(_145_),
    .X(_147_));
 sky130_fd_sc_hd__and2_1 _560_ (.A(_146_),
    .B(_147_),
    .X(_148_));
 sky130_fd_sc_hd__xnor2_1 _561_ (.A(_118_),
    .B(_148_),
    .Y(_149_));
 sky130_fd_sc_hd__o21ba_1 _562_ (.A1(_396_),
    .A2(_149_),
    .B1_N(_116_),
    .X(_150_));
 sky130_fd_sc_hd__a22o_1 _563_ (.A1(_113_),
    .A2(_117_),
    .B1(_123_),
    .B2(_145_),
    .X(_151_));
 sky130_fd_sc_hd__or2_1 _564_ (.A(_089_),
    .B(_121_),
    .X(_152_));
 sky130_fd_sc_hd__o21a_1 _565_ (.A1(_124_),
    .A2(_142_),
    .B1(_143_),
    .X(_153_));
 sky130_fd_sc_hd__or4_2 _566_ (.A(\FB5.q ),
    .B(\FB4.q ),
    .C(\FB6.q ),
    .D(_054_),
    .X(_154_));
 sky130_fd_sc_hd__a21boi_4 _567_ (.A1(\FC.q ),
    .A2(_154_),
    .B1_N(\FB7.q ),
    .Y(_155_));
 sky130_fd_sc_hd__inv_2 _568_ (.A(_155_),
    .Y(_156_));
 sky130_fd_sc_hd__or4b_2 _569_ (.A(_383_),
    .B(_393_),
    .C(_126_),
    .D_N(_155_),
    .X(_157_));
 sky130_fd_sc_hd__a2bb2o_1 _570_ (.A1_N(_393_),
    .A2_N(_126_),
    .B1(_155_),
    .B2(\FA0.q ),
    .X(_158_));
 sky130_fd_sc_hd__or4_2 _571_ (.A(_404_),
    .B(_038_),
    .C(_056_),
    .D(_096_),
    .X(_159_));
 sky130_fd_sc_hd__a2bb2o_1 _572_ (.A1_N(_038_),
    .A2_N(_056_),
    .B1(_095_),
    .B2(_403_),
    .X(_160_));
 sky130_fd_sc_hd__nand4_1 _573_ (.A(_157_),
    .B(_158_),
    .C(_159_),
    .D(_160_),
    .Y(_161_));
 sky130_fd_sc_hd__a22o_1 _574_ (.A1(_157_),
    .A2(_158_),
    .B1(_159_),
    .B2(_160_),
    .X(_162_));
 sky130_fd_sc_hd__and3_1 _575_ (.A(_130_),
    .B(_161_),
    .C(_162_),
    .X(_163_));
 sky130_fd_sc_hd__a21oi_1 _576_ (.A1(_161_),
    .A2(_162_),
    .B1(_130_),
    .Y(_164_));
 sky130_fd_sc_hd__nor2_1 _577_ (.A(_163_),
    .B(_164_),
    .Y(_165_));
 sky130_fd_sc_hd__nand2_1 _578_ (.A(_097_),
    .B(_131_),
    .Y(_166_));
 sky130_fd_sc_hd__or3b_2 _579_ (.A(_163_),
    .B(_164_),
    .C_N(_166_),
    .X(_167_));
 sky130_fd_sc_hd__xnor2_2 _580_ (.A(_165_),
    .B(_166_),
    .Y(_168_));
 sky130_fd_sc_hd__or4_4 _581_ (.A(_400_),
    .B(_033_),
    .C(_061_),
    .D(_102_),
    .X(_169_));
 sky130_fd_sc_hd__a2bb2o_1 _582_ (.A1_N(_033_),
    .A2_N(_061_),
    .B1(_101_),
    .B2(_399_),
    .X(_170_));
 sky130_fd_sc_hd__or4_2 _583_ (.A(\FA5.q ),
    .B(\FA4.q ),
    .C(\FA6.q ),
    .D(_059_),
    .X(_171_));
 sky130_fd_sc_hd__a21boi_4 _584_ (.A1(\FC.q ),
    .A2(_171_),
    .B1_N(\FA7.q ),
    .Y(_172_));
 sky130_fd_sc_hd__or4b_4 _585_ (.A(_384_),
    .B(_389_),
    .C(_136_),
    .D_N(_172_),
    .X(_173_));
 sky130_fd_sc_hd__a2bb2o_1 _586_ (.A1_N(_389_),
    .A2_N(_136_),
    .B1(_172_),
    .B2(\FB0.q ),
    .X(_174_));
 sky130_fd_sc_hd__and4_1 _587_ (.A(_169_),
    .B(_170_),
    .C(_173_),
    .D(_174_),
    .X(_175_));
 sky130_fd_sc_hd__nand4_1 _588_ (.A(_169_),
    .B(_170_),
    .C(_173_),
    .D(_174_),
    .Y(_176_));
 sky130_fd_sc_hd__a22o_1 _589_ (.A1(_169_),
    .A2(_170_),
    .B1(_173_),
    .B2(_174_),
    .X(_177_));
 sky130_fd_sc_hd__nand3_1 _590_ (.A(_139_),
    .B(_176_),
    .C(_177_),
    .Y(_178_));
 sky130_fd_sc_hd__a21o_1 _591_ (.A1(_176_),
    .A2(_177_),
    .B1(_139_),
    .X(_179_));
 sky130_fd_sc_hd__nand2_1 _592_ (.A(_103_),
    .B(_140_),
    .Y(_180_));
 sky130_fd_sc_hd__and3_1 _593_ (.A(_178_),
    .B(_179_),
    .C(_180_),
    .X(_181_));
 sky130_fd_sc_hd__a21oi_1 _594_ (.A1(_178_),
    .A2(_179_),
    .B1(_180_),
    .Y(_182_));
 sky130_fd_sc_hd__or2_1 _595_ (.A(_181_),
    .B(_182_),
    .X(_183_));
 sky130_fd_sc_hd__nor2_1 _596_ (.A(_168_),
    .B(_183_),
    .Y(_184_));
 sky130_fd_sc_hd__nand2_1 _597_ (.A(_168_),
    .B(_183_),
    .Y(_185_));
 sky130_fd_sc_hd__xor2_1 _598_ (.A(_168_),
    .B(_183_),
    .X(_186_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(_153_),
    .B(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a31o_1 _600_ (.A1(_081_),
    .A2(_119_),
    .A3(_152_),
    .B1(_187_),
    .X(_188_));
 sky130_fd_sc_hd__inv_2 _601_ (.A(_188_),
    .Y(_189_));
 sky130_fd_sc_hd__and4_1 _602_ (.A(_081_),
    .B(_119_),
    .C(_152_),
    .D(_187_),
    .X(_190_));
 sky130_fd_sc_hd__a211o_1 _603_ (.A1(_147_),
    .A2(_151_),
    .B1(_189_),
    .C1(_190_),
    .X(_191_));
 sky130_fd_sc_hd__o211ai_1 _604_ (.A1(_189_),
    .A2(_190_),
    .B1(_147_),
    .C1(_151_),
    .Y(_192_));
 sky130_fd_sc_hd__nand2_1 _605_ (.A(_191_),
    .B(_192_),
    .Y(_193_));
 sky130_fd_sc_hd__o21a_1 _606_ (.A1(_396_),
    .A2(_193_),
    .B1(_150_),
    .X(_194_));
 sky130_fd_sc_hd__or2_1 _607_ (.A(_056_),
    .B(_061_),
    .X(_195_));
 sky130_fd_sc_hd__a31o_1 _608_ (.A1(_147_),
    .A2(_151_),
    .A3(_188_),
    .B1(_190_),
    .X(_196_));
 sky130_fd_sc_hd__o21ai_1 _609_ (.A1(_153_),
    .A2(_184_),
    .B1(_185_),
    .Y(_197_));
 sky130_fd_sc_hd__nor2_1 _610_ (.A(_404_),
    .B(_126_),
    .Y(_198_));
 sky130_fd_sc_hd__o211a_1 _611_ (.A1(_404_),
    .A2(_056_),
    .B1(_095_),
    .C1(_037_),
    .X(_199_));
 sky130_fd_sc_hd__and4_1 _612_ (.A(_392_),
    .B(_127_),
    .C(_155_),
    .D(_199_),
    .X(_200_));
 sky130_fd_sc_hd__a31o_1 _613_ (.A1(_392_),
    .A2(_127_),
    .A3(_155_),
    .B1(_199_),
    .X(_201_));
 sky130_fd_sc_hd__and2b_1 _614_ (.A_N(_200_),
    .B(_201_),
    .X(_202_));
 sky130_fd_sc_hd__a21bo_1 _615_ (.A1(_130_),
    .A2(_162_),
    .B1_N(_161_),
    .X(_203_));
 sky130_fd_sc_hd__xor2_2 _616_ (.A(_202_),
    .B(_203_),
    .X(_204_));
 sky130_fd_sc_hd__xnor2_2 _617_ (.A(_167_),
    .B(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__and2_1 _618_ (.A(_198_),
    .B(_205_),
    .X(_206_));
 sky130_fd_sc_hd__xnor2_2 _619_ (.A(_198_),
    .B(_205_),
    .Y(_207_));
 sky130_fd_sc_hd__nor2_1 _620_ (.A(_400_),
    .B(_136_),
    .Y(_208_));
 sky130_fd_sc_hd__nor2_1 _621_ (.A(_033_),
    .B(_102_),
    .Y(_209_));
 sky130_fd_sc_hd__o211a_1 _622_ (.A1(_384_),
    .A2(_136_),
    .B1(_172_),
    .C1(_388_),
    .X(_210_));
 sky130_fd_sc_hd__and3_1 _623_ (.A(_134_),
    .B(_209_),
    .C(_210_),
    .X(_211_));
 sky130_fd_sc_hd__a32oi_4 _624_ (.A1(_388_),
    .A2(_137_),
    .A3(_172_),
    .B1(_209_),
    .B2(_134_),
    .Y(_212_));
 sky130_fd_sc_hd__nor2_1 _625_ (.A(_211_),
    .B(_212_),
    .Y(_213_));
 sky130_fd_sc_hd__a21oi_1 _626_ (.A1(_139_),
    .A2(_177_),
    .B1(_175_),
    .Y(_214_));
 sky130_fd_sc_hd__xnor2_2 _627_ (.A(_213_),
    .B(_214_),
    .Y(_215_));
 sky130_fd_sc_hd__xor2_1 _628_ (.A(_181_),
    .B(_215_),
    .X(_216_));
 sky130_fd_sc_hd__and2_1 _629_ (.A(_208_),
    .B(_216_),
    .X(_217_));
 sky130_fd_sc_hd__xnor2_1 _630_ (.A(_208_),
    .B(_216_),
    .Y(_218_));
 sky130_fd_sc_hd__or2_1 _631_ (.A(_207_),
    .B(_218_),
    .X(_219_));
 sky130_fd_sc_hd__and2_1 _632_ (.A(_207_),
    .B(_218_),
    .X(_220_));
 sky130_fd_sc_hd__xnor2_1 _633_ (.A(_207_),
    .B(_218_),
    .Y(_221_));
 sky130_fd_sc_hd__xnor2_1 _634_ (.A(_197_),
    .B(_221_),
    .Y(_222_));
 sky130_fd_sc_hd__a311o_1 _635_ (.A1(_147_),
    .A2(_151_),
    .A3(_188_),
    .B1(_190_),
    .C1(_222_),
    .X(_223_));
 sky130_fd_sc_hd__xnor2_1 _636_ (.A(_196_),
    .B(_222_),
    .Y(_224_));
 sky130_fd_sc_hd__nor2_1 _637_ (.A(_195_),
    .B(_224_),
    .Y(_225_));
 sky130_fd_sc_hd__and2_1 _638_ (.A(_195_),
    .B(_224_),
    .X(_226_));
 sky130_fd_sc_hd__or2_1 _639_ (.A(_225_),
    .B(_226_),
    .X(_227_));
 sky130_fd_sc_hd__o21ai_1 _640_ (.A1(_396_),
    .A2(_227_),
    .B1(_194_),
    .Y(_228_));
 sky130_fd_sc_hd__and4bb_1 _641_ (.A_N(_056_),
    .B_N(_061_),
    .C(_095_),
    .D(_101_),
    .X(_229_));
 sky130_fd_sc_hd__o22a_1 _642_ (.A1(_061_),
    .A2(_096_),
    .B1(_102_),
    .B2(_056_),
    .X(_230_));
 sky130_fd_sc_hd__nor2_1 _643_ (.A(_229_),
    .B(_230_),
    .Y(_231_));
 sky130_fd_sc_hd__a21o_1 _644_ (.A1(_197_),
    .A2(_219_),
    .B1(_220_),
    .X(_232_));
 sky130_fd_sc_hd__or4_1 _645_ (.A(_404_),
    .B(_038_),
    .C(_126_),
    .D(_156_),
    .X(_233_));
 sky130_fd_sc_hd__a2bb2o_1 _646_ (.A1_N(_038_),
    .A2_N(_126_),
    .B1(_155_),
    .B2(_403_),
    .X(_234_));
 sky130_fd_sc_hd__and2_1 _647_ (.A(_233_),
    .B(_234_),
    .X(_235_));
 sky130_fd_sc_hd__or2_1 _648_ (.A(_157_),
    .B(_159_),
    .X(_236_));
 sky130_fd_sc_hd__nand2_1 _649_ (.A(_157_),
    .B(_159_),
    .Y(_237_));
 sky130_fd_sc_hd__a41o_1 _650_ (.A1(_157_),
    .A2(_158_),
    .A3(_159_),
    .A4(_160_),
    .B1(_200_),
    .X(_238_));
 sky130_fd_sc_hd__a22o_1 _651_ (.A1(_236_),
    .A2(_237_),
    .B1(_238_),
    .B2(_201_),
    .X(_239_));
 sky130_fd_sc_hd__nand3b_1 _652_ (.A_N(_167_),
    .B(_204_),
    .C(_239_),
    .Y(_240_));
 sky130_fd_sc_hd__a31o_1 _653_ (.A1(_165_),
    .A2(_166_),
    .A3(_204_),
    .B1(_239_),
    .X(_241_));
 sky130_fd_sc_hd__nand3_1 _654_ (.A(_235_),
    .B(_240_),
    .C(_241_),
    .Y(_242_));
 sky130_fd_sc_hd__a21o_1 _655_ (.A1(_240_),
    .A2(_241_),
    .B1(_235_),
    .X(_243_));
 sky130_fd_sc_hd__and3_1 _656_ (.A(_206_),
    .B(_242_),
    .C(_243_),
    .X(_244_));
 sky130_fd_sc_hd__a21oi_1 _657_ (.A1(_242_),
    .A2(_243_),
    .B1(_206_),
    .Y(_245_));
 sky130_fd_sc_hd__a2bb2oi_1 _658_ (.A1_N(_033_),
    .A2_N(_136_),
    .B1(_172_),
    .B2(_399_),
    .Y(_246_));
 sky130_fd_sc_hd__a31oi_1 _659_ (.A1(_412_),
    .A2(_172_),
    .A3(_208_),
    .B1(_246_),
    .Y(_247_));
 sky130_fd_sc_hd__xnor2_1 _660_ (.A(_169_),
    .B(_173_),
    .Y(_248_));
 sky130_fd_sc_hd__nor2_1 _661_ (.A(_175_),
    .B(_211_),
    .Y(_249_));
 sky130_fd_sc_hd__o21ai_2 _662_ (.A1(_212_),
    .A2(_249_),
    .B1(_248_),
    .Y(_250_));
 sky130_fd_sc_hd__nand3_2 _663_ (.A(_181_),
    .B(_215_),
    .C(_250_),
    .Y(_251_));
 sky130_fd_sc_hd__a21o_1 _664_ (.A1(_181_),
    .A2(_215_),
    .B1(_250_),
    .X(_252_));
 sky130_fd_sc_hd__nand3_1 _665_ (.A(_247_),
    .B(_251_),
    .C(_252_),
    .Y(_253_));
 sky130_fd_sc_hd__a21o_1 _666_ (.A1(_251_),
    .A2(_252_),
    .B1(_247_),
    .X(_254_));
 sky130_fd_sc_hd__nand3_1 _667_ (.A(_217_),
    .B(_253_),
    .C(_254_),
    .Y(_255_));
 sky130_fd_sc_hd__a21o_1 _668_ (.A1(_253_),
    .A2(_254_),
    .B1(_217_),
    .X(_256_));
 sky130_fd_sc_hd__or4bb_2 _669_ (.A(_244_),
    .B(_245_),
    .C_N(_255_),
    .D_N(_256_),
    .X(_257_));
 sky130_fd_sc_hd__a2bb2o_1 _670_ (.A1_N(_244_),
    .A2_N(_245_),
    .B1(_255_),
    .B2(_256_),
    .X(_258_));
 sky130_fd_sc_hd__a21o_1 _671_ (.A1(_257_),
    .A2(_258_),
    .B1(_232_),
    .X(_259_));
 sky130_fd_sc_hd__nand3_1 _672_ (.A(_232_),
    .B(_257_),
    .C(_258_),
    .Y(_260_));
 sky130_fd_sc_hd__a21o_1 _673_ (.A1(_259_),
    .A2(_260_),
    .B1(_223_),
    .X(_261_));
 sky130_fd_sc_hd__nand3_1 _674_ (.A(_223_),
    .B(_259_),
    .C(_260_),
    .Y(_262_));
 sky130_fd_sc_hd__and3_1 _675_ (.A(_231_),
    .B(_261_),
    .C(_262_),
    .X(_263_));
 sky130_fd_sc_hd__a21o_1 _676_ (.A1(_261_),
    .A2(_262_),
    .B1(_231_),
    .X(_264_));
 sky130_fd_sc_hd__and2b_1 _677_ (.A_N(_263_),
    .B(_264_),
    .X(_265_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(_225_),
    .B(_265_),
    .Y(_266_));
 sky130_fd_sc_hd__o21ba_1 _679_ (.A1(_396_),
    .A2(_266_),
    .B1_N(_228_),
    .X(_267_));
 sky130_fd_sc_hd__o21a_1 _680_ (.A1(_225_),
    .A2(_263_),
    .B1(_264_),
    .X(_268_));
 sky130_fd_sc_hd__o21a_1 _681_ (.A1(_157_),
    .A2(_159_),
    .B1(_240_),
    .X(_269_));
 sky130_fd_sc_hd__o211a_1 _682_ (.A1(_404_),
    .A2(_126_),
    .B1(_155_),
    .C1(_037_),
    .X(_270_));
 sky130_fd_sc_hd__xnor2_1 _683_ (.A(_269_),
    .B(_270_),
    .Y(_271_));
 sky130_fd_sc_hd__a21bo_1 _684_ (.A1(_206_),
    .A2(_243_),
    .B1_N(_242_),
    .X(_272_));
 sky130_fd_sc_hd__xnor2_1 _685_ (.A(_271_),
    .B(_272_),
    .Y(_273_));
 sky130_fd_sc_hd__o21ai_2 _686_ (.A1(_169_),
    .A2(_173_),
    .B1(_251_),
    .Y(_274_));
 sky130_fd_sc_hd__o211a_1 _687_ (.A1(_400_),
    .A2(_136_),
    .B1(_172_),
    .C1(_412_),
    .X(_275_));
 sky130_fd_sc_hd__xnor2_1 _688_ (.A(_274_),
    .B(_275_),
    .Y(_276_));
 sky130_fd_sc_hd__a21bo_1 _689_ (.A1(_217_),
    .A2(_254_),
    .B1_N(_253_),
    .X(_277_));
 sky130_fd_sc_hd__and2b_1 _690_ (.A_N(_276_),
    .B(_277_),
    .X(_278_));
 sky130_fd_sc_hd__xor2_1 _691_ (.A(_276_),
    .B(_277_),
    .X(_279_));
 sky130_fd_sc_hd__nor2_1 _692_ (.A(_273_),
    .B(_279_),
    .Y(_280_));
 sky130_fd_sc_hd__xor2_1 _693_ (.A(_273_),
    .B(_279_),
    .X(_281_));
 sky130_fd_sc_hd__a21boi_1 _694_ (.A1(_232_),
    .A2(_257_),
    .B1_N(_258_),
    .Y(_282_));
 sky130_fd_sc_hd__xor2_1 _695_ (.A(_281_),
    .B(_282_),
    .X(_283_));
 sky130_fd_sc_hd__nand2b_1 _696_ (.A_N(_261_),
    .B(_283_),
    .Y(_284_));
 sky130_fd_sc_hd__xnor2_1 _697_ (.A(_261_),
    .B(_283_),
    .Y(_285_));
 sky130_fd_sc_hd__nor2_1 _698_ (.A(_061_),
    .B(_126_),
    .Y(_286_));
 sky130_fd_sc_hd__nor2_1 _699_ (.A(_056_),
    .B(_136_),
    .Y(_287_));
 sky130_fd_sc_hd__nor2_1 _700_ (.A(_096_),
    .B(_102_),
    .Y(_288_));
 sky130_fd_sc_hd__a211o_1 _701_ (.A1(_195_),
    .A2(_288_),
    .B1(_287_),
    .C1(_286_),
    .X(_289_));
 sky130_fd_sc_hd__nand2_1 _702_ (.A(_286_),
    .B(_287_),
    .Y(_290_));
 sky130_fd_sc_hd__o211a_1 _703_ (.A1(_286_),
    .A2(_287_),
    .B1(_288_),
    .C1(_195_),
    .X(_291_));
 sky130_fd_sc_hd__inv_2 _704_ (.A(_291_),
    .Y(_292_));
 sky130_fd_sc_hd__and3_1 _705_ (.A(_289_),
    .B(_290_),
    .C(_292_),
    .X(_293_));
 sky130_fd_sc_hd__and2_1 _706_ (.A(_285_),
    .B(_293_),
    .X(_294_));
 sky130_fd_sc_hd__or2_1 _707_ (.A(_285_),
    .B(_293_),
    .X(_295_));
 sky130_fd_sc_hd__and2b_1 _708_ (.A_N(_294_),
    .B(_295_),
    .X(_296_));
 sky130_fd_sc_hd__xnor2_1 _709_ (.A(_268_),
    .B(_296_),
    .Y(_297_));
 sky130_fd_sc_hd__o21ai_2 _710_ (.A1(_396_),
    .A2(_297_),
    .B1(_267_),
    .Y(_298_));
 sky130_fd_sc_hd__o21a_1 _711_ (.A1(_268_),
    .A2(_294_),
    .B1(_295_),
    .X(_299_));
 sky130_fd_sc_hd__o41a_1 _712_ (.A1(_038_),
    .A2(_156_),
    .A3(_198_),
    .A4(_269_),
    .B1(_233_),
    .X(_300_));
 sky130_fd_sc_hd__a21boi_1 _713_ (.A1(_271_),
    .A2(_272_),
    .B1_N(_300_),
    .Y(_301_));
 sky130_fd_sc_hd__o211a_1 _714_ (.A1(_208_),
    .A2(_274_),
    .B1(_412_),
    .C1(_172_),
    .X(_302_));
 sky130_fd_sc_hd__nor2_1 _715_ (.A(_278_),
    .B(_302_),
    .Y(_303_));
 sky130_fd_sc_hd__nor2_1 _716_ (.A(_301_),
    .B(_303_),
    .Y(_304_));
 sky130_fd_sc_hd__xor2_1 _717_ (.A(_301_),
    .B(_303_),
    .X(_305_));
 sky130_fd_sc_hd__a21oi_1 _718_ (.A1(_281_),
    .A2(_282_),
    .B1(_280_),
    .Y(_306_));
 sky130_fd_sc_hd__and2b_1 _719_ (.A_N(_306_),
    .B(_305_),
    .X(_307_));
 sky130_fd_sc_hd__xor2_1 _720_ (.A(_305_),
    .B(_306_),
    .X(_308_));
 sky130_fd_sc_hd__nor2_1 _721_ (.A(_284_),
    .B(_308_),
    .Y(_309_));
 sky130_fd_sc_hd__xor2_1 _722_ (.A(_284_),
    .B(_308_),
    .X(_310_));
 sky130_fd_sc_hd__or4_1 _723_ (.A(_061_),
    .B(_102_),
    .C(_126_),
    .D(_156_),
    .X(_311_));
 sky130_fd_sc_hd__o22ai_1 _724_ (.A1(_102_),
    .A2(_126_),
    .B1(_156_),
    .B2(_061_),
    .Y(_312_));
 sky130_fd_sc_hd__and2_1 _725_ (.A(_311_),
    .B(_312_),
    .X(_313_));
 sky130_fd_sc_hd__or4b_1 _726_ (.A(_056_),
    .B(_096_),
    .C(_136_),
    .D_N(_172_),
    .X(_314_));
 sky130_fd_sc_hd__a2bb2o_1 _727_ (.A1_N(_096_),
    .A2_N(_136_),
    .B1(_172_),
    .B2(_057_),
    .X(_315_));
 sky130_fd_sc_hd__and2_1 _728_ (.A(_314_),
    .B(_315_),
    .X(_316_));
 sky130_fd_sc_hd__nand2_1 _729_ (.A(_313_),
    .B(_316_),
    .Y(_317_));
 sky130_fd_sc_hd__nor2_1 _730_ (.A(_313_),
    .B(_316_),
    .Y(_318_));
 sky130_fd_sc_hd__or2_1 _731_ (.A(_313_),
    .B(_316_),
    .X(_319_));
 sky130_fd_sc_hd__and2_1 _732_ (.A(_317_),
    .B(_319_),
    .X(_320_));
 sky130_fd_sc_hd__xnor2_1 _733_ (.A(_290_),
    .B(_320_),
    .Y(_321_));
 sky130_fd_sc_hd__o21ai_1 _734_ (.A1(_229_),
    .A2(_291_),
    .B1(_321_),
    .Y(_322_));
 sky130_fd_sc_hd__or3_1 _735_ (.A(_229_),
    .B(_291_),
    .C(_321_),
    .X(_323_));
 sky130_fd_sc_hd__and2_1 _736_ (.A(_322_),
    .B(_323_),
    .X(_324_));
 sky130_fd_sc_hd__and2_1 _737_ (.A(_310_),
    .B(_324_),
    .X(_325_));
 sky130_fd_sc_hd__or2_1 _738_ (.A(_310_),
    .B(_324_),
    .X(_326_));
 sky130_fd_sc_hd__xor2_1 _739_ (.A(_310_),
    .B(_324_),
    .X(_327_));
 sky130_fd_sc_hd__xnor2_1 _740_ (.A(_299_),
    .B(_327_),
    .Y(_328_));
 sky130_fd_sc_hd__nor2_1 _741_ (.A(_396_),
    .B(_328_),
    .Y(_329_));
 sky130_fd_sc_hd__nor2_2 _742_ (.A(_126_),
    .B(_136_),
    .Y(_330_));
 sky130_fd_sc_hd__or3_1 _743_ (.A(_102_),
    .B(_156_),
    .C(_286_),
    .X(_331_));
 sky130_fd_sc_hd__or3b_1 _744_ (.A(_096_),
    .B(_287_),
    .C_N(_172_),
    .X(_332_));
 sky130_fd_sc_hd__or2_1 _745_ (.A(_331_),
    .B(_332_),
    .X(_333_));
 sky130_fd_sc_hd__and2_1 _746_ (.A(_331_),
    .B(_332_),
    .X(_334_));
 sky130_fd_sc_hd__nand2_1 _747_ (.A(_331_),
    .B(_332_),
    .Y(_335_));
 sky130_fd_sc_hd__nand2_1 _748_ (.A(_333_),
    .B(_335_),
    .Y(_336_));
 sky130_fd_sc_hd__o21a_1 _749_ (.A1(_290_),
    .A2(_318_),
    .B1(_317_),
    .X(_337_));
 sky130_fd_sc_hd__xnor2_1 _750_ (.A(_336_),
    .B(_337_),
    .Y(_338_));
 sky130_fd_sc_hd__nor2_1 _751_ (.A(_322_),
    .B(_338_),
    .Y(_339_));
 sky130_fd_sc_hd__and2_1 _752_ (.A(_322_),
    .B(_338_),
    .X(_340_));
 sky130_fd_sc_hd__nor2_1 _753_ (.A(_339_),
    .B(_340_),
    .Y(_341_));
 sky130_fd_sc_hd__xor2_1 _754_ (.A(_330_),
    .B(_341_),
    .X(_342_));
 sky130_fd_sc_hd__o31a_1 _755_ (.A1(_304_),
    .A2(_307_),
    .A3(_309_),
    .B1(_342_),
    .X(_343_));
 sky130_fd_sc_hd__nor4_1 _756_ (.A(_304_),
    .B(_307_),
    .C(_309_),
    .D(_342_),
    .Y(_344_));
 sky130_fd_sc_hd__or2_1 _757_ (.A(_343_),
    .B(_344_),
    .X(_345_));
 sky130_fd_sc_hd__a21o_1 _758_ (.A1(_299_),
    .A2(_326_),
    .B1(_325_),
    .X(_346_));
 sky130_fd_sc_hd__xnor2_1 _759_ (.A(_345_),
    .B(_346_),
    .Y(_347_));
 sky130_fd_sc_hd__a211o_1 _760_ (.A1(_395_),
    .A2(_347_),
    .B1(_329_),
    .C1(_298_),
    .X(_348_));
 sky130_fd_sc_hd__nand3_1 _761_ (.A(_155_),
    .B(_172_),
    .C(_330_),
    .Y(_349_));
 sky130_fd_sc_hd__nand2b_1 _762_ (.A_N(_126_),
    .B(_172_),
    .Y(_350_));
 sky130_fd_sc_hd__o21ai_1 _763_ (.A1(_136_),
    .A2(_156_),
    .B1(_350_),
    .Y(_351_));
 sky130_fd_sc_hd__nor2_1 _764_ (.A(_311_),
    .B(_314_),
    .Y(_352_));
 sky130_fd_sc_hd__and2_1 _765_ (.A(_311_),
    .B(_314_),
    .X(_353_));
 sky130_fd_sc_hd__nor2_1 _766_ (.A(_352_),
    .B(_353_),
    .Y(_354_));
 sky130_fd_sc_hd__a21oi_1 _767_ (.A1(_317_),
    .A2(_333_),
    .B1(_334_),
    .Y(_355_));
 sky130_fd_sc_hd__o21a_1 _768_ (.A1(_354_),
    .A2(_355_),
    .B1(_339_),
    .X(_356_));
 sky130_fd_sc_hd__nor3_1 _769_ (.A(_339_),
    .B(_354_),
    .C(_355_),
    .Y(_357_));
 sky130_fd_sc_hd__nor2_1 _770_ (.A(_356_),
    .B(_357_),
    .Y(_358_));
 sky130_fd_sc_hd__and3_1 _771_ (.A(_349_),
    .B(_351_),
    .C(_358_),
    .X(_359_));
 sky130_fd_sc_hd__a21oi_1 _772_ (.A1(_349_),
    .A2(_351_),
    .B1(_358_),
    .Y(_360_));
 sky130_fd_sc_hd__nor2_1 _773_ (.A(_359_),
    .B(_360_),
    .Y(_361_));
 sky130_fd_sc_hd__and3_1 _774_ (.A(_330_),
    .B(_341_),
    .C(_361_),
    .X(_362_));
 sky130_fd_sc_hd__a21oi_1 _775_ (.A1(_330_),
    .A2(_341_),
    .B1(_361_),
    .Y(_363_));
 sky130_fd_sc_hd__nor2_1 _776_ (.A(_362_),
    .B(_363_),
    .Y(_364_));
 sky130_fd_sc_hd__a211o_1 _777_ (.A1(_299_),
    .A2(_326_),
    .B1(_343_),
    .C1(_325_),
    .X(_365_));
 sky130_fd_sc_hd__nand2b_1 _778_ (.A_N(_344_),
    .B(_365_),
    .Y(_366_));
 sky130_fd_sc_hd__and3b_1 _779_ (.A_N(_344_),
    .B(_364_),
    .C(_365_),
    .X(_367_));
 sky130_fd_sc_hd__xnor2_2 _780_ (.A(_364_),
    .B(_366_),
    .Y(_368_));
 sky130_fd_sc_hd__nor2_1 _781_ (.A(_352_),
    .B(_356_),
    .Y(_369_));
 sky130_fd_sc_hd__o211a_1 _782_ (.A1(_126_),
    .A2(_136_),
    .B1(_155_),
    .C1(_172_),
    .X(_370_));
 sky130_fd_sc_hd__xnor2_1 _783_ (.A(_369_),
    .B(_370_),
    .Y(_371_));
 sky130_fd_sc_hd__o21a_1 _784_ (.A1(_359_),
    .A2(_362_),
    .B1(_371_),
    .X(_372_));
 sky130_fd_sc_hd__nor3_1 _785_ (.A(_359_),
    .B(_362_),
    .C(_371_),
    .Y(_373_));
 sky130_fd_sc_hd__nor2_1 _786_ (.A(_372_),
    .B(_373_),
    .Y(_374_));
 sky130_fd_sc_hd__o311a_1 _787_ (.A1(_330_),
    .A2(_352_),
    .A3(_356_),
    .B1(_172_),
    .C1(_155_),
    .X(_375_));
 sky130_fd_sc_hd__a211o_1 _788_ (.A1(_367_),
    .A2(_374_),
    .B1(_375_),
    .C1(_372_),
    .X(_376_));
 sky130_fd_sc_hd__a211o_1 _789_ (.A1(_395_),
    .A2(_368_),
    .B1(_376_),
    .C1(_348_),
    .X(\FP15.d ));
 sky130_fd_sc_hd__xor2_1 _790_ (.A(_367_),
    .B(_374_),
    .X(_377_));
 sky130_fd_sc_hd__a211o_1 _791_ (.A1(_395_),
    .A2(_368_),
    .B1(_377_),
    .C1(_348_),
    .X(\FP14.d ));
 sky130_fd_sc_hd__xor2_1 _792_ (.A(_348_),
    .B(_368_),
    .X(\FP13.d ));
 sky130_fd_sc_hd__or3_1 _793_ (.A(_298_),
    .B(_329_),
    .C(_347_),
    .X(_378_));
 sky130_fd_sc_hd__o21ai_1 _794_ (.A1(_298_),
    .A2(_329_),
    .B1(_347_),
    .Y(_379_));
 sky130_fd_sc_hd__and2_1 _795_ (.A(_378_),
    .B(_379_),
    .X(\FP12.d ));
 sky130_fd_sc_hd__xnor2_1 _796_ (.A(_298_),
    .B(_328_),
    .Y(\FP11.d ));
 sky130_fd_sc_hd__xor2_1 _797_ (.A(_267_),
    .B(_297_),
    .X(\FP10.d ));
 sky130_fd_sc_hd__xnor2_1 _798_ (.A(_228_),
    .B(_266_),
    .Y(\FP9.d ));
 sky130_fd_sc_hd__xor2_1 _799_ (.A(_194_),
    .B(_227_),
    .X(\FP8.d ));
 sky130_fd_sc_hd__xor2_1 _800_ (.A(_150_),
    .B(_193_),
    .X(\FP7.d ));
 sky130_fd_sc_hd__xnor2_1 _801_ (.A(_116_),
    .B(_149_),
    .Y(\FP6.d ));
 sky130_fd_sc_hd__xor2_1 _802_ (.A(_080_),
    .B(_115_),
    .X(\FP5.d ));
 sky130_fd_sc_hd__xor2_1 _803_ (.A(_053_),
    .B(_079_),
    .X(\FP4.d ));
 sky130_fd_sc_hd__xnor2_1 _804_ (.A(_410_),
    .B(_052_),
    .Y(\FP3.d ));
 sky130_fd_sc_hd__nor2_1 _805_ (.A(_409_),
    .B(_043_),
    .Y(_380_));
 sky130_fd_sc_hd__xnor2_1 _806_ (.A(_397_),
    .B(_380_),
    .Y(\FP2.d ));
 sky130_fd_sc_hd__nand2_1 _807_ (.A(\FP0.d ),
    .B(_395_),
    .Y(_381_));
 sky130_fd_sc_hd__nor2_1 _808_ (.A(_394_),
    .B(_047_),
    .Y(_382_));
 sky130_fd_sc_hd__xnor2_1 _809_ (.A(_381_),
    .B(_382_),
    .Y(\FP1.d ));
 sky130_fd_sc_hd__inv_2 _810_ (.A(net19),
    .Y(_001_));
 sky130_fd_sc_hd__inv_2 _811_ (.A(net19),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _812_ (.A(net19),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _813_ (.A(net19),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _814_ (.A(net19),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _815_ (.A(net19),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _816_ (.A(net19),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _817_ (.A(net19),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _818_ (.A(net19),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _819_ (.A(net19),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _820_ (.A(net19),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _821_ (.A(net19),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _822_ (.A(net19),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _823_ (.A(net19),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _824_ (.A(net19),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _825_ (.A(net19),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _826_ (.A(net19),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _827_ (.A(net19),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _828_ (.A(net19),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _829_ (.A(net19),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _830_ (.A(net19),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _831_ (.A(net19),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _832_ (.A(net19),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _833_ (.A(net19),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _834_ (.A(net19),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _835_ (.A(net19),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _836_ (.A(net19),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _837_ (.A(net19),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _838_ (.A(net19),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _839_ (.A(net19),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _840_ (.A(net19),
    .Y(_031_));
 sky130_fd_sc_hd__inv_2 _841_ (.A(net19),
    .Y(_032_));
 sky130_fd_sc_hd__dfrtp_1 _842_ (.CLK(net17),
    .D(\FP0.d ),
    .RESET_B(_000_),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _843_ (.CLK(net17),
    .D(\FP1.d ),
    .RESET_B(_001_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_2 _844_ (.CLK(net17),
    .D(\FP2.d ),
    .RESET_B(_002_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _845_ (.CLK(net17),
    .D(\FP3.d ),
    .RESET_B(_003_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _846_ (.CLK(net17),
    .D(\FP4.d ),
    .RESET_B(_004_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _847_ (.CLK(net17),
    .D(\FP5.d ),
    .RESET_B(_005_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _848_ (.CLK(net17),
    .D(\FP6.d ),
    .RESET_B(_006_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _849_ (.CLK(net17),
    .D(\FP7.d ),
    .RESET_B(_007_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _850_ (.CLK(net17),
    .D(\FP8.d ),
    .RESET_B(_008_),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _851_ (.CLK(net17),
    .D(\FP9.d ),
    .RESET_B(_009_),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _852_ (.CLK(net17),
    .D(\FP10.d ),
    .RESET_B(_010_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _853_ (.CLK(net17),
    .D(\FP11.d ),
    .RESET_B(_011_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _854_ (.CLK(net17),
    .D(\FP12.d ),
    .RESET_B(_012_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _855_ (.CLK(net17),
    .D(\FP13.d ),
    .RESET_B(_013_),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_2 _856_ (.CLK(net17),
    .D(\FP14.d ),
    .RESET_B(_014_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_2 _857_ (.CLK(net17),
    .D(\FP15.d ),
    .RESET_B(_015_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_4 _858_ (.CLK(net17),
    .D(net1),
    .RESET_B(_016_),
    .Q(\FA0.q ));
 sky130_fd_sc_hd__dfrtp_4 _859_ (.CLK(net17),
    .D(net2),
    .RESET_B(_017_),
    .Q(\FA1.q ));
 sky130_fd_sc_hd__dfrtp_4 _860_ (.CLK(net17),
    .D(net3),
    .RESET_B(_018_),
    .Q(\FA2.q ));
 sky130_fd_sc_hd__dfrtp_4 _861_ (.CLK(net17),
    .D(net4),
    .RESET_B(_019_),
    .Q(\FA3.q ));
 sky130_fd_sc_hd__dfrtp_4 _862_ (.CLK(net17),
    .D(net5),
    .RESET_B(_020_),
    .Q(\FA4.q ));
 sky130_fd_sc_hd__dfrtp_4 _863_ (.CLK(net17),
    .D(net6),
    .RESET_B(_021_),
    .Q(\FA5.q ));
 sky130_fd_sc_hd__dfrtp_4 _864_ (.CLK(net17),
    .D(net7),
    .RESET_B(_022_),
    .Q(\FA6.q ));
 sky130_fd_sc_hd__dfrtp_2 _865_ (.CLK(net17),
    .D(net8),
    .RESET_B(_023_),
    .Q(\FA7.q ));
 sky130_fd_sc_hd__dfrtp_4 _866_ (.CLK(net17),
    .D(net9),
    .RESET_B(_024_),
    .Q(\FB0.q ));
 sky130_fd_sc_hd__dfrtp_4 _867_ (.CLK(net17),
    .D(net10),
    .RESET_B(_025_),
    .Q(\FB1.q ));
 sky130_fd_sc_hd__dfrtp_4 _868_ (.CLK(net17),
    .D(net11),
    .RESET_B(_026_),
    .Q(\FB2.q ));
 sky130_fd_sc_hd__dfrtp_4 _869_ (.CLK(net17),
    .D(net12),
    .RESET_B(_027_),
    .Q(\FB3.q ));
 sky130_fd_sc_hd__dfrtp_4 _870_ (.CLK(net17),
    .D(net13),
    .RESET_B(_028_),
    .Q(\FB4.q ));
 sky130_fd_sc_hd__dfrtp_4 _871_ (.CLK(net17),
    .D(net14),
    .RESET_B(_029_),
    .Q(\FB5.q ));
 sky130_fd_sc_hd__dfrtp_2 _872_ (.CLK(net17),
    .D(net15),
    .RESET_B(_030_),
    .Q(\FB6.q ));
 sky130_fd_sc_hd__dfrtp_4 _873_ (.CLK(net17),
    .D(net16),
    .RESET_B(_031_),
    .Q(\FB7.q ));
 sky130_fd_sc_hd__dfrtp_4 _874_ (.CLK(net17),
    .D(net18),
    .RESET_B(_032_),
    .Q(\FC.q ));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_8 input17 (.A(clk),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(control),
    .X(net18));
 sky130_fd_sc_hd__buf_12 input19 (.A(rst),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(p[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(p[10]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(p[11]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(p[12]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(p[13]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(p[14]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(p[15]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(p[1]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(p[2]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(p[3]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(p[4]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(p[5]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(p[6]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(p[7]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(p[8]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(p[9]));
endmodule

