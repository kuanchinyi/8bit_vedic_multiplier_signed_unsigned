magic
tech sky130A
magscale 1 2
timestamp 1726994193
<< viali >>
rect 1409 36125 1443 36159
rect 33149 36125 33183 36159
rect 34345 36057 34379 36091
rect 1593 35989 1627 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 34069 34017 34103 34051
rect 34529 33949 34563 33983
rect 1409 32861 1443 32895
rect 1593 32725 1627 32759
rect 34069 31841 34103 31875
rect 34437 31773 34471 31807
rect 1409 30685 1443 30719
rect 1593 30549 1627 30583
rect 34069 29665 34103 29699
rect 34529 29597 34563 29631
rect 34529 28713 34563 28747
rect 21097 28577 21131 28611
rect 1409 28509 1443 28543
rect 19441 28509 19475 28543
rect 19625 28509 19659 28543
rect 19901 28509 19935 28543
rect 20085 28509 20119 28543
rect 21189 28509 21223 28543
rect 32781 28509 32815 28543
rect 19809 28441 19843 28475
rect 33057 28441 33091 28475
rect 1593 28373 1627 28407
rect 19901 28373 19935 28407
rect 21557 28373 21591 28407
rect 32597 28373 32631 28407
rect 34437 28169 34471 28203
rect 19257 28101 19291 28135
rect 19901 28101 19935 28135
rect 21005 28101 21039 28135
rect 31309 28101 31343 28135
rect 18981 28033 19015 28067
rect 19625 28033 19659 28067
rect 19993 28033 20027 28067
rect 20361 28033 20395 28067
rect 21097 28033 21131 28067
rect 22569 28033 22603 28067
rect 30849 28033 30883 28067
rect 31033 28033 31067 28067
rect 19257 27965 19291 27999
rect 19533 27965 19567 27999
rect 20085 27965 20119 27999
rect 20177 27965 20211 27999
rect 20637 27965 20671 27999
rect 22477 27965 22511 27999
rect 32689 27965 32723 27999
rect 32965 27965 32999 27999
rect 19073 27897 19107 27931
rect 20545 27897 20579 27931
rect 19349 27829 19383 27863
rect 20821 27829 20855 27863
rect 22845 27829 22879 27863
rect 30113 27829 30147 27863
rect 30665 27829 30699 27863
rect 30941 27829 30975 27863
rect 31769 27829 31803 27863
rect 32597 27829 32631 27863
rect 34713 27829 34747 27863
rect 4058 27625 4092 27659
rect 19901 27625 19935 27659
rect 25218 27625 25252 27659
rect 33701 27625 33735 27659
rect 34161 27625 34195 27659
rect 19717 27557 19751 27591
rect 23581 27557 23615 27591
rect 26709 27557 26743 27591
rect 30113 27557 30147 27591
rect 33149 27557 33183 27591
rect 15301 27489 15335 27523
rect 15669 27489 15703 27523
rect 23673 27489 23707 27523
rect 29837 27489 29871 27523
rect 30481 27489 30515 27523
rect 30573 27489 30607 27523
rect 30849 27489 30883 27523
rect 31677 27489 31711 27523
rect 3801 27421 3835 27455
rect 14841 27421 14875 27455
rect 15117 27421 15151 27455
rect 15393 27421 15427 27455
rect 15485 27421 15519 27455
rect 17417 27421 17451 27455
rect 17601 27421 17635 27455
rect 20177 27421 20211 27455
rect 23397 27421 23431 27455
rect 23489 27421 23523 27455
rect 24869 27421 24903 27455
rect 24961 27421 24995 27455
rect 27169 27421 27203 27455
rect 29745 27421 29779 27455
rect 30205 27421 30239 27455
rect 30389 27421 30423 27455
rect 30665 27421 30699 27455
rect 31033 27421 31067 27455
rect 31125 27421 31159 27455
rect 31401 27421 31435 27455
rect 33425 27421 33459 27455
rect 33609 27421 33643 27455
rect 34253 27421 34287 27455
rect 14933 27353 14967 27387
rect 18245 27353 18279 27387
rect 33333 27353 33367 27387
rect 5549 27285 5583 27319
rect 5825 27285 5859 27319
rect 15669 27285 15703 27319
rect 17509 27285 17543 27319
rect 18521 27285 18555 27319
rect 27077 27285 27111 27319
rect 27261 27285 27295 27319
rect 30849 27285 30883 27319
rect 4169 27081 4203 27115
rect 17693 27081 17727 27115
rect 22569 27081 22603 27115
rect 23305 27081 23339 27115
rect 24501 27081 24535 27115
rect 25973 27081 26007 27115
rect 26709 27081 26743 27115
rect 28733 27081 28767 27115
rect 31493 27081 31527 27115
rect 33149 27081 33183 27115
rect 15945 27013 15979 27047
rect 16957 27013 16991 27047
rect 17141 27013 17175 27047
rect 19349 27013 19383 27047
rect 32781 27013 32815 27047
rect 4077 26945 4111 26979
rect 14841 26945 14875 26979
rect 15485 26945 15519 26979
rect 16129 26945 16163 26979
rect 16313 26945 16347 26979
rect 16773 26945 16807 26979
rect 17233 26945 17267 26979
rect 17417 26945 17451 26979
rect 17785 26945 17819 26979
rect 17877 26945 17911 26979
rect 18061 26945 18095 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 18613 26945 18647 26979
rect 18705 26945 18739 26979
rect 18797 26945 18831 26979
rect 19533 26945 19567 26979
rect 19625 26945 19659 26979
rect 20085 26945 20119 26979
rect 20269 26945 20303 26979
rect 20361 26945 20395 26979
rect 20637 26945 20671 26979
rect 21833 26945 21867 26979
rect 22017 26945 22051 26979
rect 22385 26945 22419 26979
rect 24041 26945 24075 26979
rect 24715 26945 24749 26979
rect 24869 26945 24903 26979
rect 25789 26945 25823 26979
rect 25881 26945 25915 26979
rect 26985 26945 27019 26979
rect 29009 26945 29043 26979
rect 30113 26945 30147 26979
rect 31125 26945 31159 26979
rect 33701 26945 33735 26979
rect 34713 26945 34747 26979
rect 14749 26877 14783 26911
rect 15393 26877 15427 26911
rect 18245 26877 18279 26911
rect 20177 26877 20211 26911
rect 20545 26877 20579 26911
rect 22109 26877 22143 26911
rect 22201 26877 22235 26911
rect 23765 26877 23799 26911
rect 23949 26877 23983 26911
rect 27261 26877 27295 26911
rect 30205 26877 30239 26911
rect 31033 26877 31067 26911
rect 15209 26809 15243 26843
rect 15853 26809 15887 26843
rect 18981 26809 19015 26843
rect 23489 26809 23523 26843
rect 30481 26809 30515 26843
rect 3617 26741 3651 26775
rect 4629 26741 4663 26775
rect 19349 26741 19383 26775
rect 24317 26741 24351 26775
rect 28917 26741 28951 26775
rect 29377 26741 29411 26775
rect 5825 26537 5859 26571
rect 15025 26537 15059 26571
rect 16865 26537 16899 26571
rect 18613 26537 18647 26571
rect 20177 26537 20211 26571
rect 20361 26537 20395 26571
rect 21465 26537 21499 26571
rect 21649 26537 21683 26571
rect 22017 26537 22051 26571
rect 22293 26537 22327 26571
rect 26893 26537 26927 26571
rect 28825 26537 28859 26571
rect 30849 26537 30883 26571
rect 34529 26537 34563 26571
rect 7021 26469 7055 26503
rect 11345 26469 11379 26503
rect 25237 26469 25271 26503
rect 1685 26401 1719 26435
rect 3801 26401 3835 26435
rect 9229 26401 9263 26435
rect 13001 26401 13035 26435
rect 13461 26401 13495 26435
rect 18153 26401 18187 26435
rect 22753 26401 22787 26435
rect 24777 26401 24811 26435
rect 27077 26401 27111 26435
rect 1409 26333 1443 26367
rect 6837 26333 6871 26367
rect 8953 26333 8987 26367
rect 12909 26333 12943 26367
rect 13369 26333 13403 26367
rect 13645 26333 13679 26367
rect 15209 26333 15243 26367
rect 15485 26333 15519 26367
rect 16773 26333 16807 26367
rect 16957 26333 16991 26367
rect 17634 26333 17668 26367
rect 18061 26333 18095 26367
rect 18245 26333 18279 26367
rect 18429 26333 18463 26367
rect 20361 26333 20395 26367
rect 20545 26333 20579 26367
rect 21373 26333 21407 26367
rect 21557 26333 21591 26367
rect 21833 26333 21867 26367
rect 22201 26333 22235 26367
rect 22477 26333 22511 26367
rect 22661 26333 22695 26367
rect 24869 26333 24903 26367
rect 32781 26333 32815 26367
rect 3433 26265 3467 26299
rect 4077 26265 4111 26299
rect 10977 26265 11011 26299
rect 13829 26265 13863 26299
rect 15393 26265 15427 26299
rect 17759 26265 17793 26299
rect 27353 26265 27387 26299
rect 30481 26265 30515 26299
rect 30665 26265 30699 26299
rect 33057 26265 33091 26299
rect 5549 26197 5583 26231
rect 13277 26197 13311 26231
rect 17509 26197 17543 26231
rect 31401 26197 31435 26231
rect 32597 26197 32631 26231
rect 1869 25993 1903 26027
rect 4721 25993 4755 26027
rect 6101 25993 6135 26027
rect 9597 25993 9631 26027
rect 13277 25993 13311 26027
rect 17601 25993 17635 26027
rect 17877 25993 17911 26027
rect 19809 25993 19843 26027
rect 21465 25993 21499 26027
rect 21833 25993 21867 26027
rect 22201 25993 22235 26027
rect 29653 25993 29687 26027
rect 31401 25993 31435 26027
rect 33885 25993 33919 26027
rect 34345 25993 34379 26027
rect 2329 25925 2363 25959
rect 3985 25925 4019 25959
rect 16957 25925 16991 25959
rect 19993 25925 20027 25959
rect 28181 25925 28215 25959
rect 29837 25925 29871 25959
rect 34069 25925 34103 25959
rect 1409 25857 1443 25891
rect 1961 25857 1995 25891
rect 4077 25857 4111 25891
rect 4353 25857 4387 25891
rect 4629 25857 4663 25891
rect 5089 25857 5123 25891
rect 5917 25857 5951 25891
rect 9505 25857 9539 25891
rect 12817 25857 12851 25891
rect 12909 25857 12943 25891
rect 13093 25857 13127 25891
rect 13645 25857 13679 25891
rect 16129 25857 16163 25891
rect 16773 25857 16807 25891
rect 18243 25879 18277 25913
rect 20177 25857 20211 25891
rect 20269 25857 20303 25891
rect 20361 25857 20395 25891
rect 20545 25857 20579 25891
rect 21189 25857 21223 25891
rect 21833 25857 21867 25891
rect 22017 25857 22051 25891
rect 22109 25857 22143 25891
rect 22293 25857 22327 25891
rect 29929 25857 29963 25891
rect 31033 25857 31067 25891
rect 31493 25857 31527 25891
rect 31677 25857 31711 25891
rect 34161 25857 34195 25891
rect 34437 25857 34471 25891
rect 34713 25857 34747 25891
rect 2053 25789 2087 25823
rect 5733 25789 5767 25823
rect 13553 25789 13587 25823
rect 15945 25789 15979 25823
rect 16405 25789 16439 25823
rect 17877 25789 17911 25823
rect 17969 25789 18003 25823
rect 18153 25789 18187 25823
rect 20821 25789 20855 25823
rect 21281 25789 21315 25823
rect 27905 25789 27939 25823
rect 31125 25789 31159 25823
rect 31585 25789 31619 25823
rect 32137 25789 32171 25823
rect 32413 25789 32447 25823
rect 3801 25721 3835 25755
rect 14013 25721 14047 25755
rect 1593 25653 1627 25687
rect 9965 25653 9999 25687
rect 14657 25653 14691 25687
rect 15117 25653 15151 25687
rect 16313 25653 16347 25687
rect 17141 25653 17175 25687
rect 20729 25653 20763 25687
rect 27721 25653 27755 25687
rect 30205 25653 30239 25687
rect 5457 25449 5491 25483
rect 8401 25449 8435 25483
rect 10701 25449 10735 25483
rect 16497 25449 16531 25483
rect 18981 25449 19015 25483
rect 20453 25449 20487 25483
rect 21741 25449 21775 25483
rect 22385 25449 22419 25483
rect 23121 25449 23155 25483
rect 26433 25449 26467 25483
rect 14749 25381 14783 25415
rect 16405 25381 16439 25415
rect 20821 25381 20855 25415
rect 24961 25381 24995 25415
rect 31217 25381 31251 25415
rect 5365 25313 5399 25347
rect 11069 25313 11103 25347
rect 11897 25313 11931 25347
rect 13001 25313 13035 25347
rect 16589 25313 16623 25347
rect 20913 25313 20947 25347
rect 24501 25313 24535 25347
rect 25329 25313 25363 25347
rect 25789 25313 25823 25347
rect 28273 25313 28307 25347
rect 30941 25313 30975 25347
rect 34069 25313 34103 25347
rect 5549 25245 5583 25279
rect 5641 25245 5675 25279
rect 12081 25245 12115 25279
rect 15577 25245 15611 25279
rect 16313 25245 16347 25279
rect 18797 25245 18831 25279
rect 18981 25245 19015 25279
rect 20637 25245 20671 25279
rect 21925 25245 21959 25279
rect 22201 25245 22235 25279
rect 22293 25245 22327 25279
rect 22661 25245 22695 25279
rect 22753 25245 22787 25279
rect 23305 25245 23339 25279
rect 23489 25245 23523 25279
rect 24593 25245 24627 25279
rect 25421 25245 25455 25279
rect 26525 25245 26559 25279
rect 30849 25245 30883 25279
rect 34345 25245 34379 25279
rect 10333 25177 10367 25211
rect 26801 25177 26835 25211
rect 2145 25109 2179 25143
rect 3985 25109 4019 25143
rect 5181 25109 5215 25143
rect 14381 25109 14415 25143
rect 15117 25109 15151 25143
rect 16221 25109 16255 25143
rect 17509 25109 17543 25143
rect 22109 25109 22143 25143
rect 32045 25109 32079 25143
rect 11161 24905 11195 24939
rect 11529 24905 11563 24939
rect 12357 24905 12391 24939
rect 12541 24905 12575 24939
rect 14565 24905 14599 24939
rect 14933 24905 14967 24939
rect 15393 24905 15427 24939
rect 16681 24905 16715 24939
rect 23213 24905 23247 24939
rect 23949 24905 23983 24939
rect 24593 24905 24627 24939
rect 25329 24905 25363 24939
rect 30481 24905 30515 24939
rect 31217 24905 31251 24939
rect 34161 24905 34195 24939
rect 15301 24837 15335 24871
rect 15561 24837 15595 24871
rect 15761 24837 15795 24871
rect 17509 24837 17543 24871
rect 15071 24803 15105 24837
rect 1409 24769 1443 24803
rect 3893 24769 3927 24803
rect 4077 24769 4111 24803
rect 4169 24769 4203 24803
rect 4261 24769 4295 24803
rect 4813 24769 4847 24803
rect 5825 24769 5859 24803
rect 6561 24769 6595 24803
rect 8401 24769 8435 24803
rect 10333 24769 10367 24803
rect 11069 24769 11103 24803
rect 11253 24769 11287 24803
rect 11529 24769 11563 24803
rect 11713 24769 11747 24803
rect 12173 24769 12207 24803
rect 12357 24769 12391 24803
rect 12449 24769 12483 24803
rect 12633 24769 12667 24803
rect 13737 24769 13771 24803
rect 14657 24769 14691 24803
rect 14841 24769 14875 24803
rect 16865 24769 16899 24803
rect 16957 24769 16991 24803
rect 17049 24769 17083 24803
rect 18613 24769 18647 24803
rect 18797 24769 18831 24803
rect 18889 24769 18923 24803
rect 19073 24769 19107 24803
rect 19349 24769 19383 24803
rect 23397 24769 23431 24803
rect 23627 24769 23661 24803
rect 24133 24769 24167 24803
rect 24225 24769 24259 24803
rect 24317 24769 24351 24803
rect 24501 24769 24535 24803
rect 24593 24769 24627 24803
rect 24777 24769 24811 24803
rect 25145 24769 25179 24803
rect 25329 24769 25363 24803
rect 26985 24769 27019 24803
rect 29009 24769 29043 24803
rect 30849 24769 30883 24803
rect 30941 24769 30975 24803
rect 4537 24701 4571 24735
rect 4721 24701 4755 24735
rect 5733 24701 5767 24735
rect 6193 24701 6227 24735
rect 6837 24701 6871 24735
rect 8677 24701 8711 24735
rect 10885 24701 10919 24735
rect 18429 24701 18463 24735
rect 23489 24701 23523 24735
rect 23765 24701 23799 24735
rect 23857 24701 23891 24735
rect 30757 24701 30791 24735
rect 31217 24701 31251 24735
rect 32413 24701 32447 24735
rect 32689 24701 32723 24735
rect 3433 24633 3467 24667
rect 12909 24633 12943 24667
rect 13369 24633 13403 24667
rect 14841 24633 14875 24667
rect 16129 24633 16163 24667
rect 17233 24633 17267 24667
rect 18981 24633 19015 24667
rect 31033 24633 31067 24667
rect 1593 24565 1627 24599
rect 3709 24565 3743 24599
rect 5181 24565 5215 24599
rect 8309 24565 8343 24599
rect 10149 24565 10183 24599
rect 11989 24565 12023 24599
rect 14105 24565 14139 24599
rect 15117 24565 15151 24599
rect 15577 24565 15611 24599
rect 16405 24565 16439 24599
rect 18245 24565 18279 24599
rect 28273 24565 28307 24599
rect 30849 24565 30883 24599
rect 31585 24565 31619 24599
rect 31953 24565 31987 24599
rect 34437 24565 34471 24599
rect 4537 24361 4571 24395
rect 5549 24361 5583 24395
rect 5733 24361 5767 24395
rect 9045 24361 9079 24395
rect 9505 24361 9539 24395
rect 10057 24361 10091 24395
rect 14749 24361 14783 24395
rect 15209 24361 15243 24395
rect 15485 24361 15519 24395
rect 18429 24361 18463 24395
rect 19349 24361 19383 24395
rect 27629 24361 27663 24395
rect 31217 24361 31251 24395
rect 33517 24361 33551 24395
rect 15853 24293 15887 24327
rect 17049 24293 17083 24327
rect 21005 24293 21039 24327
rect 33333 24293 33367 24327
rect 1593 24225 1627 24259
rect 1869 24225 1903 24259
rect 3617 24225 3651 24259
rect 4445 24225 4479 24259
rect 14381 24225 14415 24259
rect 16773 24225 16807 24259
rect 17141 24225 17175 24259
rect 27445 24225 27479 24259
rect 31033 24225 31067 24259
rect 31493 24225 31527 24259
rect 3985 24157 4019 24191
rect 4353 24157 4387 24191
rect 8769 24157 8803 24191
rect 9137 24157 9171 24191
rect 9413 24157 9447 24191
rect 10609 24157 10643 24191
rect 11437 24157 11471 24191
rect 12081 24157 12115 24191
rect 12541 24157 12575 24191
rect 13737 24157 13771 24191
rect 13921 24157 13955 24191
rect 14106 24157 14140 24191
rect 14197 24157 14231 24191
rect 14473 24157 14507 24191
rect 14657 24157 14691 24191
rect 14933 24157 14967 24191
rect 15085 24157 15119 24191
rect 15301 24157 15335 24191
rect 15393 24157 15427 24191
rect 15577 24157 15611 24191
rect 16037 24157 16071 24191
rect 16405 24157 16439 24191
rect 16681 24157 16715 24191
rect 17417 24157 17451 24191
rect 18153 24157 18187 24191
rect 18337 24157 18371 24191
rect 18613 24157 18647 24191
rect 19257 24157 19291 24191
rect 19441 24157 19475 24191
rect 19901 24157 19935 24191
rect 20361 24157 20395 24191
rect 20637 24157 20671 24191
rect 20729 24157 20763 24191
rect 27537 24157 27571 24191
rect 30941 24157 30975 24191
rect 31401 24157 31435 24191
rect 31585 24157 31619 24191
rect 33425 24157 33459 24191
rect 3893 24089 3927 24123
rect 5365 24089 5399 24123
rect 13185 24089 13219 24123
rect 13553 24089 13587 24123
rect 13829 24089 13863 24123
rect 16129 24089 16163 24123
rect 17509 24089 17543 24123
rect 17693 24089 17727 24123
rect 20177 24089 20211 24123
rect 20821 24089 20855 24123
rect 21005 24089 21039 24123
rect 4721 24021 4755 24055
rect 5181 24021 5215 24055
rect 5570 24021 5604 24055
rect 10517 24021 10551 24055
rect 12817 24021 12851 24055
rect 14381 24021 14415 24055
rect 14565 24021 14599 24055
rect 16221 24021 16255 24055
rect 17325 24021 17359 24055
rect 18981 24021 19015 24055
rect 20545 24021 20579 24055
rect 31953 24021 31987 24055
rect 4077 23817 4111 23851
rect 15025 23817 15059 23851
rect 15945 23817 15979 23851
rect 16405 23817 16439 23851
rect 21281 23817 21315 23851
rect 23857 23817 23891 23851
rect 25697 23817 25731 23851
rect 27537 23817 27571 23851
rect 29561 23817 29595 23851
rect 1685 23749 1719 23783
rect 8493 23749 8527 23783
rect 9321 23749 9355 23783
rect 12633 23749 12667 23783
rect 13001 23749 13035 23783
rect 23305 23749 23339 23783
rect 23397 23749 23431 23783
rect 28089 23749 28123 23783
rect 29745 23749 29779 23783
rect 6377 23681 6411 23715
rect 9045 23681 9079 23715
rect 12541 23681 12575 23715
rect 12725 23681 12759 23715
rect 12817 23681 12851 23715
rect 13093 23681 13127 23715
rect 13185 23681 13219 23715
rect 13829 23681 13863 23715
rect 14565 23681 14599 23715
rect 15485 23681 15519 23715
rect 15669 23681 15703 23715
rect 18429 23681 18463 23715
rect 18613 23681 18647 23715
rect 20177 23681 20211 23715
rect 20729 23681 20763 23715
rect 21005 23681 21039 23715
rect 21097 23681 21131 23715
rect 21453 23681 21487 23715
rect 21649 23681 21683 23715
rect 21833 23681 21867 23715
rect 22017 23681 22051 23715
rect 22569 23681 22603 23715
rect 22845 23681 22879 23715
rect 22937 23681 22971 23715
rect 23213 23681 23247 23715
rect 23673 23681 23707 23715
rect 25329 23681 25363 23715
rect 27169 23681 27203 23715
rect 27813 23681 27847 23715
rect 29837 23681 29871 23715
rect 1409 23613 1443 23647
rect 13553 23613 13587 23647
rect 15117 23613 15151 23647
rect 15209 23613 15243 23647
rect 17325 23613 17359 23647
rect 20085 23613 20119 23647
rect 20545 23613 20579 23647
rect 20821 23613 20855 23647
rect 23581 23613 23615 23647
rect 25421 23613 25455 23647
rect 26709 23613 26743 23647
rect 27077 23613 27111 23647
rect 3157 23545 3191 23579
rect 11897 23545 11931 23579
rect 13369 23545 13403 23579
rect 14473 23545 14507 23579
rect 14657 23545 14691 23579
rect 15577 23545 15611 23579
rect 21465 23545 21499 23579
rect 22201 23545 22235 23579
rect 26341 23545 26375 23579
rect 3525 23477 3559 23511
rect 4629 23477 4663 23511
rect 6561 23477 6595 23511
rect 8861 23477 8895 23511
rect 9873 23477 9907 23511
rect 11253 23477 11287 23511
rect 12357 23477 12391 23511
rect 16957 23477 16991 23511
rect 23397 23477 23431 23511
rect 26249 23477 26283 23511
rect 30113 23477 30147 23511
rect 2329 23273 2363 23307
rect 4905 23273 4939 23307
rect 6193 23273 6227 23307
rect 8493 23273 8527 23307
rect 13461 23273 13495 23307
rect 14841 23273 14875 23307
rect 15669 23273 15703 23307
rect 18521 23273 18555 23307
rect 20177 23273 20211 23307
rect 21005 23273 21039 23307
rect 22937 23273 22971 23307
rect 24685 23273 24719 23307
rect 26801 23273 26835 23307
rect 27721 23273 27755 23307
rect 4537 23205 4571 23239
rect 5089 23205 5123 23239
rect 15301 23205 15335 23239
rect 21373 23205 21407 23239
rect 24133 23205 24167 23239
rect 24869 23205 24903 23239
rect 4261 23137 4295 23171
rect 5273 23137 5307 23171
rect 5733 23137 5767 23171
rect 7021 23137 7055 23171
rect 9229 23137 9263 23171
rect 10701 23137 10735 23171
rect 14197 23137 14231 23171
rect 17969 23137 18003 23171
rect 23397 23137 23431 23171
rect 23673 23137 23707 23171
rect 34069 23137 34103 23171
rect 2237 23069 2271 23103
rect 4169 23069 4203 23103
rect 5365 23069 5399 23103
rect 5825 23069 5859 23103
rect 6009 23069 6043 23103
rect 6745 23069 6779 23103
rect 8769 23069 8803 23103
rect 8953 23069 8987 23103
rect 10977 23069 11011 23103
rect 12081 23069 12115 23103
rect 12725 23069 12759 23103
rect 14565 23069 14599 23103
rect 14657 23069 14691 23103
rect 18521 23069 18555 23103
rect 18613 23069 18647 23103
rect 19901 23069 19935 23103
rect 20453 23069 20487 23103
rect 20637 23069 20671 23103
rect 20729 23069 20763 23103
rect 21281 23069 21315 23103
rect 22753 23069 22787 23103
rect 23765 23069 23799 23103
rect 24133 23069 24167 23103
rect 24501 23069 24535 23103
rect 24777 23069 24811 23103
rect 25145 23069 25179 23103
rect 25237 23069 25271 23103
rect 25605 23069 25639 23103
rect 26065 23069 26099 23103
rect 26433 23069 26467 23103
rect 26801 23069 26835 23103
rect 26985 23069 27019 23103
rect 34345 23069 34379 23103
rect 4721 23001 4755 23035
rect 8677 23001 8711 23035
rect 11805 23001 11839 23035
rect 12265 23001 12299 23035
rect 14289 23001 14323 23035
rect 18245 23001 18279 23035
rect 20177 23001 20211 23035
rect 20269 23001 20303 23035
rect 21189 23001 21223 23035
rect 22385 23001 22419 23035
rect 22569 23001 22603 23035
rect 24593 23001 24627 23035
rect 2789 22933 2823 22967
rect 3617 22933 3651 22967
rect 4931 22933 4965 22967
rect 13093 22933 13127 22967
rect 13921 22933 13955 22967
rect 17417 22933 17451 22967
rect 19993 22933 20027 22967
rect 20821 22933 20855 22967
rect 20989 22933 21023 22967
rect 22661 22933 22695 22967
rect 4353 22729 4387 22763
rect 5089 22729 5123 22763
rect 9965 22729 9999 22763
rect 24133 22729 24167 22763
rect 2145 22661 2179 22695
rect 3985 22661 4019 22695
rect 4201 22661 4235 22695
rect 6653 22661 6687 22695
rect 8309 22661 8343 22695
rect 16405 22661 16439 22695
rect 18429 22661 18463 22695
rect 22569 22661 22603 22695
rect 24593 22661 24627 22695
rect 5273 22593 5307 22627
rect 5365 22593 5399 22627
rect 8401 22593 8435 22627
rect 8861 22593 8895 22627
rect 9873 22593 9907 22627
rect 10333 22593 10367 22627
rect 12081 22593 12115 22627
rect 12357 22593 12391 22627
rect 15393 22593 15427 22627
rect 16957 22593 16991 22627
rect 17141 22593 17175 22627
rect 17693 22593 17727 22627
rect 18061 22593 18095 22627
rect 18245 22593 18279 22627
rect 22385 22593 22419 22627
rect 24225 22593 24259 22627
rect 24317 22593 24351 22627
rect 24961 22593 24995 22627
rect 25329 22593 25363 22627
rect 25421 22593 25455 22627
rect 1869 22525 1903 22559
rect 5089 22525 5123 22559
rect 6377 22525 6411 22559
rect 8125 22525 8159 22559
rect 9413 22525 9447 22559
rect 12449 22525 12483 22559
rect 23857 22525 23891 22559
rect 3617 22457 3651 22491
rect 10793 22457 10827 22491
rect 12725 22457 12759 22491
rect 17509 22457 17543 22491
rect 18521 22457 18555 22491
rect 4169 22389 4203 22423
rect 4997 22389 5031 22423
rect 14933 22389 14967 22423
rect 17049 22389 17083 22423
rect 22753 22389 22787 22423
rect 23949 22389 23983 22423
rect 2973 22185 3007 22219
rect 3617 22185 3651 22219
rect 4721 22185 4755 22219
rect 4997 22185 5031 22219
rect 8309 22185 8343 22219
rect 14565 22185 14599 22219
rect 15393 22185 15427 22219
rect 15669 22185 15703 22219
rect 20729 22185 20763 22219
rect 21281 22185 21315 22219
rect 21465 22185 21499 22219
rect 22569 22185 22603 22219
rect 23673 22185 23707 22219
rect 23857 22185 23891 22219
rect 32578 22185 32612 22219
rect 34069 22185 34103 22219
rect 16405 22117 16439 22151
rect 16773 22117 16807 22151
rect 18613 22117 18647 22151
rect 24685 22117 24719 22151
rect 31585 22117 31619 22151
rect 15209 22049 15243 22083
rect 17233 22049 17267 22083
rect 17325 22049 17359 22083
rect 18153 22049 18187 22083
rect 19441 22049 19475 22083
rect 31125 22049 31159 22083
rect 31677 22049 31711 22083
rect 32321 22049 32355 22083
rect 1409 21981 1443 22015
rect 2789 21981 2823 22015
rect 2881 21981 2915 22015
rect 4629 21981 4663 22015
rect 4813 21981 4847 22015
rect 13829 21981 13863 22015
rect 14289 21981 14323 22015
rect 14657 21981 14691 22015
rect 15301 21981 15335 22015
rect 15485 21981 15519 22015
rect 15577 21981 15611 22015
rect 15761 21981 15795 22015
rect 16221 21981 16255 22015
rect 16313 21981 16347 22015
rect 16497 21981 16531 22015
rect 16681 21981 16715 22015
rect 17785 21981 17819 22015
rect 18245 21981 18279 22015
rect 19533 21981 19567 22015
rect 21005 21981 21039 22015
rect 21925 21981 21959 22015
rect 22063 21981 22097 22015
rect 22293 21981 22327 22015
rect 22569 21981 22603 22015
rect 22753 21981 22787 22015
rect 23029 21981 23063 22015
rect 23397 21981 23431 22015
rect 24409 21981 24443 22015
rect 24593 21981 24627 22015
rect 31217 21981 31251 22015
rect 31861 21981 31895 22015
rect 21327 21947 21361 21981
rect 16037 21913 16071 21947
rect 17601 21913 17635 21947
rect 20729 21913 20763 21947
rect 21097 21913 21131 21947
rect 22197 21913 22231 21947
rect 23489 21913 23523 21947
rect 32045 21913 32079 21947
rect 1593 21845 1627 21879
rect 4169 21845 4203 21879
rect 7849 21845 7883 21879
rect 8585 21845 8619 21879
rect 9597 21845 9631 21879
rect 11897 21845 11931 21879
rect 13185 21845 13219 21879
rect 13553 21845 13587 21879
rect 14105 21845 14139 21879
rect 17141 21845 17175 21879
rect 17969 21845 18003 21879
rect 20361 21845 20395 21879
rect 20913 21845 20947 21879
rect 22477 21845 22511 21879
rect 23689 21845 23723 21879
rect 9873 21641 9907 21675
rect 11345 21641 11379 21675
rect 11621 21641 11655 21675
rect 11989 21641 12023 21675
rect 13277 21641 13311 21675
rect 17049 21641 17083 21675
rect 17417 21641 17451 21675
rect 18153 21641 18187 21675
rect 20913 21641 20947 21675
rect 23397 21641 23431 21675
rect 26801 21641 26835 21675
rect 30297 21641 30331 21675
rect 31125 21641 31159 21675
rect 31585 21641 31619 21675
rect 33333 21641 33367 21675
rect 2605 21573 2639 21607
rect 10057 21573 10091 21607
rect 10977 21573 11011 21607
rect 14105 21573 14139 21607
rect 28365 21573 28399 21607
rect 28825 21573 28859 21607
rect 30481 21573 30515 21607
rect 2329 21505 2363 21539
rect 4445 21505 4479 21539
rect 4629 21505 4663 21539
rect 4721 21505 4755 21539
rect 4813 21505 4847 21539
rect 5365 21505 5399 21539
rect 8401 21505 8435 21539
rect 9229 21505 9263 21539
rect 9965 21505 9999 21539
rect 10149 21505 10183 21539
rect 10333 21505 10367 21539
rect 11529 21505 11563 21539
rect 11805 21505 11839 21539
rect 13369 21505 13403 21539
rect 13461 21505 13495 21539
rect 13645 21505 13679 21539
rect 13737 21505 13771 21539
rect 14013 21505 14047 21539
rect 14197 21505 14231 21539
rect 17233 21505 17267 21539
rect 17509 21505 17543 21539
rect 17785 21505 17819 21539
rect 17969 21505 18003 21539
rect 18245 21505 18279 21539
rect 18521 21505 18555 21539
rect 20453 21505 20487 21539
rect 20545 21505 20579 21539
rect 20729 21505 20763 21539
rect 22569 21505 22603 21539
rect 23305 21505 23339 21539
rect 23581 21505 23615 21539
rect 25421 21505 25455 21539
rect 26433 21505 26467 21539
rect 28549 21505 28583 21539
rect 30573 21505 30607 21539
rect 30849 21505 30883 21539
rect 31125 21505 31159 21539
rect 31309 21505 31343 21539
rect 33241 21505 33275 21539
rect 4077 21437 4111 21471
rect 5089 21437 5123 21471
rect 5273 21437 5307 21471
rect 6377 21437 6411 21471
rect 6653 21437 6687 21471
rect 8125 21437 8159 21471
rect 10609 21437 10643 21471
rect 17693 21437 17727 21471
rect 22477 21437 22511 21471
rect 22937 21437 22971 21471
rect 25329 21437 25363 21471
rect 26341 21437 26375 21471
rect 5733 21369 5767 21403
rect 18337 21369 18371 21403
rect 23581 21369 23615 21403
rect 25789 21369 25823 21403
rect 10425 21301 10459 21335
rect 10517 21301 10551 21335
rect 13921 21301 13955 21335
rect 14473 21301 14507 21335
rect 15117 21301 15151 21335
rect 15577 21301 15611 21335
rect 18705 21301 18739 21335
rect 32413 21301 32447 21335
rect 33149 21301 33183 21335
rect 3157 21097 3191 21131
rect 3341 21097 3375 21131
rect 4353 21097 4387 21131
rect 5641 21097 5675 21131
rect 7389 21097 7423 21131
rect 10149 21097 10183 21131
rect 17325 21097 17359 21131
rect 17877 21097 17911 21131
rect 23029 21097 23063 21131
rect 26433 21097 26467 21131
rect 5457 21029 5491 21063
rect 9597 21029 9631 21063
rect 11345 21029 11379 21063
rect 13369 21029 13403 21063
rect 5089 20961 5123 20995
rect 5365 20961 5399 20995
rect 11989 20961 12023 20995
rect 12725 20961 12759 20995
rect 15025 20961 15059 20995
rect 15577 20961 15611 20995
rect 20361 20961 20395 20995
rect 25145 20961 25179 20995
rect 3249 20893 3283 20927
rect 4997 20893 5031 20927
rect 7297 20893 7331 20927
rect 9873 20893 9907 20927
rect 10701 20893 10735 20927
rect 10793 20893 10827 20927
rect 11161 20893 11195 20927
rect 11253 20893 11287 20927
rect 11713 20893 11747 20927
rect 12081 20893 12115 20927
rect 12265 20893 12299 20927
rect 13001 20893 13035 20927
rect 14381 20893 14415 20927
rect 14565 20893 14599 20927
rect 14657 20893 14691 20927
rect 14841 20893 14875 20927
rect 14933 20893 14967 20927
rect 15209 20893 15243 20927
rect 15485 20893 15519 20927
rect 15669 20893 15703 20927
rect 17233 20893 17267 20927
rect 17417 20893 17451 20927
rect 17693 20893 17727 20927
rect 17877 20893 17911 20927
rect 21189 20893 21223 20927
rect 21373 20893 21407 20927
rect 21741 20893 21775 20927
rect 24961 20893 24995 20927
rect 25513 20893 25547 20927
rect 25605 20893 25639 20927
rect 25789 20893 25823 20927
rect 25973 20893 26007 20927
rect 26249 20893 26283 20927
rect 33333 20893 33367 20927
rect 5825 20825 5859 20859
rect 6101 20825 6135 20859
rect 8309 20825 8343 20859
rect 9505 20825 9539 20859
rect 9965 20825 9999 20859
rect 10517 20825 10551 20859
rect 11069 20825 11103 20859
rect 11621 20825 11655 20859
rect 12173 20825 12207 20859
rect 14473 20825 14507 20859
rect 34345 20825 34379 20859
rect 5615 20757 5649 20791
rect 7757 20757 7791 20791
rect 8769 20757 8803 20791
rect 9781 20757 9815 20791
rect 10977 20757 11011 20791
rect 11529 20757 11563 20791
rect 12909 20757 12943 20791
rect 13921 20757 13955 20791
rect 15393 20757 15427 20791
rect 15945 20757 15979 20791
rect 9689 20553 9723 20587
rect 11069 20553 11103 20587
rect 11621 20553 11655 20587
rect 12817 20553 12851 20587
rect 14289 20553 14323 20587
rect 15025 20553 15059 20587
rect 15577 20553 15611 20587
rect 17601 20553 17635 20587
rect 20913 20553 20947 20587
rect 22293 20553 22327 20587
rect 24593 20553 24627 20587
rect 33977 20553 34011 20587
rect 6653 20485 6687 20519
rect 12081 20485 12115 20519
rect 21373 20485 21407 20519
rect 24869 20485 24903 20519
rect 6377 20417 6411 20451
rect 8309 20417 8343 20451
rect 9965 20417 9999 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 12633 20417 12667 20451
rect 12817 20417 12851 20451
rect 13088 20417 13122 20451
rect 13185 20417 13219 20451
rect 13277 20417 13311 20451
rect 13405 20417 13439 20451
rect 13553 20417 13587 20451
rect 13645 20417 13679 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 14105 20417 14139 20451
rect 15209 20417 15243 20451
rect 15761 20417 15795 20451
rect 17233 20417 17267 20451
rect 17417 20417 17451 20451
rect 18061 20417 18095 20451
rect 18981 20417 19015 20451
rect 20453 20417 20487 20451
rect 20545 20417 20579 20451
rect 20637 20417 20671 20451
rect 21005 20417 21039 20451
rect 21189 20417 21223 20451
rect 22937 20417 22971 20451
rect 23121 20417 23155 20451
rect 23397 20417 23431 20451
rect 24777 20417 24811 20451
rect 24961 20417 24995 20451
rect 25145 20417 25179 20451
rect 25237 20417 25271 20451
rect 26249 20417 26283 20451
rect 8125 20349 8159 20383
rect 9137 20349 9171 20383
rect 10057 20349 10091 20383
rect 10333 20349 10367 20383
rect 15485 20349 15519 20383
rect 16037 20349 16071 20383
rect 17969 20349 18003 20383
rect 18889 20349 18923 20383
rect 19809 20349 19843 20383
rect 20729 20349 20763 20383
rect 26157 20349 26191 20383
rect 32229 20349 32263 20383
rect 32505 20349 32539 20383
rect 12449 20281 12483 20315
rect 12909 20281 12943 20315
rect 13921 20281 13955 20315
rect 14933 20281 14967 20315
rect 18429 20281 18463 20315
rect 15393 20213 15427 20247
rect 15945 20213 15979 20247
rect 16405 20213 16439 20247
rect 17049 20213 17083 20247
rect 22569 20213 22603 20247
rect 23029 20213 23063 20247
rect 26525 20213 26559 20247
rect 31953 20213 31987 20247
rect 7389 20009 7423 20043
rect 8309 20009 8343 20043
rect 11069 20009 11103 20043
rect 13185 20009 13219 20043
rect 14289 20009 14323 20043
rect 14933 20009 14967 20043
rect 16313 20009 16347 20043
rect 16957 20009 16991 20043
rect 17141 20009 17175 20043
rect 20821 20009 20855 20043
rect 21649 20009 21683 20043
rect 24961 20009 24995 20043
rect 25881 20009 25915 20043
rect 26065 20009 26099 20043
rect 30113 20009 30147 20043
rect 31677 20009 31711 20043
rect 32045 20009 32079 20043
rect 33333 20009 33367 20043
rect 20913 19941 20947 19975
rect 31585 19941 31619 19975
rect 17509 19873 17543 19907
rect 23397 19873 23431 19907
rect 24225 19873 24259 19907
rect 27261 19873 27295 19907
rect 31125 19873 31159 19907
rect 31769 19873 31803 19907
rect 1409 19805 1443 19839
rect 7297 19805 7331 19839
rect 11805 19805 11839 19839
rect 11897 19805 11931 19839
rect 13369 19805 13403 19839
rect 13461 19805 13495 19839
rect 13737 19805 13771 19839
rect 13829 19805 13863 19839
rect 20361 19805 20395 19839
rect 20637 19805 20671 19839
rect 22109 19805 22143 19839
rect 22385 19805 22419 19839
rect 22569 19805 22603 19839
rect 22661 19805 22695 19839
rect 22845 19805 22879 19839
rect 25237 19805 25271 19839
rect 25421 19805 25455 19839
rect 25605 19805 25639 19839
rect 25697 19805 25731 19839
rect 26893 19805 26927 19839
rect 27077 19805 27111 19839
rect 27353 19805 27387 19839
rect 29745 19805 29779 19839
rect 31217 19805 31251 19839
rect 31677 19805 31711 19839
rect 33241 19805 33275 19839
rect 11437 19737 11471 19771
rect 12725 19737 12759 19771
rect 13553 19737 13587 19771
rect 16773 19737 16807 19771
rect 20453 19737 20487 19771
rect 21097 19737 21131 19771
rect 21281 19737 21315 19771
rect 22477 19737 22511 19771
rect 25329 19737 25363 19771
rect 26249 19737 26283 19771
rect 26985 19737 27019 19771
rect 1593 19669 1627 19703
rect 7757 19669 7791 19703
rect 12081 19669 12115 19703
rect 13093 19669 13127 19703
rect 15485 19669 15519 19703
rect 16681 19669 16715 19703
rect 16983 19669 17017 19703
rect 23029 19669 23063 19703
rect 26065 19669 26099 19703
rect 27721 19669 27755 19703
rect 29653 19669 29687 19703
rect 33149 19669 33183 19703
rect 9873 19465 9907 19499
rect 10241 19465 10275 19499
rect 11989 19465 12023 19499
rect 12081 19465 12115 19499
rect 13829 19465 13863 19499
rect 16497 19465 16531 19499
rect 16865 19465 16899 19499
rect 17509 19465 17543 19499
rect 17969 19465 18003 19499
rect 25506 19465 25540 19499
rect 28365 19465 28399 19499
rect 30205 19465 30239 19499
rect 31125 19465 31159 19499
rect 9965 19397 9999 19431
rect 14933 19397 14967 19431
rect 16773 19397 16807 19431
rect 25421 19397 25455 19431
rect 28733 19397 28767 19431
rect 10057 19329 10091 19363
rect 12449 19329 12483 19363
rect 12633 19329 12667 19363
rect 12725 19329 12759 19363
rect 12909 19329 12943 19363
rect 13737 19329 13771 19363
rect 13921 19329 13955 19363
rect 15117 19329 15151 19363
rect 15761 19329 15795 19363
rect 18061 19329 18095 19363
rect 18797 19329 18831 19363
rect 18889 19329 18923 19363
rect 19073 19329 19107 19363
rect 20637 19329 20671 19363
rect 22109 19329 22143 19363
rect 25329 19329 25363 19363
rect 25605 19329 25639 19363
rect 28457 19329 28491 19363
rect 31400 19351 31434 19385
rect 10517 19261 10551 19295
rect 11529 19261 11563 19295
rect 11713 19261 11747 19295
rect 11805 19261 11839 19295
rect 12173 19261 12207 19295
rect 15485 19261 15519 19295
rect 15669 19261 15703 19295
rect 16865 19261 16899 19295
rect 17693 19261 17727 19295
rect 17785 19261 17819 19295
rect 18153 19261 18187 19295
rect 20545 19261 20579 19295
rect 22017 19261 22051 19295
rect 22937 19261 22971 19295
rect 31033 19261 31067 19295
rect 31125 19261 31159 19295
rect 9597 19193 9631 19227
rect 9689 19193 9723 19227
rect 12265 19193 12299 19227
rect 12541 19193 12575 19227
rect 13553 19193 13587 19227
rect 15301 19193 15335 19227
rect 21005 19193 21039 19227
rect 9229 19125 9263 19159
rect 10977 19125 11011 19159
rect 11253 19125 11287 19159
rect 13277 19125 13311 19159
rect 14289 19125 14323 19159
rect 16129 19125 16163 19159
rect 17325 19125 17359 19159
rect 19257 19125 19291 19159
rect 23213 19125 23247 19159
rect 31309 19125 31343 19159
rect 12541 18921 12575 18955
rect 14381 18921 14415 18955
rect 14933 18921 14967 18955
rect 15669 18921 15703 18955
rect 16129 18921 16163 18955
rect 17141 18921 17175 18955
rect 19073 18921 19107 18955
rect 25513 18921 25547 18955
rect 26801 18921 26835 18955
rect 31309 18921 31343 18955
rect 9505 18853 9539 18887
rect 15853 18853 15887 18887
rect 20361 18853 20395 18887
rect 25973 18853 26007 18887
rect 27721 18853 27755 18887
rect 28641 18853 28675 18887
rect 12173 18785 12207 18819
rect 12265 18785 12299 18819
rect 12357 18785 12391 18819
rect 16773 18785 16807 18819
rect 19257 18785 19291 18819
rect 19625 18785 19659 18819
rect 19901 18785 19935 18819
rect 27905 18785 27939 18819
rect 28089 18785 28123 18819
rect 31677 18785 31711 18819
rect 32137 18785 32171 18819
rect 34069 18785 34103 18819
rect 9413 18717 9447 18751
rect 9505 18717 9539 18751
rect 9781 18717 9815 18751
rect 10333 18717 10367 18751
rect 12081 18717 12115 18751
rect 15761 18717 15795 18751
rect 15945 18717 15979 18751
rect 16037 18717 16071 18751
rect 16221 18717 16255 18751
rect 17049 18717 17083 18751
rect 17233 18717 17267 18751
rect 18245 18717 18279 18751
rect 18429 18717 18463 18751
rect 18521 18717 18555 18751
rect 18889 18717 18923 18751
rect 19717 18717 19751 18751
rect 19993 18717 20027 18751
rect 20177 18717 20211 18751
rect 22385 18717 22419 18751
rect 22569 18717 22603 18751
rect 22753 18717 22787 18751
rect 24961 18717 24995 18751
rect 25237 18717 25271 18751
rect 25605 18717 25639 18751
rect 25697 18717 25731 18751
rect 26985 18717 27019 18751
rect 27077 18717 27111 18751
rect 27261 18717 27295 18751
rect 27353 18717 27387 18751
rect 27445 18717 27479 18751
rect 28181 18717 28215 18751
rect 28917 18717 28951 18751
rect 29377 18717 29411 18751
rect 29561 18717 29595 18751
rect 31585 18717 31619 18751
rect 32045 18717 32079 18751
rect 32229 18717 32263 18751
rect 32505 18717 32539 18751
rect 34529 18717 34563 18751
rect 15301 18649 15335 18683
rect 15485 18649 15519 18683
rect 18705 18649 18739 18683
rect 18797 18649 18831 18683
rect 22477 18649 22511 18683
rect 23765 18649 23799 18683
rect 25973 18649 26007 18683
rect 28641 18649 28675 18683
rect 29837 18649 29871 18683
rect 13185 18581 13219 18615
rect 13461 18581 13495 18615
rect 13921 18581 13955 18615
rect 17601 18581 17635 18615
rect 18429 18581 18463 18615
rect 19349 18581 19383 18615
rect 19441 18581 19475 18615
rect 22017 18581 22051 18615
rect 25789 18581 25823 18615
rect 28549 18581 28583 18615
rect 28825 18581 28859 18615
rect 31953 18581 31987 18615
rect 4169 18377 4203 18411
rect 9413 18377 9447 18411
rect 12081 18377 12115 18411
rect 14749 18377 14783 18411
rect 15117 18377 15151 18411
rect 18889 18377 18923 18411
rect 19073 18377 19107 18411
rect 19441 18377 19475 18411
rect 19809 18377 19843 18411
rect 22845 18377 22879 18411
rect 30113 18377 30147 18411
rect 30297 18377 30331 18411
rect 34529 18377 34563 18411
rect 1685 18309 1719 18343
rect 10241 18309 10275 18343
rect 10885 18309 10919 18343
rect 11529 18309 11563 18343
rect 13369 18309 13403 18343
rect 15301 18309 15335 18343
rect 18797 18309 18831 18343
rect 19533 18309 19567 18343
rect 33057 18309 33091 18343
rect 3341 18241 3375 18275
rect 3433 18241 3467 18275
rect 9045 18241 9079 18275
rect 9873 18241 9907 18275
rect 10149 18241 10183 18275
rect 10977 18241 11011 18275
rect 11161 18241 11195 18275
rect 11713 18241 11747 18275
rect 11989 18241 12023 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 12633 18241 12667 18275
rect 12909 18241 12943 18275
rect 13001 18241 13035 18275
rect 13553 18241 13587 18275
rect 14013 18241 14047 18275
rect 14657 18241 14691 18275
rect 14841 18241 14875 18275
rect 15209 18241 15243 18275
rect 15485 18241 15519 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 16129 18241 16163 18275
rect 18613 18241 18647 18275
rect 18889 18241 18923 18275
rect 18981 18241 19015 18275
rect 19257 18241 19291 18275
rect 19717 18241 19751 18275
rect 19809 18241 19843 18275
rect 22753 18241 22787 18275
rect 22937 18241 22971 18275
rect 23213 18241 23247 18275
rect 30205 18241 30239 18275
rect 1409 18173 1443 18207
rect 11897 18173 11931 18207
rect 13829 18173 13863 18207
rect 14381 18173 14415 18207
rect 22293 18173 22327 18207
rect 32781 18173 32815 18207
rect 3157 18037 3191 18071
rect 3709 18037 3743 18071
rect 9781 18037 9815 18071
rect 10701 18037 10735 18071
rect 12449 18037 12483 18071
rect 12725 18037 12759 18071
rect 13185 18037 13219 18071
rect 13737 18037 13771 18071
rect 14197 18037 14231 18071
rect 14473 18037 14507 18071
rect 16957 18037 16991 18071
rect 22569 18037 22603 18071
rect 32689 18037 32723 18071
rect 4077 17833 4111 17867
rect 4353 17833 4387 17867
rect 10609 17833 10643 17867
rect 11069 17833 11103 17867
rect 11989 17833 12023 17867
rect 13277 17833 13311 17867
rect 14381 17833 14415 17867
rect 15025 17833 15059 17867
rect 19625 17833 19659 17867
rect 20729 17833 20763 17867
rect 27353 17833 27387 17867
rect 27721 17833 27755 17867
rect 28273 17833 28307 17867
rect 33793 17833 33827 17867
rect 11529 17765 11563 17799
rect 11621 17765 11655 17799
rect 11897 17765 11931 17799
rect 13185 17765 13219 17799
rect 14749 17765 14783 17799
rect 23029 17765 23063 17799
rect 28825 17765 28859 17799
rect 3985 17697 4019 17731
rect 5457 17697 5491 17731
rect 5733 17697 5767 17731
rect 12081 17697 12115 17731
rect 20177 17697 20211 17731
rect 22569 17697 22603 17731
rect 23213 17697 23247 17731
rect 24593 17697 24627 17731
rect 1409 17629 1443 17663
rect 3893 17629 3927 17663
rect 4169 17629 4203 17663
rect 5365 17629 5399 17663
rect 6193 17629 6227 17663
rect 6285 17629 6319 17663
rect 11805 17629 11839 17663
rect 12541 17629 12575 17663
rect 12725 17629 12759 17663
rect 13001 17629 13035 17663
rect 13553 17629 13587 17663
rect 13645 17629 13679 17663
rect 13737 17629 13771 17663
rect 13921 17629 13955 17663
rect 16589 17629 16623 17663
rect 16865 17629 16899 17663
rect 19809 17629 19843 17663
rect 19993 17629 20027 17663
rect 20453 17629 20487 17663
rect 20545 17629 20579 17663
rect 21005 17629 21039 17663
rect 21189 17629 21223 17663
rect 21465 17629 21499 17663
rect 22201 17629 22235 17663
rect 22477 17629 22511 17663
rect 22661 17629 22695 17663
rect 22753 17629 22787 17663
rect 23121 17629 23155 17663
rect 23305 17629 23339 17663
rect 23581 17629 23615 17663
rect 23765 17629 23799 17663
rect 24685 17629 24719 17663
rect 27629 17629 27663 17663
rect 27721 17629 27755 17663
rect 27813 17629 27847 17663
rect 27997 17629 28031 17663
rect 28549 17629 28583 17663
rect 28641 17629 28675 17663
rect 33701 17629 33735 17663
rect 9965 17561 9999 17595
rect 11161 17561 11195 17595
rect 20085 17561 20119 17595
rect 23029 17561 23063 17595
rect 27353 17561 27387 17595
rect 28089 17561 28123 17595
rect 28825 17561 28859 17595
rect 1593 17493 1627 17527
rect 6469 17493 6503 17527
rect 6745 17493 6779 17527
rect 9321 17493 9355 17527
rect 10241 17493 10275 17527
rect 12449 17493 12483 17527
rect 17601 17493 17635 17527
rect 20821 17493 20855 17527
rect 22845 17493 22879 17527
rect 23397 17493 23431 17527
rect 25513 17493 25547 17527
rect 27537 17493 27571 17527
rect 28289 17493 28323 17527
rect 28457 17493 28491 17527
rect 33609 17493 33643 17527
rect 3525 17289 3559 17323
rect 23489 17289 23523 17323
rect 25697 17289 25731 17323
rect 27813 17289 27847 17323
rect 29285 17289 29319 17323
rect 31493 17289 31527 17323
rect 6837 17221 6871 17255
rect 9137 17221 9171 17255
rect 10149 17221 10183 17255
rect 10885 17221 10919 17255
rect 13277 17221 13311 17255
rect 13553 17221 13587 17255
rect 18337 17221 18371 17255
rect 21097 17221 21131 17255
rect 21281 17221 21315 17255
rect 21465 17221 21499 17255
rect 27445 17221 27479 17255
rect 3893 17153 3927 17187
rect 4997 17153 5031 17187
rect 6929 17153 6963 17187
rect 9229 17153 9263 17187
rect 9321 17153 9355 17187
rect 11989 17153 12023 17187
rect 12265 17153 12299 17187
rect 12633 17153 12667 17187
rect 12796 17153 12830 17187
rect 12909 17153 12943 17187
rect 13001 17153 13035 17187
rect 15853 17153 15887 17187
rect 16313 17153 16347 17187
rect 16497 17153 16531 17187
rect 20453 17153 20487 17187
rect 23121 17153 23155 17187
rect 23305 17153 23339 17187
rect 25237 17153 25271 17187
rect 26157 17153 26191 17187
rect 27353 17153 27387 17187
rect 27629 17153 27663 17187
rect 28641 17153 28675 17187
rect 28825 17153 28859 17187
rect 29377 17153 29411 17187
rect 31677 17153 31711 17187
rect 31861 17153 31895 17187
rect 3801 17085 3835 17119
rect 5089 17085 5123 17119
rect 7205 17085 7239 17119
rect 7481 17085 7515 17119
rect 8953 17085 8987 17119
rect 15761 17085 15795 17119
rect 18245 17085 18279 17119
rect 18337 17085 18371 17119
rect 20545 17085 20579 17119
rect 24777 17085 24811 17119
rect 25053 17085 25087 17119
rect 25145 17085 25179 17119
rect 25881 17085 25915 17119
rect 25973 17085 26007 17119
rect 26065 17085 26099 17119
rect 29653 17085 29687 17119
rect 31125 17085 31159 17119
rect 5365 17017 5399 17051
rect 12173 17017 12207 17051
rect 16221 17017 16255 17051
rect 18797 17017 18831 17051
rect 20821 17017 20855 17051
rect 24593 17017 24627 17051
rect 28641 17017 28675 17051
rect 4261 16949 4295 16983
rect 7021 16949 7055 16983
rect 11161 16949 11195 16983
rect 11713 16949 11747 16983
rect 16405 16949 16439 16983
rect 25605 16949 25639 16983
rect 3801 16745 3835 16779
rect 5181 16745 5215 16779
rect 8217 16745 8251 16779
rect 8677 16745 8711 16779
rect 11621 16745 11655 16779
rect 12357 16745 12391 16779
rect 12817 16745 12851 16779
rect 16497 16745 16531 16779
rect 19257 16745 19291 16779
rect 20453 16745 20487 16779
rect 22477 16745 22511 16779
rect 23581 16745 23615 16779
rect 25513 16745 25547 16779
rect 26249 16745 26283 16779
rect 30389 16745 30423 16779
rect 32873 16745 32907 16779
rect 21373 16677 21407 16711
rect 29285 16677 29319 16711
rect 30757 16677 30791 16711
rect 32321 16677 32355 16711
rect 1685 16609 1719 16643
rect 4077 16609 4111 16643
rect 6469 16609 6503 16643
rect 9689 16609 9723 16643
rect 11069 16609 11103 16643
rect 11989 16609 12023 16643
rect 15209 16609 15243 16643
rect 15853 16609 15887 16643
rect 16037 16609 16071 16643
rect 25789 16609 25823 16643
rect 32045 16609 32079 16643
rect 32505 16609 32539 16643
rect 1409 16541 1443 16575
rect 3433 16541 3467 16575
rect 3977 16541 4011 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 4445 16541 4479 16575
rect 4537 16541 4571 16575
rect 4700 16541 4734 16575
rect 4813 16538 4847 16572
rect 4905 16541 4939 16575
rect 6193 16541 6227 16575
rect 14197 16541 14231 16575
rect 14381 16541 14415 16575
rect 15761 16541 15795 16575
rect 15945 16541 15979 16575
rect 16129 16541 16163 16575
rect 16313 16541 16347 16575
rect 16681 16541 16715 16575
rect 16865 16541 16899 16575
rect 17141 16541 17175 16575
rect 17325 16541 17359 16575
rect 18613 16541 18647 16575
rect 18889 16541 18923 16575
rect 19441 16541 19475 16575
rect 19717 16541 19751 16575
rect 19901 16541 19935 16575
rect 20821 16541 20855 16575
rect 21005 16541 21039 16575
rect 23949 16541 23983 16575
rect 24133 16541 24167 16575
rect 24593 16541 24627 16575
rect 24869 16541 24903 16575
rect 25053 16541 25087 16575
rect 25329 16541 25363 16575
rect 25881 16541 25915 16575
rect 29745 16541 29779 16575
rect 30021 16541 30055 16575
rect 30297 16541 30331 16575
rect 31953 16541 31987 16575
rect 32413 16541 32447 16575
rect 32597 16541 32631 16575
rect 34529 16541 34563 16575
rect 3341 16473 3375 16507
rect 8953 16473 8987 16507
rect 24041 16473 24075 16507
rect 33609 16473 33643 16507
rect 3157 16405 3191 16439
rect 7941 16405 7975 16439
rect 18521 16405 18555 16439
rect 18705 16405 18739 16439
rect 19073 16405 19107 16439
rect 21005 16405 21039 16439
rect 10333 16201 10367 16235
rect 10977 16201 11011 16235
rect 12357 16201 12391 16235
rect 13645 16201 13679 16235
rect 14013 16201 14047 16235
rect 14289 16201 14323 16235
rect 18245 16201 18279 16235
rect 19257 16201 19291 16235
rect 22937 16201 22971 16235
rect 25237 16201 25271 16235
rect 27445 16201 27479 16235
rect 27813 16201 27847 16235
rect 34713 16201 34747 16235
rect 3341 16133 3375 16167
rect 12541 16133 12575 16167
rect 13369 16133 13403 16167
rect 19073 16133 19107 16167
rect 22753 16133 22787 16167
rect 33241 16133 33275 16167
rect 6377 16065 6411 16099
rect 9965 16065 9999 16099
rect 11069 16065 11103 16099
rect 11161 16065 11195 16099
rect 11345 16065 11379 16099
rect 11713 16065 11747 16099
rect 12449 16065 12483 16099
rect 12725 16065 12759 16099
rect 13829 16065 13863 16099
rect 14013 16065 14047 16099
rect 14105 16065 14139 16099
rect 14289 16065 14323 16099
rect 14657 16065 14691 16099
rect 18429 16065 18463 16099
rect 18613 16065 18647 16099
rect 19257 16065 19291 16099
rect 19441 16065 19475 16099
rect 19717 16065 19751 16099
rect 22201 16065 22235 16099
rect 22661 16065 22695 16099
rect 22845 16065 22879 16099
rect 22937 16065 22971 16099
rect 23121 16065 23155 16099
rect 23397 16065 23431 16099
rect 24777 16065 24811 16099
rect 27353 16065 27387 16099
rect 27629 16065 27663 16099
rect 28181 16065 28215 16099
rect 11805 15997 11839 16031
rect 12173 15997 12207 16031
rect 22109 15997 22143 16031
rect 22569 15997 22603 16031
rect 27997 15997 28031 16031
rect 32965 15997 32999 16031
rect 10701 15929 10735 15963
rect 10793 15929 10827 15963
rect 16313 15929 16347 15963
rect 3709 15861 3743 15895
rect 4353 15861 4387 15895
rect 6561 15861 6595 15895
rect 11989 15861 12023 15895
rect 15669 15861 15703 15895
rect 17877 15861 17911 15895
rect 18521 15861 18555 15895
rect 20177 15861 20211 15895
rect 23857 15861 23891 15895
rect 25053 15861 25087 15895
rect 28365 15861 28399 15895
rect 32781 15861 32815 15895
rect 3617 15657 3651 15691
rect 4813 15657 4847 15691
rect 9137 15657 9171 15691
rect 13461 15657 13495 15691
rect 15945 15657 15979 15691
rect 22845 15657 22879 15691
rect 33977 15657 34011 15691
rect 16589 15589 16623 15623
rect 20453 15589 20487 15623
rect 23121 15589 23155 15623
rect 27261 15589 27295 15623
rect 1869 15521 1903 15555
rect 15117 15521 15151 15555
rect 21005 15521 21039 15555
rect 21741 15521 21775 15555
rect 23581 15521 23615 15555
rect 24685 15521 24719 15555
rect 28089 15521 28123 15555
rect 29837 15521 29871 15555
rect 30113 15521 30147 15555
rect 30481 15521 30515 15555
rect 1409 15453 1443 15487
rect 3985 15453 4019 15487
rect 7481 15453 7515 15487
rect 7849 15453 7883 15487
rect 8309 15453 8343 15487
rect 14197 15453 14231 15487
rect 14381 15453 14415 15487
rect 15301 15453 15335 15487
rect 15485 15453 15519 15487
rect 15577 15453 15611 15487
rect 15669 15453 15703 15487
rect 16037 15453 16071 15487
rect 16221 15453 16255 15487
rect 16405 15453 16439 15487
rect 16497 15453 16531 15487
rect 17141 15453 17175 15487
rect 17233 15453 17267 15487
rect 17785 15453 17819 15487
rect 18153 15453 18187 15487
rect 19533 15453 19567 15487
rect 19625 15453 19659 15487
rect 20361 15453 20395 15487
rect 20453 15453 20487 15487
rect 20913 15453 20947 15487
rect 23489 15453 23523 15487
rect 23673 15453 23707 15487
rect 23771 15453 23805 15487
rect 23949 15453 23983 15487
rect 25973 15453 26007 15487
rect 26985 15453 27019 15487
rect 27353 15453 27387 15487
rect 27905 15453 27939 15487
rect 28181 15453 28215 15487
rect 28641 15453 28675 15487
rect 29193 15453 29227 15487
rect 29745 15453 29779 15487
rect 30573 15453 30607 15487
rect 33793 15453 33827 15487
rect 33885 15453 33919 15487
rect 4859 15419 4893 15453
rect 2145 15385 2179 15419
rect 3893 15385 3927 15419
rect 4445 15385 4479 15419
rect 4629 15385 4663 15419
rect 18981 15385 19015 15419
rect 19809 15385 19843 15419
rect 23857 15385 23891 15419
rect 25513 15385 25547 15419
rect 27261 15385 27295 15419
rect 1593 15317 1627 15351
rect 4997 15317 5031 15351
rect 7389 15317 7423 15351
rect 8217 15317 8251 15351
rect 8677 15317 8711 15351
rect 10517 15317 10551 15351
rect 11345 15317 11379 15351
rect 11621 15317 11655 15351
rect 12081 15317 12115 15351
rect 12449 15317 12483 15351
rect 19257 15317 19291 15351
rect 19441 15317 19475 15351
rect 22293 15317 22327 15351
rect 26065 15317 26099 15351
rect 27077 15317 27111 15351
rect 30205 15317 30239 15351
rect 3801 15113 3835 15147
rect 5733 15113 5767 15147
rect 13461 15113 13495 15147
rect 15025 15113 15059 15147
rect 15945 15113 15979 15147
rect 18981 15113 19015 15147
rect 19809 15113 19843 15147
rect 21189 15113 21223 15147
rect 22937 15113 22971 15147
rect 23765 15113 23799 15147
rect 26617 15113 26651 15147
rect 27629 15113 27663 15147
rect 28365 15113 28399 15147
rect 28733 15113 28767 15147
rect 29837 15113 29871 15147
rect 1685 15045 1719 15079
rect 4445 15045 4479 15079
rect 7297 15045 7331 15079
rect 9873 15045 9907 15079
rect 12265 15045 12299 15079
rect 16865 15045 16899 15079
rect 18153 15045 18187 15079
rect 22109 15045 22143 15079
rect 25605 15045 25639 15079
rect 30297 15045 30331 15079
rect 1409 14977 1443 15011
rect 4813 14977 4847 15011
rect 5549 14977 5583 15011
rect 9045 14977 9079 15011
rect 11621 14977 11655 15011
rect 11805 14977 11839 15011
rect 13093 14977 13127 15011
rect 14933 14977 14967 15011
rect 15209 14977 15243 15011
rect 15393 14977 15427 15011
rect 16313 14977 16347 15011
rect 17141 14977 17175 15011
rect 17325 14977 17359 15011
rect 18061 14977 18095 15011
rect 18245 14977 18279 15011
rect 18521 14977 18555 15011
rect 19165 14977 19199 15011
rect 19349 14977 19383 15011
rect 20453 14977 20487 15011
rect 20821 14977 20855 15011
rect 23305 14977 23339 15011
rect 25237 14977 25271 15011
rect 25329 14977 25363 15011
rect 25513 14977 25547 15011
rect 25697 14977 25731 15011
rect 25973 14977 26007 15011
rect 26065 14977 26099 15011
rect 26249 14977 26283 15011
rect 26341 14977 26375 15011
rect 26433 14977 26467 15011
rect 27813 14977 27847 15011
rect 27905 14977 27939 15011
rect 28089 14977 28123 15011
rect 28181 14977 28215 15011
rect 28273 14977 28307 15011
rect 28549 14977 28583 15011
rect 30021 14977 30055 15011
rect 3157 14909 3191 14943
rect 4905 14909 4939 14943
rect 7021 14909 7055 14943
rect 8769 14909 8803 14943
rect 11253 14909 11287 14943
rect 13185 14909 13219 14943
rect 17049 14909 17083 14943
rect 17509 14909 17543 14943
rect 17693 14909 17727 14943
rect 18613 14909 18647 14943
rect 18705 14909 18739 14943
rect 18797 14909 18831 14943
rect 19165 14841 19199 14875
rect 21557 14841 21591 14875
rect 25881 14841 25915 14875
rect 4077 14773 4111 14807
rect 5181 14773 5215 14807
rect 11621 14773 11655 14807
rect 15301 14773 15335 14807
rect 16221 14773 16255 14807
rect 20085 14773 20119 14807
rect 31769 14773 31803 14807
rect 3617 14569 3651 14603
rect 4629 14569 4663 14603
rect 8309 14569 8343 14603
rect 10885 14569 10919 14603
rect 15669 14569 15703 14603
rect 16129 14569 16163 14603
rect 16681 14569 16715 14603
rect 17693 14569 17727 14603
rect 18153 14569 18187 14603
rect 19625 14569 19659 14603
rect 21005 14569 21039 14603
rect 25237 14569 25271 14603
rect 25421 14569 25455 14603
rect 30665 14569 30699 14603
rect 30941 14569 30975 14603
rect 19809 14501 19843 14535
rect 20913 14501 20947 14535
rect 21465 14501 21499 14535
rect 27537 14501 27571 14535
rect 1869 14433 1903 14467
rect 4261 14433 4295 14467
rect 6469 14433 6503 14467
rect 9689 14433 9723 14467
rect 15577 14433 15611 14467
rect 16221 14433 16255 14467
rect 18429 14433 18463 14467
rect 18889 14433 18923 14467
rect 22017 14433 22051 14467
rect 22477 14433 22511 14467
rect 23213 14433 23247 14467
rect 24869 14433 24903 14467
rect 27169 14433 27203 14467
rect 34069 14433 34103 14467
rect 3985 14365 4019 14399
rect 6193 14365 6227 14399
rect 10977 14365 11011 14399
rect 11161 14365 11195 14399
rect 11621 14365 11655 14399
rect 12081 14365 12115 14399
rect 14939 14365 14973 14399
rect 15117 14365 15151 14399
rect 15663 14365 15697 14399
rect 15853 14365 15887 14399
rect 16681 14365 16715 14399
rect 16773 14365 16807 14399
rect 17969 14365 18003 14399
rect 18153 14365 18187 14399
rect 18337 14365 18371 14399
rect 18521 14365 18555 14399
rect 19257 14365 19291 14399
rect 19993 14365 20027 14399
rect 20177 14365 20211 14399
rect 20269 14365 20303 14399
rect 20361 14365 20395 14399
rect 20545 14365 20579 14399
rect 20729 14365 20763 14399
rect 20821 14365 20855 14399
rect 21741 14365 21775 14399
rect 21833 14365 21867 14399
rect 22385 14365 22419 14399
rect 23397 14365 23431 14399
rect 23489 14365 23523 14399
rect 23673 14365 23707 14399
rect 23765 14365 23799 14399
rect 25605 14365 25639 14399
rect 26065 14365 26099 14399
rect 26341 14365 26375 14399
rect 26801 14365 26835 14399
rect 30849 14365 30883 14399
rect 34529 14365 34563 14399
rect 2145 14297 2179 14331
rect 3893 14297 3927 14331
rect 8953 14297 8987 14331
rect 11345 14297 11379 14331
rect 16313 14297 16347 14331
rect 16957 14297 16991 14331
rect 19625 14297 19659 14331
rect 21097 14297 21131 14331
rect 7941 14229 7975 14263
rect 10517 14229 10551 14263
rect 15025 14229 15059 14263
rect 15301 14229 15335 14263
rect 15945 14229 15979 14263
rect 16497 14229 16531 14263
rect 17325 14229 17359 14263
rect 21649 14229 21683 14263
rect 23949 14229 23983 14263
rect 25237 14229 25271 14263
rect 2329 14025 2363 14059
rect 9045 14025 9079 14059
rect 11069 14025 11103 14059
rect 16313 14025 16347 14059
rect 16773 14025 16807 14059
rect 16957 14025 16991 14059
rect 17601 14025 17635 14059
rect 18061 14025 18095 14059
rect 19809 14025 19843 14059
rect 19993 14025 20027 14059
rect 20085 14025 20119 14059
rect 20821 14025 20855 14059
rect 22201 14025 22235 14059
rect 22293 14025 22327 14059
rect 22477 14025 22511 14059
rect 23121 14025 23155 14059
rect 24869 14025 24903 14059
rect 25529 14025 25563 14059
rect 25697 14025 25731 14059
rect 31953 14025 31987 14059
rect 34897 14025 34931 14059
rect 6653 13957 6687 13991
rect 8309 13957 8343 13991
rect 18337 13957 18371 13991
rect 19349 13957 19383 13991
rect 20729 13957 20763 13991
rect 21557 13957 21591 13991
rect 22109 13957 22143 13991
rect 24133 13957 24167 13991
rect 25329 13957 25363 13991
rect 2237 13889 2271 13923
rect 3985 13889 4019 13923
rect 6377 13889 6411 13923
rect 8401 13889 8435 13923
rect 10149 13889 10183 13923
rect 11805 13889 11839 13923
rect 12081 13889 12115 13923
rect 13001 13889 13035 13923
rect 14657 13889 14691 13923
rect 14841 13889 14875 13923
rect 14933 13889 14967 13923
rect 16129 13889 16163 13923
rect 16405 13889 16439 13923
rect 16681 13889 16715 13923
rect 17049 13889 17083 13923
rect 19441 13889 19475 13923
rect 21281 13889 21315 13923
rect 23765 13889 23799 13923
rect 23949 13889 23983 13923
rect 24685 13889 24719 13923
rect 28365 13889 28399 13923
rect 31585 13889 31619 13923
rect 32321 13889 32355 13923
rect 4077 13821 4111 13855
rect 8125 13821 8159 13855
rect 10701 13821 10735 13855
rect 12633 13821 12667 13855
rect 13093 13821 13127 13855
rect 16865 13821 16899 13855
rect 18797 13821 18831 13855
rect 20269 13821 20303 13855
rect 20361 13821 20395 13855
rect 22753 13821 22787 13855
rect 24501 13821 24535 13855
rect 28273 13821 28307 13855
rect 28733 13821 28767 13855
rect 31677 13821 31711 13855
rect 32229 13821 32263 13855
rect 32965 13821 32999 13855
rect 33149 13821 33183 13855
rect 33425 13821 33459 13855
rect 4353 13753 4387 13787
rect 13369 13753 13403 13787
rect 20913 13753 20947 13787
rect 21925 13753 21959 13787
rect 32689 13753 32723 13787
rect 2789 13685 2823 13719
rect 4813 13685 4847 13719
rect 8769 13685 8803 13719
rect 14749 13685 14783 13719
rect 16129 13685 16163 13719
rect 19809 13685 19843 13719
rect 23489 13685 23523 13719
rect 25513 13685 25547 13719
rect 31677 13685 31711 13719
rect 4261 13481 4295 13515
rect 14841 13481 14875 13515
rect 15761 13481 15795 13515
rect 16405 13481 16439 13515
rect 16589 13481 16623 13515
rect 18153 13481 18187 13515
rect 18889 13481 18923 13515
rect 19533 13481 19567 13515
rect 20545 13481 20579 13515
rect 21281 13481 21315 13515
rect 21649 13481 21683 13515
rect 23029 13481 23063 13515
rect 23673 13481 23707 13515
rect 27261 13481 27295 13515
rect 28549 13481 28583 13515
rect 31493 13481 31527 13515
rect 31953 13481 31987 13515
rect 34161 13481 34195 13515
rect 22201 13413 22235 13447
rect 31861 13413 31895 13447
rect 1409 13345 1443 13379
rect 4537 13345 4571 13379
rect 4629 13345 4663 13379
rect 5641 13345 5675 13379
rect 5825 13345 5859 13379
rect 6285 13345 6319 13379
rect 9229 13345 9263 13379
rect 10701 13345 10735 13379
rect 11897 13345 11931 13379
rect 17049 13345 17083 13379
rect 21833 13345 21867 13379
rect 29101 13345 29135 13379
rect 32045 13345 32079 13379
rect 32321 13345 32355 13379
rect 4445 13277 4479 13311
rect 4721 13277 4755 13311
rect 4905 13277 4939 13311
rect 4997 13277 5031 13311
rect 5181 13277 5215 13311
rect 5273 13277 5307 13311
rect 5365 13277 5399 13311
rect 5917 13277 5951 13311
rect 8953 13277 8987 13311
rect 10885 13277 10919 13311
rect 11437 13277 11471 13311
rect 12265 13277 12299 13311
rect 12357 13277 12391 13311
rect 12541 13277 12575 13311
rect 14565 13277 14599 13311
rect 14703 13277 14737 13311
rect 15025 13277 15059 13311
rect 15209 13277 15243 13311
rect 15301 13277 15335 13311
rect 15485 13277 15519 13311
rect 15577 13277 15611 13311
rect 16589 13277 16623 13311
rect 16773 13277 16807 13311
rect 16861 13277 16895 13311
rect 16957 13277 16991 13311
rect 17141 13277 17175 13311
rect 18337 13277 18371 13311
rect 18613 13277 18647 13311
rect 18705 13277 18739 13311
rect 19901 13277 19935 13311
rect 20913 13277 20947 13311
rect 22017 13277 22051 13311
rect 27445 13277 27479 13311
rect 27537 13277 27571 13311
rect 27721 13277 27755 13311
rect 27813 13277 27847 13311
rect 28089 13277 28123 13311
rect 28181 13277 28215 13311
rect 28273 13277 28307 13311
rect 28365 13277 28399 13311
rect 29009 13277 29043 13311
rect 29745 13277 29779 13311
rect 31769 13277 31803 13311
rect 34069 13277 34103 13311
rect 1685 13209 1719 13243
rect 4077 13209 4111 13243
rect 14933 13209 14967 13243
rect 18521 13209 18555 13243
rect 20269 13209 20303 13243
rect 24041 13209 24075 13243
rect 30021 13209 30055 13243
rect 3157 13141 3191 13175
rect 3525 13141 3559 13175
rect 13093 13141 13127 13175
rect 17601 13141 17635 13175
rect 22569 13141 22603 13175
rect 23305 13141 23339 13175
rect 29377 13141 29411 13175
rect 33977 13141 34011 13175
rect 1593 12937 1627 12971
rect 2421 12937 2455 12971
rect 2881 12937 2915 12971
rect 3525 12937 3559 12971
rect 3893 12937 3927 12971
rect 6535 12937 6569 12971
rect 8861 12937 8895 12971
rect 9137 12937 9171 12971
rect 9413 12937 9447 12971
rect 14381 12937 14415 12971
rect 15117 12937 15151 12971
rect 15945 12937 15979 12971
rect 16313 12937 16347 12971
rect 17693 12937 17727 12971
rect 19165 12937 19199 12971
rect 19349 12937 19383 12971
rect 20085 12937 20119 12971
rect 20269 12937 20303 12971
rect 21465 12937 21499 12971
rect 22753 12937 22787 12971
rect 23305 12937 23339 12971
rect 27997 12937 28031 12971
rect 28641 12937 28675 12971
rect 29561 12937 29595 12971
rect 30573 12937 30607 12971
rect 30757 12937 30791 12971
rect 31585 12937 31619 12971
rect 4077 12869 4111 12903
rect 5457 12869 5491 12903
rect 6745 12869 6779 12903
rect 7389 12869 7423 12903
rect 10517 12869 10551 12903
rect 11345 12869 11379 12903
rect 13803 12869 13837 12903
rect 19717 12869 19751 12903
rect 21005 12869 21039 12903
rect 23121 12869 23155 12903
rect 27629 12869 27663 12903
rect 27829 12869 27863 12903
rect 1409 12801 1443 12835
rect 2513 12801 2547 12835
rect 4261 12801 4295 12835
rect 4353 12801 4387 12835
rect 5825 12801 5859 12835
rect 9321 12801 9355 12835
rect 10149 12801 10183 12835
rect 11621 12801 11655 12835
rect 11897 12801 11931 12835
rect 12449 12801 12483 12835
rect 13645 12801 13679 12835
rect 13921 12801 13955 12835
rect 14013 12801 14047 12835
rect 14105 12801 14139 12835
rect 14289 12801 14323 12835
rect 14749 12801 14783 12835
rect 15025 12801 15059 12835
rect 15209 12801 15243 12835
rect 16129 12801 16163 12835
rect 16405 12801 16439 12835
rect 17049 12801 17083 12835
rect 17325 12801 17359 12835
rect 17877 12801 17911 12835
rect 18061 12801 18095 12835
rect 18521 12801 18555 12835
rect 18613 12801 18647 12835
rect 18797 12801 18831 12835
rect 18889 12801 18923 12835
rect 19257 12801 19291 12835
rect 19901 12801 19935 12835
rect 19993 12801 20027 12835
rect 22017 12801 22051 12835
rect 22201 12801 22235 12835
rect 23213 12801 23247 12835
rect 23857 12801 23891 12835
rect 24133 12801 24167 12835
rect 24501 12801 24535 12835
rect 25053 12801 25087 12835
rect 25237 12801 25271 12835
rect 25605 12801 25639 12835
rect 26157 12801 26191 12835
rect 27169 12801 27203 12835
rect 27261 12801 27295 12835
rect 27353 12801 27387 12835
rect 28273 12801 28307 12835
rect 30665 12801 30699 12835
rect 31769 12801 31803 12835
rect 31953 12801 31987 12835
rect 32321 12801 32355 12835
rect 5917 12733 5951 12767
rect 6193 12733 6227 12767
rect 7113 12733 7147 12767
rect 11989 12733 12023 12767
rect 12541 12733 12575 12767
rect 13185 12733 13219 12767
rect 14565 12733 14599 12767
rect 14657 12733 14691 12767
rect 14841 12733 14875 12767
rect 18245 12733 18279 12767
rect 18981 12733 19015 12767
rect 20545 12733 20579 12767
rect 21925 12733 21959 12767
rect 22109 12733 22143 12767
rect 22385 12733 22419 12767
rect 25145 12733 25179 12767
rect 26065 12733 26099 12767
rect 26525 12733 26559 12767
rect 27077 12733 27111 12767
rect 27537 12733 27571 12767
rect 28365 12733 28399 12767
rect 31861 12733 31895 12767
rect 32229 12733 32263 12767
rect 4537 12665 4571 12699
rect 6377 12665 6411 12699
rect 19533 12665 19567 12699
rect 22937 12665 22971 12699
rect 32689 12665 32723 12699
rect 4169 12597 4203 12631
rect 6561 12597 6595 12631
rect 9873 12597 9907 12631
rect 16129 12597 16163 12631
rect 18337 12597 18371 12631
rect 23489 12597 23523 12631
rect 27813 12597 27847 12631
rect 28457 12597 28491 12631
rect 34621 12597 34655 12631
rect 3157 12393 3191 12427
rect 8217 12393 8251 12427
rect 8677 12393 8711 12427
rect 11529 12393 11563 12427
rect 14105 12393 14139 12427
rect 16405 12393 16439 12427
rect 17509 12393 17543 12427
rect 18153 12393 18187 12427
rect 20085 12393 20119 12427
rect 20269 12393 20303 12427
rect 22293 12393 22327 12427
rect 25053 12393 25087 12427
rect 27261 12393 27295 12427
rect 4261 12325 4295 12359
rect 22753 12325 22787 12359
rect 24593 12325 24627 12359
rect 25605 12325 25639 12359
rect 1409 12257 1443 12291
rect 14933 12257 14967 12291
rect 15577 12257 15611 12291
rect 15669 12257 15703 12291
rect 19809 12257 19843 12291
rect 26341 12257 26375 12291
rect 29837 12257 29871 12291
rect 33057 12257 33091 12291
rect 3433 12189 3467 12223
rect 3985 12189 4019 12223
rect 6285 12189 6319 12223
rect 7021 12189 7055 12223
rect 8125 12189 8159 12223
rect 12449 12189 12483 12223
rect 12633 12189 12667 12223
rect 14289 12189 14323 12223
rect 14565 12189 14599 12223
rect 15071 12189 15105 12223
rect 15301 12189 15335 12223
rect 15393 12189 15427 12223
rect 16037 12189 16071 12223
rect 16592 12167 16626 12201
rect 16681 12189 16715 12223
rect 16865 12189 16899 12223
rect 16957 12189 16991 12223
rect 17049 12189 17083 12223
rect 17325 12189 17359 12223
rect 17877 12189 17911 12223
rect 18613 12189 18647 12223
rect 18705 12189 18739 12223
rect 18797 12189 18831 12223
rect 18981 12189 19015 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 19993 12189 20027 12223
rect 20269 12189 20303 12223
rect 20361 12189 20395 12223
rect 21097 12189 21131 12223
rect 21189 12189 21223 12223
rect 21465 12189 21499 12223
rect 21649 12189 21683 12223
rect 21833 12189 21867 12223
rect 21925 12189 21959 12223
rect 22569 12189 22603 12223
rect 22753 12189 22787 12223
rect 23029 12189 23063 12223
rect 23213 12189 23247 12223
rect 23397 12189 23431 12223
rect 23489 12189 23523 12223
rect 23581 12189 23615 12223
rect 24133 12189 24167 12223
rect 25789 12189 25823 12223
rect 25895 12189 25929 12223
rect 26065 12189 26099 12223
rect 26157 12189 26191 12223
rect 26709 12189 26743 12223
rect 26893 12189 26927 12223
rect 27077 12189 27111 12223
rect 27353 12189 27387 12223
rect 29561 12189 29595 12223
rect 32689 12189 32723 12223
rect 32781 12189 32815 12223
rect 34713 12189 34747 12223
rect 1685 12121 1719 12155
rect 3341 12121 3375 12155
rect 15209 12121 15243 12155
rect 15853 12121 15887 12155
rect 17141 12121 17175 12155
rect 23121 12121 23155 12155
rect 25145 12121 25179 12155
rect 25329 12121 25363 12155
rect 26985 12121 27019 12155
rect 29377 12121 29411 12155
rect 34805 12121 34839 12155
rect 3893 12053 3927 12087
rect 6469 12053 6503 12087
rect 7205 12053 7239 12087
rect 14473 12053 14507 12087
rect 18337 12053 18371 12087
rect 20637 12053 20671 12087
rect 20729 12053 20763 12087
rect 21373 12053 21407 12087
rect 22845 12053 22879 12087
rect 23765 12053 23799 12087
rect 23857 12053 23891 12087
rect 23949 12053 23983 12087
rect 27445 12053 27479 12087
rect 31309 12053 31343 12087
rect 34529 12053 34563 12087
rect 4261 11849 4295 11883
rect 13093 11849 13127 11883
rect 13369 11849 13403 11883
rect 13921 11849 13955 11883
rect 17141 11849 17175 11883
rect 17785 11849 17819 11883
rect 19349 11849 19383 11883
rect 21833 11849 21867 11883
rect 22201 11849 22235 11883
rect 22293 11849 22327 11883
rect 23305 11849 23339 11883
rect 24685 11849 24719 11883
rect 25421 11849 25455 11883
rect 26433 11849 26467 11883
rect 27629 11849 27663 11883
rect 28365 11849 28399 11883
rect 30941 11849 30975 11883
rect 32321 11849 32355 11883
rect 7941 11781 7975 11815
rect 9597 11781 9631 11815
rect 10793 11781 10827 11815
rect 16681 11781 16715 11815
rect 17325 11781 17359 11815
rect 21189 11781 21223 11815
rect 21373 11781 21407 11815
rect 22845 11781 22879 11815
rect 25053 11781 25087 11815
rect 30665 11781 30699 11815
rect 2513 11713 2547 11747
rect 9689 11713 9723 11747
rect 10241 11713 10275 11747
rect 13553 11713 13587 11747
rect 13737 11713 13771 11747
rect 16037 11713 16071 11747
rect 16313 11713 16347 11747
rect 16497 11713 16531 11747
rect 16957 11713 16991 11747
rect 17233 11713 17267 11747
rect 17417 11713 17451 11747
rect 18429 11713 18463 11747
rect 18613 11713 18647 11747
rect 20729 11713 20763 11747
rect 21097 11713 21131 11747
rect 22661 11713 22695 11747
rect 22937 11703 22971 11737
rect 24041 11713 24075 11747
rect 24317 11713 24351 11747
rect 26341 11713 26375 11747
rect 26985 11713 27019 11747
rect 27169 11713 27203 11747
rect 27261 11713 27295 11747
rect 27353 11713 27387 11747
rect 27721 11713 27755 11747
rect 27814 11713 27848 11747
rect 27997 11713 28031 11747
rect 28089 11713 28123 11747
rect 28186 11713 28220 11747
rect 28733 11713 28767 11747
rect 30757 11713 30791 11747
rect 31033 11713 31067 11747
rect 31401 11713 31435 11747
rect 31677 11713 31711 11747
rect 34713 11713 34747 11747
rect 2789 11645 2823 11679
rect 4629 11645 4663 11679
rect 7665 11645 7699 11679
rect 9413 11645 9447 11679
rect 16773 11645 16807 11679
rect 18797 11645 18831 11679
rect 22477 11645 22511 11679
rect 26709 11645 26743 11679
rect 29009 11645 29043 11679
rect 31769 11645 31803 11679
rect 31953 11645 31987 11679
rect 34437 11645 34471 11679
rect 16175 11577 16209 11611
rect 16405 11577 16439 11611
rect 19993 11577 20027 11611
rect 21373 11577 21407 11611
rect 10057 11509 10091 11543
rect 16681 11509 16715 11543
rect 18337 11509 18371 11543
rect 19625 11509 19659 11543
rect 20361 11509 20395 11543
rect 22661 11509 22695 11543
rect 23581 11509 23615 11543
rect 26617 11509 26651 11543
rect 26801 11509 26835 11543
rect 30481 11509 30515 11543
rect 31861 11509 31895 11543
rect 1593 11305 1627 11339
rect 18153 11305 18187 11339
rect 18521 11305 18555 11339
rect 20177 11305 20211 11339
rect 21005 11305 21039 11339
rect 22293 11305 22327 11339
rect 22661 11305 22695 11339
rect 24225 11305 24259 11339
rect 27813 11305 27847 11339
rect 28641 11305 28675 11339
rect 31493 11305 31527 11339
rect 31769 11305 31803 11339
rect 18889 11237 18923 11271
rect 21373 11237 21407 11271
rect 21741 11237 21775 11271
rect 25881 11237 25915 11271
rect 32413 11237 32447 11271
rect 23397 11169 23431 11203
rect 23581 11169 23615 11203
rect 31401 11169 31435 11203
rect 31953 11169 31987 11203
rect 33057 11169 33091 11203
rect 34529 11169 34563 11203
rect 1409 11101 1443 11135
rect 22109 11101 22143 11135
rect 22293 11101 22327 11135
rect 23029 11101 23063 11135
rect 23213 11101 23247 11135
rect 23489 11101 23523 11135
rect 23949 11101 23983 11135
rect 24409 11101 24443 11135
rect 24777 11101 24811 11135
rect 25145 11101 25179 11135
rect 25513 11101 25547 11135
rect 25973 11101 26007 11135
rect 26893 11101 26927 11135
rect 27077 11101 27111 11135
rect 27261 11101 27295 11135
rect 27445 11101 27479 11135
rect 27629 11101 27663 11135
rect 31585 11101 31619 11135
rect 32045 11101 32079 11135
rect 32781 11101 32815 11135
rect 34713 11101 34747 11135
rect 9597 11033 9631 11067
rect 20453 11033 20487 11067
rect 23765 11033 23799 11067
rect 23857 11033 23891 11067
rect 26985 11033 27019 11067
rect 27537 11033 27571 11067
rect 30389 11033 30423 11067
rect 31309 11033 31343 11067
rect 34805 11033 34839 11067
rect 10609 10761 10643 10795
rect 23581 10761 23615 10795
rect 27445 10761 27479 10795
rect 29377 10761 29411 10795
rect 31309 10761 31343 10795
rect 32689 10761 32723 10795
rect 32965 10761 32999 10795
rect 25881 10693 25915 10727
rect 9321 10625 9355 10659
rect 18705 10625 18739 10659
rect 19257 10625 19291 10659
rect 20453 10625 20487 10659
rect 20637 10625 20671 10659
rect 20729 10625 20763 10659
rect 20913 10625 20947 10659
rect 21373 10625 21407 10659
rect 22109 10625 22143 10659
rect 22293 10625 22327 10659
rect 22569 10625 22603 10659
rect 23029 10625 23063 10659
rect 23213 10625 23247 10659
rect 24685 10625 24719 10659
rect 24869 10625 24903 10659
rect 24961 10625 24995 10659
rect 25605 10625 25639 10659
rect 25789 10625 25823 10659
rect 25973 10625 26007 10659
rect 26249 10625 26283 10659
rect 26433 10625 26467 10659
rect 27169 10625 27203 10659
rect 29837 10625 29871 10659
rect 30021 10625 30055 10659
rect 31585 10625 31619 10659
rect 31769 10625 31803 10659
rect 31861 10625 31895 10659
rect 21189 10557 21223 10591
rect 22661 10557 22695 10591
rect 23121 10557 23155 10591
rect 23857 10557 23891 10591
rect 24225 10557 24259 10591
rect 25237 10557 25271 10591
rect 27077 10557 27111 10591
rect 27261 10557 27295 10591
rect 11805 10489 11839 10523
rect 21557 10489 21591 10523
rect 22937 10489 22971 10523
rect 25513 10489 25547 10523
rect 26157 10489 26191 10523
rect 26341 10489 26375 10523
rect 31677 10489 31711 10523
rect 20545 10421 20579 10455
rect 20821 10421 20855 10455
rect 22201 10421 22235 10455
rect 22569 10421 22603 10455
rect 24869 10421 24903 10455
rect 25053 10421 25087 10455
rect 30113 10421 30147 10455
rect 31401 10421 31435 10455
rect 34161 10421 34195 10455
rect 34529 10421 34563 10455
rect 4077 10217 4111 10251
rect 18705 10217 18739 10251
rect 19533 10217 19567 10251
rect 19993 10217 20027 10251
rect 21281 10217 21315 10251
rect 22017 10217 22051 10251
rect 22845 10217 22879 10251
rect 23213 10217 23247 10251
rect 23673 10217 23707 10251
rect 24593 10217 24627 10251
rect 24777 10217 24811 10251
rect 29009 10217 29043 10251
rect 31309 10217 31343 10251
rect 32505 10217 32539 10251
rect 20913 10149 20947 10183
rect 1593 10081 1627 10115
rect 18153 10081 18187 10115
rect 20637 10081 20671 10115
rect 22569 10081 22603 10115
rect 28089 10081 28123 10115
rect 31493 10081 31527 10115
rect 31953 10081 31987 10115
rect 33057 10081 33091 10115
rect 3617 10013 3651 10047
rect 18613 10013 18647 10047
rect 18797 10013 18831 10047
rect 19441 10013 19475 10047
rect 19625 10013 19659 10047
rect 20545 10013 20579 10047
rect 22201 10013 22235 10047
rect 22477 10013 22511 10047
rect 23857 10013 23891 10047
rect 24133 10013 24167 10047
rect 24225 10013 24259 10047
rect 26525 10013 26559 10047
rect 26985 10013 27019 10047
rect 28181 10013 28215 10047
rect 29193 10013 29227 10047
rect 29561 10013 29595 10047
rect 31585 10013 31619 10047
rect 32045 10013 32079 10047
rect 32229 10013 32263 10047
rect 32781 10013 32815 10047
rect 34713 10013 34747 10047
rect 1869 9945 1903 9979
rect 18521 9945 18555 9979
rect 24409 9945 24443 9979
rect 24609 9945 24643 9979
rect 29837 9945 29871 9979
rect 34805 9945 34839 9979
rect 21557 9877 21591 9911
rect 25053 9877 25087 9911
rect 25421 9877 25455 9911
rect 28549 9877 28583 9911
rect 29285 9877 29319 9911
rect 32229 9877 32263 9911
rect 34529 9877 34563 9911
rect 3249 9673 3283 9707
rect 23121 9673 23155 9707
rect 24041 9673 24075 9707
rect 24409 9673 24443 9707
rect 2789 9605 2823 9639
rect 18337 9605 18371 9639
rect 22385 9605 22419 9639
rect 22845 9605 22879 9639
rect 27445 9605 27479 9639
rect 28825 9605 28859 9639
rect 2881 9537 2915 9571
rect 23397 9537 23431 9571
rect 23673 9537 23707 9571
rect 24777 9537 24811 9571
rect 27353 9537 27387 9571
rect 27537 9537 27571 9571
rect 32321 9537 32355 9571
rect 32781 9537 32815 9571
rect 34713 9537 34747 9571
rect 22109 9469 22143 9503
rect 28457 9469 28491 9503
rect 28549 9469 28583 9503
rect 30297 9469 30331 9503
rect 32229 9469 32263 9503
rect 34437 9469 34471 9503
rect 23489 9333 23523 9367
rect 32597 9333 32631 9367
rect 32965 9333 32999 9367
rect 1593 9129 1627 9163
rect 23029 9129 23063 9163
rect 23489 9129 23523 9163
rect 27721 9061 27755 9095
rect 1409 8925 1443 8959
rect 24501 8925 24535 8959
rect 25053 8925 25087 8959
rect 26433 8925 26467 8959
rect 28457 8925 28491 8959
rect 32873 8925 32907 8959
rect 33425 8925 33459 8959
rect 33885 8925 33919 8959
rect 33057 8789 33091 8823
rect 33517 8789 33551 8823
rect 27169 8517 27203 8551
rect 32413 8517 32447 8551
rect 32781 8517 32815 8551
rect 27813 8449 27847 8483
rect 32505 8449 32539 8483
rect 34529 8449 34563 8483
rect 34805 8449 34839 8483
rect 34253 8313 34287 8347
rect 34437 8245 34471 8279
rect 32689 8041 32723 8075
rect 32781 7905 32815 7939
rect 33057 7905 33091 7939
rect 34529 7701 34563 7735
rect 34713 7361 34747 7395
rect 34437 7293 34471 7327
rect 1409 6749 1443 6783
rect 1593 6613 1627 6647
rect 34069 5729 34103 5763
rect 34345 5661 34379 5695
rect 1593 4777 1627 4811
rect 1409 4573 1443 4607
rect 34069 3553 34103 3587
rect 34437 3485 34471 3519
rect 1593 2601 1627 2635
rect 27537 2601 27571 2635
rect 9597 2465 9631 2499
rect 1409 2397 1443 2431
rect 9137 2397 9171 2431
rect 27353 2397 27387 2431
<< metal1 >>
rect 1104 36474 35248 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 35248 36474
rect 1104 36400 35248 36422
rect 934 36116 940 36168
rect 992 36156 998 36168
rect 1397 36159 1455 36165
rect 1397 36156 1409 36159
rect 992 36128 1409 36156
rect 992 36116 998 36128
rect 1397 36125 1409 36128
rect 1443 36125 1455 36159
rect 1397 36119 1455 36125
rect 33134 36116 33140 36168
rect 33192 36116 33198 36168
rect 34330 36048 34336 36100
rect 34388 36048 34394 36100
rect 1578 35980 1584 36032
rect 1636 35980 1642 36032
rect 1104 35930 35236 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 35236 35930
rect 1104 35856 35236 35878
rect 1104 35386 35248 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 35248 35386
rect 1104 35312 35248 35334
rect 934 35028 940 35080
rect 992 35068 998 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 992 35040 1409 35068
rect 992 35028 998 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 1854 34932 1860 34944
rect 1627 34904 1860 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 1854 34892 1860 34904
rect 1912 34892 1918 34944
rect 1104 34842 35236 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 35236 34842
rect 1104 34768 35236 34790
rect 1104 34298 35248 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 35248 34298
rect 1104 34224 35248 34246
rect 34057 34051 34115 34057
rect 34057 34017 34069 34051
rect 34103 34048 34115 34051
rect 34103 34020 34652 34048
rect 34103 34017 34115 34020
rect 34057 34011 34115 34017
rect 34514 33940 34520 33992
rect 34572 33940 34578 33992
rect 34624 33924 34652 34020
rect 34606 33872 34612 33924
rect 34664 33872 34670 33924
rect 1104 33754 35236 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 35236 33754
rect 1104 33680 35236 33702
rect 1104 33210 35248 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 35248 33210
rect 1104 33136 35248 33158
rect 934 32852 940 32904
rect 992 32892 998 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 992 32864 1409 32892
rect 992 32852 998 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32756 1639 32759
rect 4062 32756 4068 32768
rect 1627 32728 4068 32756
rect 1627 32725 1639 32728
rect 1581 32719 1639 32725
rect 4062 32716 4068 32728
rect 4120 32716 4126 32768
rect 1104 32666 35236 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 35236 32666
rect 1104 32592 35236 32614
rect 1104 32122 35248 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 35248 32122
rect 1104 32048 35248 32070
rect 34057 31875 34115 31881
rect 34057 31841 34069 31875
rect 34103 31841 34115 31875
rect 34057 31835 34115 31841
rect 34072 31748 34100 31835
rect 34422 31764 34428 31816
rect 34480 31764 34486 31816
rect 34054 31696 34060 31748
rect 34112 31696 34118 31748
rect 1104 31578 35236 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 35236 31578
rect 1104 31504 35236 31526
rect 1104 31034 35248 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 35248 31034
rect 1104 30960 35248 30982
rect 1394 30676 1400 30728
rect 1452 30676 1458 30728
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 2866 30580 2872 30592
rect 1627 30552 2872 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 2866 30540 2872 30552
rect 2924 30540 2930 30592
rect 1104 30490 35236 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 35236 30490
rect 1104 30416 35236 30438
rect 1104 29946 35248 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 35248 29946
rect 1104 29872 35248 29894
rect 34057 29699 34115 29705
rect 34057 29665 34069 29699
rect 34103 29696 34115 29699
rect 34103 29668 34652 29696
rect 34103 29665 34115 29668
rect 34057 29659 34115 29665
rect 34517 29631 34575 29637
rect 34517 29597 34529 29631
rect 34563 29597 34575 29631
rect 34517 29591 34575 29597
rect 34532 29492 34560 29591
rect 34624 29572 34652 29668
rect 34606 29520 34612 29572
rect 34664 29520 34670 29572
rect 34790 29492 34796 29504
rect 34532 29464 34796 29492
rect 34790 29452 34796 29464
rect 34848 29452 34854 29504
rect 1104 29402 35236 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 35236 29402
rect 1104 29328 35236 29350
rect 1104 28858 35248 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 35248 28858
rect 1104 28784 35248 28806
rect 34514 28704 34520 28756
rect 34572 28704 34578 28756
rect 19444 28648 20392 28676
rect 934 28500 940 28552
rect 992 28540 998 28552
rect 19444 28549 19472 28648
rect 1397 28543 1455 28549
rect 1397 28540 1409 28543
rect 992 28512 1409 28540
rect 992 28500 998 28512
rect 1397 28509 1409 28512
rect 1443 28509 1455 28543
rect 1397 28503 1455 28509
rect 19429 28543 19487 28549
rect 19429 28509 19441 28543
rect 19475 28509 19487 28543
rect 19429 28503 19487 28509
rect 19613 28543 19671 28549
rect 19613 28509 19625 28543
rect 19659 28540 19671 28543
rect 19889 28543 19947 28549
rect 19889 28540 19901 28543
rect 19659 28512 19901 28540
rect 19659 28509 19671 28512
rect 19613 28503 19671 28509
rect 19889 28509 19901 28512
rect 19935 28540 19947 28543
rect 19978 28540 19984 28552
rect 19935 28512 19984 28540
rect 19935 28509 19947 28512
rect 19889 28503 19947 28509
rect 19978 28500 19984 28512
rect 20036 28500 20042 28552
rect 20088 28549 20116 28648
rect 20364 28620 20392 28648
rect 20346 28568 20352 28620
rect 20404 28608 20410 28620
rect 21085 28611 21143 28617
rect 21085 28608 21097 28611
rect 20404 28580 21097 28608
rect 20404 28568 20410 28580
rect 21085 28577 21097 28580
rect 21131 28577 21143 28611
rect 21085 28571 21143 28577
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28509 20131 28543
rect 20073 28503 20131 28509
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28509 21235 28543
rect 32769 28543 32827 28549
rect 32769 28540 32781 28543
rect 21177 28503 21235 28509
rect 32600 28512 32781 28540
rect 19797 28475 19855 28481
rect 19797 28441 19809 28475
rect 19843 28472 19855 28475
rect 20162 28472 20168 28484
rect 19843 28444 20168 28472
rect 19843 28441 19855 28444
rect 19797 28435 19855 28441
rect 20162 28432 20168 28444
rect 20220 28432 20226 28484
rect 1578 28364 1584 28416
rect 1636 28364 1642 28416
rect 19334 28364 19340 28416
rect 19392 28404 19398 28416
rect 19886 28404 19892 28416
rect 19392 28376 19892 28404
rect 19392 28364 19398 28376
rect 19886 28364 19892 28376
rect 19944 28364 19950 28416
rect 19978 28364 19984 28416
rect 20036 28404 20042 28416
rect 21192 28404 21220 28503
rect 32600 28416 32628 28512
rect 32769 28509 32781 28512
rect 32815 28509 32827 28543
rect 32769 28503 32827 28509
rect 34146 28500 34152 28552
rect 34204 28500 34210 28552
rect 33042 28432 33048 28484
rect 33100 28432 33106 28484
rect 20036 28376 21220 28404
rect 20036 28364 20042 28376
rect 21542 28364 21548 28416
rect 21600 28364 21606 28416
rect 32582 28364 32588 28416
rect 32640 28364 32646 28416
rect 1104 28314 35236 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 35236 28314
rect 1104 28240 35236 28262
rect 19794 28200 19800 28212
rect 18984 28172 19800 28200
rect 18984 28073 19012 28172
rect 19794 28160 19800 28172
rect 19852 28160 19858 28212
rect 21450 28200 21456 28212
rect 19996 28172 21456 28200
rect 19245 28135 19303 28141
rect 19245 28101 19257 28135
rect 19291 28132 19303 28135
rect 19889 28135 19947 28141
rect 19291 28104 19840 28132
rect 19291 28101 19303 28104
rect 19245 28095 19303 28101
rect 18969 28067 19027 28073
rect 18969 28033 18981 28067
rect 19015 28033 19027 28067
rect 18969 28027 19027 28033
rect 19334 28024 19340 28076
rect 19392 28064 19398 28076
rect 19613 28067 19671 28073
rect 19613 28064 19625 28067
rect 19392 28036 19625 28064
rect 19392 28024 19398 28036
rect 19613 28033 19625 28036
rect 19659 28033 19671 28067
rect 19812 28064 19840 28104
rect 19889 28101 19901 28135
rect 19935 28132 19947 28135
rect 19996 28132 20024 28172
rect 21450 28160 21456 28172
rect 21508 28160 21514 28212
rect 21542 28160 21548 28212
rect 21600 28200 21606 28212
rect 21600 28172 22094 28200
rect 21600 28160 21606 28172
rect 19935 28104 20024 28132
rect 19935 28101 19947 28104
rect 19889 28095 19947 28101
rect 20070 28092 20076 28144
rect 20128 28132 20134 28144
rect 20993 28135 21051 28141
rect 20993 28132 21005 28135
rect 20128 28104 21005 28132
rect 20128 28092 20134 28104
rect 20364 28073 20392 28104
rect 20993 28101 21005 28104
rect 21039 28101 21051 28135
rect 20993 28095 21051 28101
rect 19981 28067 20039 28073
rect 19981 28064 19993 28067
rect 19812 28036 19993 28064
rect 19613 28027 19671 28033
rect 19981 28033 19993 28036
rect 20027 28033 20039 28067
rect 19981 28027 20039 28033
rect 20349 28067 20407 28073
rect 20349 28033 20361 28067
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 21082 28024 21088 28076
rect 21140 28024 21146 28076
rect 19245 27999 19303 28005
rect 19245 27965 19257 27999
rect 19291 27996 19303 27999
rect 19426 27996 19432 28008
rect 19291 27968 19432 27996
rect 19291 27965 19303 27968
rect 19245 27959 19303 27965
rect 19426 27956 19432 27968
rect 19484 27956 19490 28008
rect 19518 27956 19524 28008
rect 19576 27956 19582 28008
rect 19812 27968 20024 27996
rect 19061 27931 19119 27937
rect 19061 27897 19073 27931
rect 19107 27928 19119 27931
rect 19812 27928 19840 27968
rect 19107 27900 19840 27928
rect 19996 27928 20024 27968
rect 20070 27956 20076 28008
rect 20128 27956 20134 28008
rect 20162 27956 20168 28008
rect 20220 27996 20226 28008
rect 20625 27999 20683 28005
rect 20625 27996 20637 27999
rect 20220 27968 20637 27996
rect 20220 27956 20226 27968
rect 20625 27965 20637 27968
rect 20671 27965 20683 27999
rect 22066 27996 22094 28172
rect 34422 28160 34428 28212
rect 34480 28160 34486 28212
rect 31297 28135 31355 28141
rect 31297 28132 31309 28135
rect 30668 28104 31309 28132
rect 22554 28024 22560 28076
rect 22612 28024 22618 28076
rect 22465 27999 22523 28005
rect 22465 27996 22477 27999
rect 22066 27968 22477 27996
rect 20625 27959 20683 27965
rect 22465 27965 22477 27968
rect 22511 27965 22523 27999
rect 22465 27959 22523 27965
rect 20533 27931 20591 27937
rect 20533 27928 20545 27931
rect 19996 27900 20545 27928
rect 19107 27897 19119 27900
rect 19061 27891 19119 27897
rect 20533 27897 20545 27900
rect 20579 27897 20591 27931
rect 20533 27891 20591 27897
rect 30668 27872 30696 28104
rect 31036 28073 31064 28104
rect 31297 28101 31309 28104
rect 31343 28101 31355 28135
rect 31297 28095 31355 28101
rect 33686 28092 33692 28144
rect 33744 28092 33750 28144
rect 30837 28067 30895 28073
rect 30837 28033 30849 28067
rect 30883 28033 30895 28067
rect 30837 28027 30895 28033
rect 31021 28067 31079 28073
rect 31021 28033 31033 28067
rect 31067 28064 31079 28067
rect 31067 28036 31101 28064
rect 31067 28033 31079 28036
rect 31021 28027 31079 28033
rect 30852 27996 30880 28027
rect 32677 27999 32735 28005
rect 32677 27996 32689 27999
rect 30852 27968 31064 27996
rect 31036 27872 31064 27968
rect 32600 27968 32689 27996
rect 32600 27872 32628 27968
rect 32677 27965 32689 27968
rect 32723 27965 32735 27999
rect 32677 27959 32735 27965
rect 32950 27956 32956 28008
rect 33008 27956 33014 28008
rect 19334 27820 19340 27872
rect 19392 27820 19398 27872
rect 20806 27820 20812 27872
rect 20864 27820 20870 27872
rect 22830 27820 22836 27872
rect 22888 27820 22894 27872
rect 30101 27863 30159 27869
rect 30101 27829 30113 27863
rect 30147 27860 30159 27863
rect 30650 27860 30656 27872
rect 30147 27832 30656 27860
rect 30147 27829 30159 27832
rect 30101 27823 30159 27829
rect 30650 27820 30656 27832
rect 30708 27820 30714 27872
rect 30926 27820 30932 27872
rect 30984 27820 30990 27872
rect 31018 27820 31024 27872
rect 31076 27820 31082 27872
rect 31754 27820 31760 27872
rect 31812 27860 31818 27872
rect 32582 27860 32588 27872
rect 31812 27832 32588 27860
rect 31812 27820 31818 27832
rect 32582 27820 32588 27832
rect 32640 27820 32646 27872
rect 34698 27820 34704 27872
rect 34756 27820 34762 27872
rect 1104 27770 35248 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 35248 27770
rect 1104 27696 35248 27718
rect 2866 27616 2872 27668
rect 2924 27656 2930 27668
rect 4046 27659 4104 27665
rect 4046 27656 4058 27659
rect 2924 27628 4058 27656
rect 2924 27616 2930 27628
rect 4046 27625 4058 27628
rect 4092 27625 4104 27659
rect 4046 27619 4104 27625
rect 19426 27616 19432 27668
rect 19484 27656 19490 27668
rect 19889 27659 19947 27665
rect 19484 27628 19748 27656
rect 19484 27616 19490 27628
rect 19518 27548 19524 27600
rect 19576 27548 19582 27600
rect 19720 27597 19748 27628
rect 19889 27625 19901 27659
rect 19935 27656 19947 27659
rect 20070 27656 20076 27668
rect 19935 27628 20076 27656
rect 19935 27625 19947 27628
rect 19889 27619 19947 27625
rect 19705 27591 19763 27597
rect 19705 27557 19717 27591
rect 19751 27557 19763 27591
rect 19705 27551 19763 27557
rect 14918 27480 14924 27532
rect 14976 27520 14982 27532
rect 15289 27523 15347 27529
rect 14976 27492 15240 27520
rect 14976 27480 14982 27492
rect 3789 27455 3847 27461
rect 3789 27452 3801 27455
rect 3620 27424 3801 27452
rect 3620 27328 3648 27424
rect 3789 27421 3801 27424
rect 3835 27421 3847 27455
rect 3789 27415 3847 27421
rect 14826 27412 14832 27464
rect 14884 27412 14890 27464
rect 15102 27412 15108 27464
rect 15160 27412 15166 27464
rect 15212 27452 15240 27492
rect 15289 27489 15301 27523
rect 15335 27520 15347 27523
rect 15657 27523 15715 27529
rect 15657 27520 15669 27523
rect 15335 27492 15669 27520
rect 15335 27489 15347 27492
rect 15289 27483 15347 27489
rect 15657 27489 15669 27492
rect 15703 27489 15715 27523
rect 15657 27483 15715 27489
rect 16758 27480 16764 27532
rect 16816 27520 16822 27532
rect 19536 27520 19564 27548
rect 19904 27520 19932 27619
rect 20070 27616 20076 27628
rect 20128 27616 20134 27668
rect 21450 27616 21456 27668
rect 21508 27616 21514 27668
rect 22830 27616 22836 27668
rect 22888 27656 22894 27668
rect 25206 27659 25264 27665
rect 25206 27656 25218 27659
rect 22888 27628 25218 27656
rect 22888 27616 22894 27628
rect 25206 27625 25218 27628
rect 25252 27625 25264 27659
rect 25206 27619 25264 27625
rect 33686 27616 33692 27668
rect 33744 27616 33750 27668
rect 34146 27616 34152 27668
rect 34204 27616 34210 27668
rect 21468 27588 21496 27616
rect 23569 27591 23627 27597
rect 23569 27588 23581 27591
rect 21468 27560 23581 27588
rect 23569 27557 23581 27560
rect 23615 27557 23627 27591
rect 23569 27551 23627 27557
rect 26697 27591 26755 27597
rect 26697 27557 26709 27591
rect 26743 27588 26755 27591
rect 30101 27591 30159 27597
rect 26743 27560 30052 27588
rect 26743 27557 26755 27560
rect 26697 27551 26755 27557
rect 16816 27492 17724 27520
rect 19536 27492 19932 27520
rect 19996 27492 23612 27520
rect 16816 27480 16822 27492
rect 15381 27455 15439 27461
rect 15381 27452 15393 27455
rect 15212 27424 15393 27452
rect 15381 27421 15393 27424
rect 15427 27421 15439 27455
rect 15381 27415 15439 27421
rect 15473 27455 15531 27461
rect 15473 27421 15485 27455
rect 15519 27452 15531 27455
rect 15519 27424 15976 27452
rect 15519 27421 15531 27424
rect 15473 27415 15531 27421
rect 4154 27344 4160 27396
rect 4212 27384 4218 27396
rect 14921 27387 14979 27393
rect 4212 27356 4554 27384
rect 4212 27344 4218 27356
rect 14921 27353 14933 27387
rect 14967 27384 14979 27387
rect 15488 27384 15516 27415
rect 14967 27356 15516 27384
rect 14967 27353 14979 27356
rect 14921 27347 14979 27353
rect 15948 27328 15976 27424
rect 17310 27412 17316 27464
rect 17368 27452 17374 27464
rect 17405 27455 17463 27461
rect 17405 27452 17417 27455
rect 17368 27424 17417 27452
rect 17368 27412 17374 27424
rect 17405 27421 17417 27424
rect 17451 27421 17463 27455
rect 17405 27415 17463 27421
rect 17589 27455 17647 27461
rect 17589 27421 17601 27455
rect 17635 27421 17647 27455
rect 17696 27452 17724 27492
rect 19996 27452 20024 27492
rect 17696 27424 20024 27452
rect 17589 27415 17647 27421
rect 17604 27384 17632 27415
rect 20162 27412 20168 27464
rect 20220 27412 20226 27464
rect 23382 27452 23388 27464
rect 22066 27424 23388 27452
rect 16868 27356 17632 27384
rect 18233 27387 18291 27393
rect 16868 27328 16896 27356
rect 18233 27353 18245 27387
rect 18279 27384 18291 27387
rect 18279 27356 18736 27384
rect 18279 27353 18291 27356
rect 18233 27347 18291 27353
rect 18708 27328 18736 27356
rect 3602 27276 3608 27328
rect 3660 27276 3666 27328
rect 5534 27276 5540 27328
rect 5592 27276 5598 27328
rect 5810 27276 5816 27328
rect 5868 27276 5874 27328
rect 15654 27276 15660 27328
rect 15712 27276 15718 27328
rect 15930 27276 15936 27328
rect 15988 27276 15994 27328
rect 16850 27276 16856 27328
rect 16908 27276 16914 27328
rect 17494 27276 17500 27328
rect 17552 27276 17558 27328
rect 17954 27276 17960 27328
rect 18012 27316 18018 27328
rect 18506 27316 18512 27328
rect 18012 27288 18512 27316
rect 18012 27276 18018 27288
rect 18506 27276 18512 27288
rect 18564 27276 18570 27328
rect 18690 27276 18696 27328
rect 18748 27276 18754 27328
rect 21450 27276 21456 27328
rect 21508 27316 21514 27328
rect 22066 27316 22094 27424
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 23474 27412 23480 27464
rect 23532 27412 23538 27464
rect 23584 27452 23612 27492
rect 23658 27480 23664 27532
rect 23716 27480 23722 27532
rect 29825 27523 29883 27529
rect 29825 27489 29837 27523
rect 29871 27489 29883 27523
rect 30024 27520 30052 27560
rect 30101 27557 30113 27591
rect 30147 27588 30159 27591
rect 30147 27560 30972 27588
rect 30147 27557 30159 27560
rect 30101 27551 30159 27557
rect 30469 27523 30527 27529
rect 30469 27520 30481 27523
rect 30024 27492 30481 27520
rect 29825 27483 29883 27489
rect 30469 27489 30481 27492
rect 30515 27489 30527 27523
rect 30469 27483 30527 27489
rect 30561 27523 30619 27529
rect 30561 27489 30573 27523
rect 30607 27520 30619 27523
rect 30607 27492 30788 27520
rect 30607 27489 30619 27492
rect 30561 27483 30619 27489
rect 24857 27455 24915 27461
rect 24857 27452 24869 27455
rect 23584 27424 24869 27452
rect 24857 27421 24869 27424
rect 24903 27452 24915 27455
rect 24949 27455 25007 27461
rect 24949 27452 24961 27455
rect 24903 27424 24961 27452
rect 24903 27421 24915 27424
rect 24857 27415 24915 27421
rect 24949 27421 24961 27424
rect 24995 27421 25007 27455
rect 27157 27455 27215 27461
rect 27157 27452 27169 27455
rect 24949 27415 25007 27421
rect 27080 27424 27169 27452
rect 21508 27288 22094 27316
rect 24964 27316 24992 27415
rect 25958 27344 25964 27396
rect 26016 27344 26022 27396
rect 27080 27328 27108 27424
rect 27157 27421 27169 27424
rect 27203 27421 27215 27455
rect 27157 27415 27215 27421
rect 29730 27412 29736 27464
rect 29788 27412 29794 27464
rect 29840 27452 29868 27483
rect 30193 27455 30251 27461
rect 30193 27452 30205 27455
rect 29840 27424 30205 27452
rect 30193 27421 30205 27424
rect 30239 27421 30251 27455
rect 30193 27415 30251 27421
rect 30377 27455 30435 27461
rect 30377 27421 30389 27455
rect 30423 27421 30435 27455
rect 30377 27415 30435 27421
rect 30392 27384 30420 27415
rect 30024 27356 30420 27384
rect 30484 27384 30512 27483
rect 30650 27412 30656 27464
rect 30708 27412 30714 27464
rect 30760 27452 30788 27492
rect 30834 27480 30840 27532
rect 30892 27480 30898 27532
rect 30944 27520 30972 27560
rect 33134 27548 33140 27600
rect 33192 27548 33198 27600
rect 31665 27523 31723 27529
rect 31665 27520 31677 27523
rect 30944 27492 31677 27520
rect 31665 27489 31677 27492
rect 31711 27489 31723 27523
rect 34698 27520 34704 27532
rect 31665 27483 31723 27489
rect 34256 27492 34704 27520
rect 31018 27452 31024 27464
rect 30760 27424 31024 27452
rect 31018 27412 31024 27424
rect 31076 27412 31082 27464
rect 31113 27455 31171 27461
rect 31113 27421 31125 27455
rect 31159 27452 31171 27455
rect 31389 27455 31447 27461
rect 31159 27424 31248 27452
rect 31159 27421 31171 27424
rect 31113 27415 31171 27421
rect 31220 27396 31248 27424
rect 31389 27421 31401 27455
rect 31435 27421 31447 27455
rect 31389 27415 31447 27421
rect 31202 27384 31208 27396
rect 30484 27356 31208 27384
rect 30024 27328 30052 27356
rect 31202 27344 31208 27356
rect 31260 27344 31266 27396
rect 26694 27316 26700 27328
rect 24964 27288 26700 27316
rect 21508 27276 21514 27288
rect 26694 27276 26700 27288
rect 26752 27276 26758 27328
rect 27062 27276 27068 27328
rect 27120 27276 27126 27328
rect 27246 27276 27252 27328
rect 27304 27276 27310 27328
rect 30006 27276 30012 27328
rect 30064 27276 30070 27328
rect 30834 27276 30840 27328
rect 30892 27276 30898 27328
rect 31404 27316 31432 27415
rect 33410 27412 33416 27464
rect 33468 27452 33474 27464
rect 33597 27455 33655 27461
rect 33597 27452 33609 27455
rect 33468 27424 33609 27452
rect 33468 27412 33474 27424
rect 33597 27421 33609 27424
rect 33643 27452 33655 27455
rect 34146 27452 34152 27464
rect 33643 27424 34152 27452
rect 33643 27421 33655 27424
rect 33597 27415 33655 27421
rect 34146 27412 34152 27424
rect 34204 27452 34210 27464
rect 34256 27461 34284 27492
rect 34698 27480 34704 27492
rect 34756 27480 34762 27532
rect 34241 27455 34299 27461
rect 34241 27452 34253 27455
rect 34204 27424 34253 27452
rect 34204 27412 34210 27424
rect 34241 27421 34253 27424
rect 34287 27421 34299 27455
rect 34241 27415 34299 27421
rect 31754 27384 31760 27396
rect 31726 27344 31760 27384
rect 31812 27344 31818 27396
rect 33321 27387 33379 27393
rect 33321 27384 33333 27387
rect 32890 27356 33333 27384
rect 33321 27353 33333 27356
rect 33367 27353 33379 27387
rect 33321 27347 33379 27353
rect 31726 27316 31754 27344
rect 31404 27288 31754 27316
rect 1104 27226 35236 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 35236 27226
rect 1104 27152 35236 27174
rect 4154 27072 4160 27124
rect 4212 27072 4218 27124
rect 15654 27072 15660 27124
rect 15712 27112 15718 27124
rect 17681 27115 17739 27121
rect 15712 27084 17080 27112
rect 15712 27072 15718 27084
rect 15930 27004 15936 27056
rect 15988 27004 15994 27056
rect 16945 27047 17003 27053
rect 16945 27044 16957 27047
rect 16868 27016 16957 27044
rect 4065 26979 4123 26985
rect 4065 26945 4077 26979
rect 4111 26976 4123 26979
rect 14829 26979 14887 26985
rect 4111 26948 4660 26976
rect 4111 26945 4123 26948
rect 4065 26939 4123 26945
rect 3602 26732 3608 26784
rect 3660 26732 3666 26784
rect 4632 26781 4660 26948
rect 14829 26945 14841 26979
rect 14875 26976 14887 26979
rect 14918 26976 14924 26988
rect 14875 26948 14924 26976
rect 14875 26945 14887 26948
rect 14829 26939 14887 26945
rect 14918 26936 14924 26948
rect 14976 26936 14982 26988
rect 15473 26979 15531 26985
rect 15473 26945 15485 26979
rect 15519 26976 15531 26979
rect 16117 26979 16175 26985
rect 16117 26976 16129 26979
rect 15519 26948 16129 26976
rect 15519 26945 15531 26948
rect 15473 26939 15531 26945
rect 16117 26945 16129 26948
rect 16163 26945 16175 26979
rect 16117 26939 16175 26945
rect 14737 26911 14795 26917
rect 14737 26877 14749 26911
rect 14783 26877 14795 26911
rect 15381 26911 15439 26917
rect 15381 26908 15393 26911
rect 14737 26871 14795 26877
rect 15212 26880 15393 26908
rect 4617 26775 4675 26781
rect 4617 26741 4629 26775
rect 4663 26772 4675 26775
rect 4982 26772 4988 26784
rect 4663 26744 4988 26772
rect 4663 26741 4675 26744
rect 4617 26735 4675 26741
rect 4982 26732 4988 26744
rect 5040 26732 5046 26784
rect 14752 26772 14780 26871
rect 15212 26849 15240 26880
rect 15381 26877 15393 26880
rect 15427 26877 15439 26911
rect 15381 26871 15439 26877
rect 15197 26843 15255 26849
rect 15197 26809 15209 26843
rect 15243 26809 15255 26843
rect 15488 26840 15516 26939
rect 16298 26936 16304 26988
rect 16356 26976 16362 26988
rect 16761 26979 16819 26985
rect 16761 26976 16773 26979
rect 16356 26948 16773 26976
rect 16356 26936 16362 26948
rect 16761 26945 16773 26948
rect 16807 26945 16819 26979
rect 16761 26939 16819 26945
rect 16868 26908 16896 27016
rect 16945 27013 16957 27016
rect 16991 27013 17003 27047
rect 16945 27007 17003 27013
rect 17052 26976 17080 27084
rect 17681 27081 17693 27115
rect 17727 27112 17739 27115
rect 20070 27112 20076 27124
rect 17727 27084 20076 27112
rect 17727 27081 17739 27084
rect 17681 27075 17739 27081
rect 20070 27072 20076 27084
rect 20128 27112 20134 27124
rect 20128 27084 20300 27112
rect 20128 27072 20134 27084
rect 17129 27047 17187 27053
rect 17129 27013 17141 27047
rect 17175 27044 17187 27047
rect 19334 27044 19340 27056
rect 17175 27016 17908 27044
rect 17175 27013 17187 27016
rect 17129 27007 17187 27013
rect 17221 26979 17279 26985
rect 17221 26976 17233 26979
rect 17052 26948 17233 26976
rect 17221 26945 17233 26948
rect 17267 26945 17279 26979
rect 17221 26939 17279 26945
rect 17310 26936 17316 26988
rect 17368 26976 17374 26988
rect 17405 26979 17463 26985
rect 17405 26976 17417 26979
rect 17368 26948 17417 26976
rect 17368 26936 17374 26948
rect 17405 26945 17417 26948
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 17494 26936 17500 26988
rect 17552 26976 17558 26988
rect 17880 26985 17908 27016
rect 18340 27016 19340 27044
rect 18340 26985 18368 27016
rect 19334 27004 19340 27016
rect 19392 27004 19398 27056
rect 20272 27044 20300 27084
rect 22554 27072 22560 27124
rect 22612 27072 22618 27124
rect 23293 27115 23351 27121
rect 23293 27081 23305 27115
rect 23339 27112 23351 27115
rect 23474 27112 23480 27124
rect 23339 27084 23480 27112
rect 23339 27081 23351 27084
rect 23293 27075 23351 27081
rect 23474 27072 23480 27084
rect 23532 27072 23538 27124
rect 23658 27072 23664 27124
rect 23716 27112 23722 27124
rect 24489 27115 24547 27121
rect 24489 27112 24501 27115
rect 23716 27084 24501 27112
rect 23716 27072 23722 27084
rect 24489 27081 24501 27084
rect 24535 27081 24547 27115
rect 24489 27075 24547 27081
rect 25958 27072 25964 27124
rect 26016 27072 26022 27124
rect 26694 27072 26700 27124
rect 26752 27072 26758 27124
rect 27062 27072 27068 27124
rect 27120 27072 27126 27124
rect 27246 27072 27252 27124
rect 27304 27072 27310 27124
rect 28721 27115 28779 27121
rect 28721 27081 28733 27115
rect 28767 27112 28779 27115
rect 29730 27112 29736 27124
rect 28767 27084 29736 27112
rect 28767 27081 28779 27084
rect 28721 27075 28779 27081
rect 29730 27072 29736 27084
rect 29788 27072 29794 27124
rect 30834 27072 30840 27124
rect 30892 27072 30898 27124
rect 31481 27115 31539 27121
rect 31481 27081 31493 27115
rect 31527 27112 31539 27115
rect 32950 27112 32956 27124
rect 31527 27084 32956 27112
rect 31527 27081 31539 27084
rect 31481 27075 31539 27081
rect 32950 27072 32956 27084
rect 33008 27072 33014 27124
rect 33137 27115 33195 27121
rect 33137 27081 33149 27115
rect 33183 27112 33195 27115
rect 33410 27112 33416 27124
rect 33183 27084 33416 27112
rect 33183 27081 33195 27084
rect 33137 27075 33195 27081
rect 21634 27044 21640 27056
rect 20272 27016 20392 27044
rect 17773 26979 17831 26985
rect 17773 26976 17785 26979
rect 17552 26948 17785 26976
rect 17552 26936 17558 26948
rect 17773 26945 17785 26948
rect 17819 26945 17831 26979
rect 17773 26939 17831 26945
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26945 17923 26979
rect 17865 26939 17923 26945
rect 18049 26979 18107 26985
rect 18049 26945 18061 26979
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 18325 26979 18383 26985
rect 18325 26945 18337 26979
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18064 26908 18092 26939
rect 18414 26936 18420 26988
rect 18472 26936 18478 26988
rect 18506 26936 18512 26988
rect 18564 26976 18570 26988
rect 18601 26979 18659 26985
rect 18601 26976 18613 26979
rect 18564 26948 18613 26976
rect 18564 26936 18570 26948
rect 18601 26945 18613 26948
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18690 26936 18696 26988
rect 18748 26936 18754 26988
rect 18782 26936 18788 26988
rect 18840 26936 18846 26988
rect 19518 26936 19524 26988
rect 19576 26936 19582 26988
rect 19613 26979 19671 26985
rect 19613 26945 19625 26979
rect 19659 26945 19671 26979
rect 19613 26939 19671 26945
rect 15856 26880 16896 26908
rect 17604 26880 18092 26908
rect 18233 26911 18291 26917
rect 15856 26852 15884 26880
rect 15197 26803 15255 26809
rect 15396 26812 15516 26840
rect 15396 26784 15424 26812
rect 15838 26800 15844 26852
rect 15896 26800 15902 26852
rect 16850 26800 16856 26852
rect 16908 26840 16914 26852
rect 17604 26840 17632 26880
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 19334 26908 19340 26920
rect 18279 26880 19340 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 19334 26868 19340 26880
rect 19392 26868 19398 26920
rect 19628 26908 19656 26939
rect 20070 26936 20076 26988
rect 20128 26936 20134 26988
rect 20254 26936 20260 26988
rect 20312 26936 20318 26988
rect 20364 26985 20392 27016
rect 20640 27016 21640 27044
rect 20640 26985 20668 27016
rect 21634 27004 21640 27016
rect 21692 27044 21698 27056
rect 21692 27016 22416 27044
rect 21692 27004 21698 27016
rect 20349 26979 20407 26985
rect 20349 26945 20361 26979
rect 20395 26945 20407 26979
rect 20349 26939 20407 26945
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26945 20683 26979
rect 20625 26939 20683 26945
rect 20714 26936 20720 26988
rect 20772 26976 20778 26988
rect 20772 26948 20944 26976
rect 20772 26936 20778 26948
rect 20165 26911 20223 26917
rect 20165 26908 20177 26911
rect 19628 26880 20177 26908
rect 20165 26877 20177 26880
rect 20211 26877 20223 26911
rect 20165 26871 20223 26877
rect 20533 26911 20591 26917
rect 20533 26877 20545 26911
rect 20579 26908 20591 26911
rect 20806 26908 20812 26920
rect 20579 26880 20812 26908
rect 20579 26877 20591 26880
rect 20533 26871 20591 26877
rect 20806 26868 20812 26880
rect 20864 26868 20870 26920
rect 20916 26908 20944 26948
rect 21818 26936 21824 26988
rect 21876 26936 21882 26988
rect 22005 26979 22063 26985
rect 22005 26945 22017 26979
rect 22051 26976 22063 26979
rect 22278 26976 22284 26988
rect 22051 26948 22284 26976
rect 22051 26945 22063 26948
rect 22005 26939 22063 26945
rect 22278 26936 22284 26948
rect 22336 26936 22342 26988
rect 22388 26985 22416 27016
rect 23382 27004 23388 27056
rect 23440 27044 23446 27056
rect 27080 27044 27108 27072
rect 23440 27016 24072 27044
rect 23440 27004 23446 27016
rect 24044 26985 24072 27016
rect 25884 27016 27108 27044
rect 27264 27044 27292 27072
rect 27264 27016 27738 27044
rect 22373 26979 22431 26985
rect 22373 26945 22385 26979
rect 22419 26976 22431 26979
rect 24029 26979 24087 26985
rect 22419 26966 23428 26976
rect 22419 26948 23612 26966
rect 22419 26945 22431 26948
rect 22373 26939 22431 26945
rect 23400 26938 23612 26948
rect 24029 26945 24041 26979
rect 24075 26945 24087 26979
rect 24703 26979 24761 26985
rect 24703 26976 24715 26979
rect 24029 26939 24087 26945
rect 24136 26948 24715 26976
rect 22097 26911 22155 26917
rect 22097 26908 22109 26911
rect 20916 26880 22109 26908
rect 22097 26877 22109 26880
rect 22143 26877 22155 26911
rect 22097 26871 22155 26877
rect 22189 26911 22247 26917
rect 22189 26877 22201 26911
rect 22235 26877 22247 26911
rect 23584 26908 23612 26938
rect 23753 26911 23811 26917
rect 23753 26908 23765 26911
rect 23584 26880 23765 26908
rect 22189 26871 22247 26877
rect 23753 26877 23765 26880
rect 23799 26908 23811 26911
rect 23937 26911 23995 26917
rect 23937 26908 23949 26911
rect 23799 26880 23949 26908
rect 23799 26877 23811 26880
rect 23753 26871 23811 26877
rect 23937 26877 23949 26880
rect 23983 26908 23995 26911
rect 24136 26908 24164 26948
rect 24703 26945 24715 26948
rect 24749 26945 24761 26979
rect 24703 26939 24761 26945
rect 24854 26936 24860 26988
rect 24912 26936 24918 26988
rect 25884 26985 25912 27016
rect 25777 26979 25835 26985
rect 25777 26945 25789 26979
rect 25823 26976 25835 26979
rect 25869 26979 25927 26985
rect 25869 26976 25881 26979
rect 25823 26948 25881 26976
rect 25823 26945 25835 26948
rect 25777 26939 25835 26945
rect 25869 26945 25881 26948
rect 25915 26945 25927 26979
rect 25869 26939 25927 26945
rect 26694 26936 26700 26988
rect 26752 26976 26758 26988
rect 26878 26976 26884 26988
rect 26752 26948 26884 26976
rect 26752 26936 26758 26948
rect 26878 26936 26884 26948
rect 26936 26976 26942 26988
rect 26973 26979 27031 26985
rect 26973 26976 26985 26979
rect 26936 26948 26985 26976
rect 26936 26936 26942 26948
rect 26973 26945 26985 26948
rect 27019 26945 27031 26979
rect 26973 26939 27031 26945
rect 28997 26979 29055 26985
rect 28997 26945 29009 26979
rect 29043 26976 29055 26979
rect 30101 26979 30159 26985
rect 30101 26976 30113 26979
rect 29043 26948 29408 26976
rect 29043 26945 29055 26948
rect 28997 26939 29055 26945
rect 27249 26911 27307 26917
rect 27249 26908 27261 26911
rect 23983 26880 24164 26908
rect 27080 26880 27261 26908
rect 23983 26877 23995 26880
rect 23937 26871 23995 26877
rect 16908 26812 17632 26840
rect 18969 26843 19027 26849
rect 16908 26800 16914 26812
rect 18969 26809 18981 26843
rect 19015 26840 19027 26843
rect 22204 26840 22232 26871
rect 22370 26840 22376 26852
rect 19015 26812 22094 26840
rect 22204 26812 22376 26840
rect 19015 26809 19027 26812
rect 18969 26803 19027 26809
rect 15286 26772 15292 26784
rect 14752 26744 15292 26772
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 15378 26732 15384 26784
rect 15436 26732 15442 26784
rect 19334 26732 19340 26784
rect 19392 26732 19398 26784
rect 22066 26772 22094 26812
rect 22370 26800 22376 26812
rect 22428 26800 22434 26852
rect 23382 26800 23388 26852
rect 23440 26840 23446 26852
rect 23477 26843 23535 26849
rect 23477 26840 23489 26843
rect 23440 26812 23489 26840
rect 23440 26800 23446 26812
rect 23477 26809 23489 26812
rect 23523 26809 23535 26843
rect 27080 26840 27108 26880
rect 27249 26877 27261 26880
rect 27295 26877 27307 26911
rect 27249 26871 27307 26877
rect 23477 26803 23535 26809
rect 23584 26812 27108 26840
rect 23584 26772 23612 26812
rect 22066 26744 23612 26772
rect 24302 26732 24308 26784
rect 24360 26732 24366 26784
rect 28902 26732 28908 26784
rect 28960 26732 28966 26784
rect 29380 26781 29408 26948
rect 30024 26948 30113 26976
rect 30024 26784 30052 26948
rect 30101 26945 30113 26948
rect 30147 26945 30159 26979
rect 30101 26939 30159 26945
rect 30193 26911 30251 26917
rect 30193 26877 30205 26911
rect 30239 26908 30251 26911
rect 30852 26908 30880 27072
rect 32769 27047 32827 27053
rect 32769 27013 32781 27047
rect 32815 27044 32827 27047
rect 33152 27044 33180 27075
rect 33410 27072 33416 27084
rect 33468 27072 33474 27124
rect 32815 27016 33180 27044
rect 32815 27013 32827 27016
rect 32769 27007 32827 27013
rect 31113 26979 31171 26985
rect 31113 26945 31125 26979
rect 31159 26976 31171 26979
rect 31202 26976 31208 26988
rect 31159 26948 31208 26976
rect 31159 26945 31171 26948
rect 31113 26939 31171 26945
rect 31202 26936 31208 26948
rect 31260 26936 31266 26988
rect 33686 26936 33692 26988
rect 33744 26936 33750 26988
rect 34698 26936 34704 26988
rect 34756 26936 34762 26988
rect 30239 26880 30880 26908
rect 30239 26877 30251 26880
rect 30193 26871 30251 26877
rect 30926 26868 30932 26920
rect 30984 26908 30990 26920
rect 31021 26911 31079 26917
rect 31021 26908 31033 26911
rect 30984 26880 31033 26908
rect 30984 26868 30990 26880
rect 31021 26877 31033 26880
rect 31067 26877 31079 26911
rect 31021 26871 31079 26877
rect 30469 26843 30527 26849
rect 30469 26809 30481 26843
rect 30515 26840 30527 26843
rect 30515 26812 31754 26840
rect 30515 26809 30527 26812
rect 30469 26803 30527 26809
rect 29365 26775 29423 26781
rect 29365 26741 29377 26775
rect 29411 26772 29423 26775
rect 29914 26772 29920 26784
rect 29411 26744 29920 26772
rect 29411 26741 29423 26744
rect 29365 26735 29423 26741
rect 29914 26732 29920 26744
rect 29972 26732 29978 26784
rect 30006 26732 30012 26784
rect 30064 26732 30070 26784
rect 31726 26772 31754 26812
rect 33042 26772 33048 26784
rect 31726 26744 33048 26772
rect 33042 26732 33048 26744
rect 33100 26732 33106 26784
rect 1104 26682 35248 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 35248 26682
rect 1104 26608 35248 26630
rect 5810 26528 5816 26580
rect 5868 26528 5874 26580
rect 14826 26528 14832 26580
rect 14884 26568 14890 26580
rect 15013 26571 15071 26577
rect 15013 26568 15025 26571
rect 14884 26540 15025 26568
rect 14884 26528 14890 26540
rect 15013 26537 15025 26540
rect 15059 26537 15071 26571
rect 15013 26531 15071 26537
rect 16758 26528 16764 26580
rect 16816 26528 16822 26580
rect 16850 26528 16856 26580
rect 16908 26528 16914 26580
rect 17494 26528 17500 26580
rect 17552 26568 17558 26580
rect 17552 26540 17816 26568
rect 17552 26528 17558 26540
rect 1670 26392 1676 26444
rect 1728 26392 1734 26444
rect 3602 26432 3608 26444
rect 3344 26404 3608 26432
rect 1397 26367 1455 26373
rect 1397 26333 1409 26367
rect 1443 26333 1455 26367
rect 1397 26327 1455 26333
rect 1412 26228 1440 26327
rect 2130 26256 2136 26308
rect 2188 26256 2194 26308
rect 2038 26228 2044 26240
rect 1412 26200 2044 26228
rect 2038 26188 2044 26200
rect 2096 26228 2102 26240
rect 3344 26228 3372 26404
rect 3602 26392 3608 26404
rect 3660 26432 3666 26444
rect 3789 26435 3847 26441
rect 3789 26432 3801 26435
rect 3660 26404 3801 26432
rect 3660 26392 3666 26404
rect 3789 26401 3801 26404
rect 3835 26432 3847 26435
rect 5828 26432 5856 26528
rect 7009 26503 7067 26509
rect 7009 26469 7021 26503
rect 7055 26469 7067 26503
rect 7009 26463 7067 26469
rect 11333 26503 11391 26509
rect 11333 26469 11345 26503
rect 11379 26500 11391 26503
rect 16776 26500 16804 26528
rect 11379 26472 16804 26500
rect 11379 26469 11391 26472
rect 11333 26463 11391 26469
rect 3835 26404 5856 26432
rect 7024 26432 7052 26463
rect 9217 26435 9275 26441
rect 9217 26432 9229 26435
rect 7024 26404 9229 26432
rect 3835 26401 3847 26404
rect 3789 26395 3847 26401
rect 9217 26401 9229 26404
rect 9263 26401 9275 26435
rect 9217 26395 9275 26401
rect 9306 26392 9312 26444
rect 9364 26432 9370 26444
rect 9766 26432 9772 26444
rect 9364 26404 9772 26432
rect 9364 26392 9370 26404
rect 9766 26392 9772 26404
rect 9824 26432 9830 26444
rect 11348 26432 11376 26463
rect 9824 26404 11376 26432
rect 9824 26392 9830 26404
rect 12986 26392 12992 26444
rect 13044 26432 13050 26444
rect 13449 26435 13507 26441
rect 13449 26432 13461 26435
rect 13044 26404 13461 26432
rect 13044 26392 13050 26404
rect 13449 26401 13461 26404
rect 13495 26401 13507 26435
rect 13449 26395 13507 26401
rect 15838 26392 15844 26444
rect 15896 26432 15902 26444
rect 15896 26404 16908 26432
rect 15896 26392 15902 26404
rect 6822 26324 6828 26376
rect 6880 26324 6886 26376
rect 8941 26367 8999 26373
rect 8941 26333 8953 26367
rect 8987 26333 8999 26367
rect 8941 26327 8999 26333
rect 3421 26299 3479 26305
rect 3421 26265 3433 26299
rect 3467 26296 3479 26299
rect 3970 26296 3976 26308
rect 3467 26268 3976 26296
rect 3467 26265 3479 26268
rect 3421 26259 3479 26265
rect 3970 26256 3976 26268
rect 4028 26256 4034 26308
rect 4062 26256 4068 26308
rect 4120 26256 4126 26308
rect 4706 26256 4712 26308
rect 4764 26256 4770 26308
rect 8294 26256 8300 26308
rect 8352 26296 8358 26308
rect 8956 26296 8984 26327
rect 12894 26324 12900 26376
rect 12952 26364 12958 26376
rect 13357 26367 13415 26373
rect 13357 26364 13369 26367
rect 12952 26336 13369 26364
rect 12952 26324 12958 26336
rect 13357 26333 13369 26336
rect 13403 26333 13415 26367
rect 13357 26327 13415 26333
rect 13630 26324 13636 26376
rect 13688 26324 13694 26376
rect 14918 26324 14924 26376
rect 14976 26364 14982 26376
rect 15197 26367 15255 26373
rect 15197 26364 15209 26367
rect 14976 26336 15209 26364
rect 14976 26324 14982 26336
rect 15197 26333 15209 26336
rect 15243 26333 15255 26367
rect 15197 26327 15255 26333
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26333 15531 26367
rect 16298 26364 16304 26376
rect 15473 26327 15531 26333
rect 15948 26336 16304 26364
rect 9306 26296 9312 26308
rect 8352 26268 9312 26296
rect 8352 26256 8358 26268
rect 9306 26256 9312 26268
rect 9364 26256 9370 26308
rect 9674 26256 9680 26308
rect 9732 26256 9738 26308
rect 10686 26256 10692 26308
rect 10744 26296 10750 26308
rect 10965 26299 11023 26305
rect 10965 26296 10977 26299
rect 10744 26268 10977 26296
rect 10744 26256 10750 26268
rect 10965 26265 10977 26268
rect 11011 26265 11023 26299
rect 10965 26259 11023 26265
rect 13817 26299 13875 26305
rect 13817 26265 13829 26299
rect 13863 26296 13875 26299
rect 15378 26296 15384 26308
rect 13863 26268 15384 26296
rect 13863 26265 13875 26268
rect 13817 26259 13875 26265
rect 15378 26256 15384 26268
rect 15436 26256 15442 26308
rect 15488 26296 15516 26327
rect 15948 26308 15976 26336
rect 16298 26324 16304 26336
rect 16356 26364 16362 26376
rect 16761 26367 16819 26373
rect 16761 26364 16773 26367
rect 16356 26336 16773 26364
rect 16356 26324 16362 26336
rect 16761 26333 16773 26336
rect 16807 26333 16819 26367
rect 16880 26364 16908 26404
rect 16945 26367 17003 26373
rect 16945 26364 16957 26367
rect 16880 26336 16957 26364
rect 16761 26327 16819 26333
rect 16945 26333 16957 26336
rect 16991 26333 17003 26367
rect 17622 26367 17680 26373
rect 17622 26364 17634 26367
rect 16945 26327 17003 26333
rect 17052 26336 17634 26364
rect 15930 26296 15936 26308
rect 15488 26268 15936 26296
rect 15930 26256 15936 26268
rect 15988 26256 15994 26308
rect 17052 26296 17080 26336
rect 17622 26333 17634 26336
rect 17668 26333 17680 26367
rect 17622 26327 17680 26333
rect 17788 26305 17816 26540
rect 18414 26528 18420 26580
rect 18472 26568 18478 26580
rect 18601 26571 18659 26577
rect 18601 26568 18613 26571
rect 18472 26540 18613 26568
rect 18472 26528 18478 26540
rect 18601 26537 18613 26540
rect 18647 26537 18659 26571
rect 18601 26531 18659 26537
rect 19334 26528 19340 26580
rect 19392 26528 19398 26580
rect 20070 26528 20076 26580
rect 20128 26568 20134 26580
rect 20165 26571 20223 26577
rect 20165 26568 20177 26571
rect 20128 26540 20177 26568
rect 20128 26528 20134 26540
rect 20165 26537 20177 26540
rect 20211 26537 20223 26571
rect 20165 26531 20223 26537
rect 20346 26528 20352 26580
rect 20404 26528 20410 26580
rect 21450 26528 21456 26580
rect 21508 26528 21514 26580
rect 21637 26571 21695 26577
rect 21637 26537 21649 26571
rect 21683 26568 21695 26571
rect 21818 26568 21824 26580
rect 21683 26540 21824 26568
rect 21683 26537 21695 26540
rect 21637 26531 21695 26537
rect 21818 26528 21824 26540
rect 21876 26528 21882 26580
rect 22005 26571 22063 26577
rect 22005 26537 22017 26571
rect 22051 26568 22063 26571
rect 22094 26568 22100 26580
rect 22051 26540 22100 26568
rect 22051 26537 22063 26540
rect 22005 26531 22063 26537
rect 22094 26528 22100 26540
rect 22152 26528 22158 26580
rect 22278 26528 22284 26580
rect 22336 26528 22342 26580
rect 23382 26528 23388 26580
rect 23440 26568 23446 26580
rect 24854 26568 24860 26580
rect 23440 26540 24860 26568
rect 23440 26528 23446 26540
rect 24854 26528 24860 26540
rect 24912 26528 24918 26580
rect 26878 26528 26884 26580
rect 26936 26528 26942 26580
rect 28813 26571 28871 26577
rect 28813 26537 28825 26571
rect 28859 26568 28871 26571
rect 30006 26568 30012 26580
rect 28859 26540 30012 26568
rect 28859 26537 28871 26540
rect 28813 26531 28871 26537
rect 30006 26528 30012 26540
rect 30064 26528 30070 26580
rect 30837 26571 30895 26577
rect 30837 26537 30849 26571
rect 30883 26568 30895 26571
rect 31018 26568 31024 26580
rect 30883 26540 31024 26568
rect 30883 26537 30895 26540
rect 30837 26531 30895 26537
rect 31018 26528 31024 26540
rect 31076 26528 31082 26580
rect 34517 26571 34575 26577
rect 34517 26537 34529 26571
rect 34563 26568 34575 26571
rect 34790 26568 34796 26580
rect 34563 26540 34796 26568
rect 34563 26537 34575 26540
rect 34517 26531 34575 26537
rect 34790 26528 34796 26540
rect 34848 26528 34854 26580
rect 18141 26435 18199 26441
rect 18141 26401 18153 26435
rect 18187 26432 18199 26435
rect 18432 26432 18460 26528
rect 19352 26500 19380 26528
rect 19352 26472 24256 26500
rect 19518 26432 19524 26444
rect 18187 26404 18460 26432
rect 18524 26404 19524 26432
rect 18187 26401 18199 26404
rect 18141 26395 18199 26401
rect 18046 26324 18052 26376
rect 18104 26324 18110 26376
rect 18230 26324 18236 26376
rect 18288 26324 18294 26376
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26333 18475 26367
rect 18417 26327 18475 26333
rect 16868 26268 17080 26296
rect 17747 26299 17816 26305
rect 2096 26200 3372 26228
rect 2096 26188 2102 26200
rect 5534 26188 5540 26240
rect 5592 26188 5598 26240
rect 13262 26188 13268 26240
rect 13320 26188 13326 26240
rect 16390 26188 16396 26240
rect 16448 26228 16454 26240
rect 16868 26228 16896 26268
rect 17747 26265 17759 26299
rect 17793 26296 17816 26299
rect 18432 26296 18460 26327
rect 17793 26268 18460 26296
rect 17793 26265 17805 26268
rect 17747 26259 17805 26265
rect 16448 26200 16896 26228
rect 17497 26231 17555 26237
rect 16448 26188 16454 26200
rect 17497 26197 17509 26231
rect 17543 26228 17555 26231
rect 18524 26228 18552 26404
rect 19518 26392 19524 26404
rect 19576 26392 19582 26444
rect 19996 26404 21404 26432
rect 19996 26376 20024 26404
rect 18782 26324 18788 26376
rect 18840 26324 18846 26376
rect 19978 26324 19984 26376
rect 20036 26324 20042 26376
rect 20349 26367 20407 26373
rect 20349 26333 20361 26367
rect 20395 26364 20407 26367
rect 20438 26364 20444 26376
rect 20395 26336 20444 26364
rect 20395 26333 20407 26336
rect 20349 26327 20407 26333
rect 18800 26296 18828 26324
rect 20364 26296 20392 26327
rect 20438 26324 20444 26336
rect 20496 26324 20502 26376
rect 21376 26373 21404 26404
rect 21634 26392 21640 26444
rect 21692 26432 21698 26444
rect 22741 26435 22799 26441
rect 22741 26432 22753 26435
rect 21692 26404 22753 26432
rect 21692 26392 21698 26404
rect 20533 26367 20591 26373
rect 20533 26333 20545 26367
rect 20579 26333 20591 26367
rect 20533 26327 20591 26333
rect 21361 26367 21419 26373
rect 21361 26333 21373 26367
rect 21407 26333 21419 26367
rect 21361 26327 21419 26333
rect 20548 26296 20576 26327
rect 18800 26268 20392 26296
rect 20456 26268 20576 26296
rect 21376 26296 21404 26327
rect 21542 26324 21548 26376
rect 21600 26324 21606 26376
rect 22204 26373 22232 26404
rect 22741 26401 22753 26404
rect 22787 26401 22799 26435
rect 22741 26395 22799 26401
rect 21821 26367 21879 26373
rect 21821 26333 21833 26367
rect 21867 26333 21879 26367
rect 21821 26327 21879 26333
rect 22189 26367 22247 26373
rect 22189 26333 22201 26367
rect 22235 26364 22247 26367
rect 22235 26336 22269 26364
rect 22235 26333 22247 26336
rect 22189 26327 22247 26333
rect 21836 26296 21864 26327
rect 22370 26324 22376 26376
rect 22428 26364 22434 26376
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 22428 26336 22477 26364
rect 22428 26324 22434 26336
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 22646 26324 22652 26376
rect 22704 26324 22710 26376
rect 21376 26268 21864 26296
rect 24228 26296 24256 26472
rect 24302 26460 24308 26512
rect 24360 26460 24366 26512
rect 24320 26432 24348 26460
rect 24765 26435 24823 26441
rect 24765 26432 24777 26435
rect 24320 26404 24777 26432
rect 24765 26401 24777 26404
rect 24811 26401 24823 26435
rect 24765 26395 24823 26401
rect 24872 26373 24900 26528
rect 25225 26503 25283 26509
rect 25225 26469 25237 26503
rect 25271 26500 25283 26503
rect 26694 26500 26700 26512
rect 25271 26472 26700 26500
rect 25271 26469 25283 26472
rect 25225 26463 25283 26469
rect 26694 26460 26700 26472
rect 26752 26460 26758 26512
rect 26896 26432 26924 26528
rect 27065 26435 27123 26441
rect 27065 26432 27077 26435
rect 26896 26404 27077 26432
rect 27065 26401 27077 26404
rect 27111 26432 27123 26435
rect 27111 26404 31984 26432
rect 27111 26401 27123 26404
rect 27065 26395 27123 26401
rect 24857 26367 24915 26373
rect 24857 26333 24869 26367
rect 24903 26333 24915 26367
rect 28902 26364 28908 26376
rect 28474 26336 28908 26364
rect 24857 26327 24915 26333
rect 28902 26324 28908 26336
rect 28960 26324 28966 26376
rect 27341 26299 27399 26305
rect 27341 26296 27353 26299
rect 24228 26268 27353 26296
rect 20456 26240 20484 26268
rect 27341 26265 27353 26268
rect 27387 26265 27399 26299
rect 27341 26259 27399 26265
rect 30466 26256 30472 26308
rect 30524 26256 30530 26308
rect 30558 26256 30564 26308
rect 30616 26296 30622 26308
rect 30653 26299 30711 26305
rect 30653 26296 30665 26299
rect 30616 26268 30665 26296
rect 30616 26256 30622 26268
rect 30653 26265 30665 26268
rect 30699 26265 30711 26299
rect 30653 26259 30711 26265
rect 17543 26200 18552 26228
rect 17543 26197 17555 26200
rect 17497 26191 17555 26197
rect 20438 26188 20444 26240
rect 20496 26188 20502 26240
rect 30742 26188 30748 26240
rect 30800 26228 30806 26240
rect 31389 26231 31447 26237
rect 31389 26228 31401 26231
rect 30800 26200 31401 26228
rect 30800 26188 30806 26200
rect 31389 26197 31401 26200
rect 31435 26228 31447 26231
rect 31570 26228 31576 26240
rect 31435 26200 31576 26228
rect 31435 26197 31447 26200
rect 31389 26191 31447 26197
rect 31570 26188 31576 26200
rect 31628 26188 31634 26240
rect 31956 26228 31984 26404
rect 32582 26324 32588 26376
rect 32640 26364 32646 26376
rect 32769 26367 32827 26373
rect 32769 26364 32781 26367
rect 32640 26336 32781 26364
rect 32640 26324 32646 26336
rect 32769 26333 32781 26336
rect 32815 26333 32827 26367
rect 32769 26327 32827 26333
rect 32122 26228 32128 26240
rect 31956 26200 32128 26228
rect 32122 26188 32128 26200
rect 32180 26228 32186 26240
rect 32600 26237 32628 26324
rect 33042 26256 33048 26308
rect 33100 26256 33106 26308
rect 34330 26296 34336 26308
rect 34270 26268 34336 26296
rect 34330 26256 34336 26268
rect 34388 26256 34394 26308
rect 32585 26231 32643 26237
rect 32585 26228 32597 26231
rect 32180 26200 32597 26228
rect 32180 26188 32186 26200
rect 32585 26197 32597 26200
rect 32631 26197 32643 26231
rect 32585 26191 32643 26197
rect 1104 26138 35236 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 35236 26138
rect 1104 26064 35236 26086
rect 1857 26027 1915 26033
rect 1857 25993 1869 26027
rect 1903 26024 1915 26027
rect 2130 26024 2136 26036
rect 1903 25996 2136 26024
rect 1903 25993 1915 25996
rect 1857 25987 1915 25993
rect 2130 25984 2136 25996
rect 2188 25984 2194 26036
rect 4706 25984 4712 26036
rect 4764 25984 4770 26036
rect 6089 26027 6147 26033
rect 6089 25993 6101 26027
rect 6135 26024 6147 26027
rect 6822 26024 6828 26036
rect 6135 25996 6828 26024
rect 6135 25993 6147 25996
rect 6089 25987 6147 25993
rect 6822 25984 6828 25996
rect 6880 25984 6886 26036
rect 9585 26027 9643 26033
rect 9585 25993 9597 26027
rect 9631 26024 9643 26027
rect 9674 26024 9680 26036
rect 9631 25996 9680 26024
rect 9631 25993 9643 25996
rect 9585 25987 9643 25993
rect 9674 25984 9680 25996
rect 9732 25984 9738 26036
rect 13265 26027 13323 26033
rect 13265 25993 13277 26027
rect 13311 26024 13323 26027
rect 13630 26024 13636 26036
rect 13311 25996 13636 26024
rect 13311 25993 13323 25996
rect 13265 25987 13323 25993
rect 13630 25984 13636 25996
rect 13688 25984 13694 26036
rect 17589 26027 17647 26033
rect 17589 26024 17601 26027
rect 15672 25996 17601 26024
rect 15672 25968 15700 25996
rect 17589 25993 17601 25996
rect 17635 25993 17647 26027
rect 17589 25987 17647 25993
rect 17865 26027 17923 26033
rect 17865 25993 17877 26027
rect 17911 26024 17923 26027
rect 18046 26024 18052 26036
rect 17911 25996 18052 26024
rect 17911 25993 17923 25996
rect 17865 25987 17923 25993
rect 1578 25916 1584 25968
rect 1636 25956 1642 25968
rect 2317 25959 2375 25965
rect 2317 25956 2329 25959
rect 1636 25928 2329 25956
rect 1636 25916 1642 25928
rect 2317 25925 2329 25928
rect 2363 25925 2375 25959
rect 3973 25959 4031 25965
rect 3973 25956 3985 25959
rect 3542 25928 3985 25956
rect 2317 25919 2375 25925
rect 3973 25925 3985 25928
rect 4019 25925 4031 25959
rect 12986 25956 12992 25968
rect 3973 25919 4031 25925
rect 12820 25928 12992 25956
rect 934 25848 940 25900
rect 992 25888 998 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 992 25860 1409 25888
rect 992 25848 998 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 1949 25891 2007 25897
rect 1949 25857 1961 25891
rect 1995 25857 2007 25891
rect 4065 25891 4123 25897
rect 4065 25888 4077 25891
rect 1949 25851 2007 25857
rect 3528 25860 4077 25888
rect 1581 25687 1639 25693
rect 1581 25653 1593 25687
rect 1627 25684 1639 25687
rect 1762 25684 1768 25696
rect 1627 25656 1768 25684
rect 1627 25653 1639 25656
rect 1581 25647 1639 25653
rect 1762 25644 1768 25656
rect 1820 25644 1826 25696
rect 1964 25684 1992 25851
rect 2038 25780 2044 25832
rect 2096 25780 2102 25832
rect 2866 25684 2872 25696
rect 1964 25656 2872 25684
rect 2866 25644 2872 25656
rect 2924 25684 2930 25696
rect 3528 25684 3556 25860
rect 4065 25857 4077 25860
rect 4111 25888 4123 25891
rect 4341 25891 4399 25897
rect 4341 25888 4353 25891
rect 4111 25860 4353 25888
rect 4111 25857 4123 25860
rect 4065 25851 4123 25857
rect 4341 25857 4353 25860
rect 4387 25888 4399 25891
rect 4617 25891 4675 25897
rect 4617 25888 4629 25891
rect 4387 25860 4629 25888
rect 4387 25857 4399 25860
rect 4341 25851 4399 25857
rect 4617 25857 4629 25860
rect 4663 25888 4675 25891
rect 5077 25891 5135 25897
rect 5077 25888 5089 25891
rect 4663 25860 5089 25888
rect 4663 25857 4675 25860
rect 4617 25851 4675 25857
rect 5077 25857 5089 25860
rect 5123 25857 5135 25891
rect 5077 25851 5135 25857
rect 5902 25848 5908 25900
rect 5960 25848 5966 25900
rect 12820 25897 12848 25928
rect 12986 25916 12992 25928
rect 13044 25916 13050 25968
rect 15654 25916 15660 25968
rect 15712 25916 15718 25968
rect 16945 25959 17003 25965
rect 16945 25956 16957 25959
rect 16316 25928 16957 25956
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25888 9551 25891
rect 12805 25891 12863 25897
rect 9539 25860 9904 25888
rect 9539 25857 9551 25860
rect 9493 25851 9551 25857
rect 5721 25823 5779 25829
rect 5721 25789 5733 25823
rect 5767 25820 5779 25823
rect 5994 25820 6000 25832
rect 5767 25792 6000 25820
rect 5767 25789 5779 25792
rect 5721 25783 5779 25789
rect 5994 25780 6000 25792
rect 6052 25780 6058 25832
rect 3789 25755 3847 25761
rect 3789 25721 3801 25755
rect 3835 25752 3847 25755
rect 4614 25752 4620 25764
rect 3835 25724 4620 25752
rect 3835 25721 3847 25724
rect 3789 25715 3847 25721
rect 4614 25712 4620 25724
rect 4672 25712 4678 25764
rect 9876 25696 9904 25860
rect 12805 25857 12817 25891
rect 12851 25857 12863 25891
rect 12805 25851 12863 25857
rect 12894 25848 12900 25900
rect 12952 25848 12958 25900
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25888 13139 25891
rect 13633 25891 13691 25897
rect 13633 25888 13645 25891
rect 13127 25860 13645 25888
rect 13127 25857 13139 25860
rect 13081 25851 13139 25857
rect 13633 25857 13645 25860
rect 13679 25857 13691 25891
rect 16114 25888 16120 25900
rect 13633 25851 13691 25857
rect 14016 25860 16120 25888
rect 13262 25780 13268 25832
rect 13320 25820 13326 25832
rect 13541 25823 13599 25829
rect 13541 25820 13553 25823
rect 13320 25792 13553 25820
rect 13320 25780 13326 25792
rect 13541 25789 13553 25792
rect 13587 25789 13599 25823
rect 13541 25783 13599 25789
rect 2924 25656 3556 25684
rect 2924 25644 2930 25656
rect 9858 25644 9864 25696
rect 9916 25684 9922 25696
rect 9953 25687 10011 25693
rect 9953 25684 9965 25687
rect 9916 25656 9965 25684
rect 9916 25644 9922 25656
rect 9953 25653 9965 25656
rect 9999 25653 10011 25687
rect 13648 25684 13676 25851
rect 14016 25761 14044 25860
rect 16114 25848 16120 25860
rect 16172 25848 16178 25900
rect 15930 25780 15936 25832
rect 15988 25820 15994 25832
rect 16316 25820 16344 25928
rect 16945 25925 16957 25928
rect 16991 25925 17003 25959
rect 17604 25956 17632 25987
rect 18046 25984 18052 25996
rect 18104 25984 18110 26036
rect 18690 26024 18696 26036
rect 18156 25996 18696 26024
rect 18156 25956 18184 25996
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 19797 26027 19855 26033
rect 19797 25993 19809 26027
rect 19843 26024 19855 26027
rect 19886 26024 19892 26036
rect 19843 25996 19892 26024
rect 19843 25993 19855 25996
rect 19797 25987 19855 25993
rect 19886 25984 19892 25996
rect 19944 25984 19950 26036
rect 21082 25984 21088 26036
rect 21140 26024 21146 26036
rect 21453 26027 21511 26033
rect 21453 26024 21465 26027
rect 21140 25996 21465 26024
rect 21140 25984 21146 25996
rect 21453 25993 21465 25996
rect 21499 25993 21511 26027
rect 21453 25987 21511 25993
rect 21542 25984 21548 26036
rect 21600 26024 21606 26036
rect 21821 26027 21879 26033
rect 21821 26024 21833 26027
rect 21600 25996 21833 26024
rect 21600 25984 21606 25996
rect 21821 25993 21833 25996
rect 21867 25993 21879 26027
rect 21821 25987 21879 25993
rect 22186 25984 22192 26036
rect 22244 26024 22250 26036
rect 22646 26024 22652 26036
rect 22244 25996 22652 26024
rect 22244 25984 22250 25996
rect 22646 25984 22652 25996
rect 22704 25984 22710 26036
rect 29641 26027 29699 26033
rect 29641 25993 29653 26027
rect 29687 26024 29699 26027
rect 30558 26024 30564 26036
rect 29687 25996 30564 26024
rect 29687 25993 29699 25996
rect 29641 25987 29699 25993
rect 30558 25984 30564 25996
rect 30616 25984 30622 26036
rect 31389 26027 31447 26033
rect 31389 25993 31401 26027
rect 31435 26024 31447 26027
rect 33042 26024 33048 26036
rect 31435 25996 33048 26024
rect 31435 25993 31447 25996
rect 31389 25987 31447 25993
rect 33042 25984 33048 25996
rect 33100 25984 33106 26036
rect 33686 25984 33692 26036
rect 33744 26024 33750 26036
rect 33873 26027 33931 26033
rect 33873 26024 33885 26027
rect 33744 25996 33885 26024
rect 33744 25984 33750 25996
rect 33873 25993 33885 25996
rect 33919 25993 33931 26027
rect 33873 25987 33931 25993
rect 34330 25984 34336 26036
rect 34388 25984 34394 26036
rect 17604 25928 18184 25956
rect 16945 25919 17003 25925
rect 16758 25848 16764 25900
rect 16816 25848 16822 25900
rect 15988 25792 16344 25820
rect 16393 25823 16451 25829
rect 15988 25780 15994 25792
rect 16393 25789 16405 25823
rect 16439 25820 16451 25823
rect 16574 25820 16580 25832
rect 16439 25792 16580 25820
rect 16439 25789 16451 25792
rect 16393 25783 16451 25789
rect 16574 25780 16580 25792
rect 16632 25780 16638 25832
rect 17696 25820 17724 25928
rect 18230 25916 18236 25968
rect 18288 25916 18294 25968
rect 18874 25916 18880 25968
rect 18932 25956 18938 25968
rect 19981 25959 20039 25965
rect 19981 25956 19993 25959
rect 18932 25928 19993 25956
rect 18932 25916 18938 25928
rect 19981 25925 19993 25928
rect 20027 25956 20039 25959
rect 20027 25928 21220 25956
rect 20027 25925 20039 25928
rect 19981 25919 20039 25925
rect 18231 25913 18289 25916
rect 18231 25879 18243 25913
rect 18277 25879 18289 25913
rect 18231 25873 18289 25879
rect 17862 25820 17868 25832
rect 17696 25792 17868 25820
rect 17862 25780 17868 25792
rect 17920 25780 17926 25832
rect 17954 25780 17960 25832
rect 18012 25780 18018 25832
rect 18141 25823 18199 25829
rect 18141 25789 18153 25823
rect 18187 25820 18199 25823
rect 18892 25820 18920 25916
rect 19426 25848 19432 25900
rect 19484 25888 19490 25900
rect 20070 25888 20076 25900
rect 19484 25860 20076 25888
rect 19484 25848 19490 25860
rect 20070 25848 20076 25860
rect 20128 25888 20134 25900
rect 20165 25891 20223 25897
rect 20165 25888 20177 25891
rect 20128 25860 20177 25888
rect 20128 25848 20134 25860
rect 20165 25857 20177 25860
rect 20211 25857 20223 25891
rect 20165 25851 20223 25857
rect 20257 25891 20315 25897
rect 20257 25857 20269 25891
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 18187 25792 18920 25820
rect 20272 25820 20300 25851
rect 20346 25848 20352 25900
rect 20404 25848 20410 25900
rect 20530 25848 20536 25900
rect 20588 25848 20594 25900
rect 21192 25897 21220 25928
rect 22204 25928 23428 25956
rect 21177 25891 21235 25897
rect 21177 25857 21189 25891
rect 21223 25888 21235 25891
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 21223 25860 21833 25888
rect 21223 25857 21235 25860
rect 21177 25851 21235 25857
rect 21821 25857 21833 25860
rect 21867 25857 21879 25891
rect 22005 25891 22063 25897
rect 22005 25888 22017 25891
rect 21821 25851 21879 25857
rect 21928 25860 22017 25888
rect 21928 25832 21956 25860
rect 22005 25857 22017 25860
rect 22051 25857 22063 25891
rect 22005 25851 22063 25857
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22204 25888 22232 25928
rect 23400 25900 23428 25928
rect 26694 25916 26700 25968
rect 26752 25956 26758 25968
rect 28169 25959 28227 25965
rect 28169 25956 28181 25959
rect 26752 25928 28181 25956
rect 26752 25916 26758 25928
rect 28169 25925 28181 25928
rect 28215 25925 28227 25959
rect 29825 25959 29883 25965
rect 29825 25956 29837 25959
rect 29394 25928 29837 25956
rect 28169 25919 28227 25925
rect 29825 25925 29837 25928
rect 29871 25925 29883 25959
rect 29825 25919 29883 25925
rect 22152 25860 22232 25888
rect 22281 25891 22339 25897
rect 22152 25848 22158 25860
rect 22281 25857 22293 25891
rect 22327 25857 22339 25891
rect 22281 25851 22339 25857
rect 20438 25820 20444 25832
rect 20272 25792 20444 25820
rect 18187 25789 18199 25792
rect 18141 25783 18199 25789
rect 20438 25780 20444 25792
rect 20496 25820 20502 25832
rect 20809 25823 20867 25829
rect 20809 25820 20821 25823
rect 20496 25792 20821 25820
rect 20496 25780 20502 25792
rect 20809 25789 20821 25792
rect 20855 25789 20867 25823
rect 20809 25783 20867 25789
rect 14001 25755 14059 25761
rect 14001 25721 14013 25755
rect 14047 25721 14059 25755
rect 20824 25752 20852 25783
rect 21266 25780 21272 25832
rect 21324 25780 21330 25832
rect 21910 25780 21916 25832
rect 21968 25820 21974 25832
rect 22296 25820 22324 25851
rect 23382 25848 23388 25900
rect 23440 25848 23446 25900
rect 29914 25848 29920 25900
rect 29972 25888 29978 25900
rect 30576 25888 30604 25984
rect 30650 25916 30656 25968
rect 30708 25956 30714 25968
rect 34057 25959 34115 25965
rect 34057 25956 34069 25959
rect 30708 25928 31524 25956
rect 33626 25928 34069 25956
rect 30708 25916 30714 25928
rect 31496 25897 31524 25928
rect 34057 25925 34069 25928
rect 34103 25925 34115 25959
rect 34057 25919 34115 25925
rect 31021 25891 31079 25897
rect 31021 25888 31033 25891
rect 29972 25860 30144 25888
rect 30576 25860 31033 25888
rect 29972 25848 29978 25860
rect 27893 25823 27951 25829
rect 27893 25820 27905 25823
rect 21968 25792 22324 25820
rect 27724 25792 27905 25820
rect 21968 25780 21974 25792
rect 22370 25752 22376 25764
rect 14001 25715 14059 25721
rect 14108 25724 19012 25752
rect 20824 25724 22376 25752
rect 14108 25684 14136 25724
rect 18984 25696 19012 25724
rect 22370 25712 22376 25724
rect 22428 25712 22434 25764
rect 27724 25696 27752 25792
rect 27893 25789 27905 25792
rect 27939 25789 27951 25823
rect 27893 25783 27951 25789
rect 30116 25696 30144 25860
rect 31021 25857 31033 25860
rect 31067 25857 31079 25891
rect 31021 25851 31079 25857
rect 31481 25891 31539 25897
rect 31481 25857 31493 25891
rect 31527 25857 31539 25891
rect 31481 25851 31539 25857
rect 31665 25891 31723 25897
rect 31665 25857 31677 25891
rect 31711 25857 31723 25891
rect 31665 25851 31723 25857
rect 31113 25823 31171 25829
rect 31113 25789 31125 25823
rect 31159 25820 31171 25823
rect 31573 25823 31631 25829
rect 31573 25820 31585 25823
rect 31159 25792 31585 25820
rect 31159 25789 31171 25792
rect 31113 25783 31171 25789
rect 31573 25789 31585 25792
rect 31619 25789 31631 25823
rect 31573 25783 31631 25789
rect 31680 25752 31708 25851
rect 34146 25848 34152 25900
rect 34204 25888 34210 25900
rect 34425 25891 34483 25897
rect 34425 25888 34437 25891
rect 34204 25860 34437 25888
rect 34204 25848 34210 25860
rect 34425 25857 34437 25860
rect 34471 25888 34483 25891
rect 34701 25891 34759 25897
rect 34701 25888 34713 25891
rect 34471 25860 34713 25888
rect 34471 25857 34483 25860
rect 34425 25851 34483 25857
rect 34701 25857 34713 25860
rect 34747 25857 34759 25891
rect 34701 25851 34759 25857
rect 32122 25780 32128 25832
rect 32180 25780 32186 25832
rect 32398 25780 32404 25832
rect 32456 25780 32462 25832
rect 31588 25724 31708 25752
rect 31588 25696 31616 25724
rect 13648 25656 14136 25684
rect 9953 25647 10011 25653
rect 14642 25644 14648 25696
rect 14700 25644 14706 25696
rect 15102 25644 15108 25696
rect 15160 25644 15166 25696
rect 16298 25644 16304 25696
rect 16356 25644 16362 25696
rect 17126 25644 17132 25696
rect 17184 25644 17190 25696
rect 18966 25644 18972 25696
rect 19024 25644 19030 25696
rect 20714 25644 20720 25696
rect 20772 25644 20778 25696
rect 26878 25644 26884 25696
rect 26936 25684 26942 25696
rect 27706 25684 27712 25696
rect 26936 25656 27712 25684
rect 26936 25644 26942 25656
rect 27706 25644 27712 25656
rect 27764 25644 27770 25696
rect 30098 25644 30104 25696
rect 30156 25684 30162 25696
rect 30193 25687 30251 25693
rect 30193 25684 30205 25687
rect 30156 25656 30205 25684
rect 30156 25644 30162 25656
rect 30193 25653 30205 25656
rect 30239 25653 30251 25687
rect 30193 25647 30251 25653
rect 31570 25644 31576 25696
rect 31628 25644 31634 25696
rect 1104 25594 35248 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 35248 25594
rect 1104 25520 35248 25542
rect 5445 25483 5503 25489
rect 5445 25449 5457 25483
rect 5491 25480 5503 25483
rect 5902 25480 5908 25492
rect 5491 25452 5908 25480
rect 5491 25449 5503 25452
rect 5445 25443 5503 25449
rect 5902 25440 5908 25452
rect 5960 25440 5966 25492
rect 8294 25440 8300 25492
rect 8352 25480 8358 25492
rect 8389 25483 8447 25489
rect 8389 25480 8401 25483
rect 8352 25452 8401 25480
rect 8352 25440 8358 25452
rect 8389 25449 8401 25452
rect 8435 25449 8447 25483
rect 8389 25443 8447 25449
rect 10686 25440 10692 25492
rect 10744 25440 10750 25492
rect 16114 25440 16120 25492
rect 16172 25440 16178 25492
rect 16485 25483 16543 25489
rect 16485 25449 16497 25483
rect 16531 25480 16543 25483
rect 16758 25480 16764 25492
rect 16531 25452 16764 25480
rect 16531 25449 16543 25452
rect 16485 25443 16543 25449
rect 16758 25440 16764 25452
rect 16816 25440 16822 25492
rect 18230 25440 18236 25492
rect 18288 25440 18294 25492
rect 18966 25440 18972 25492
rect 19024 25440 19030 25492
rect 20254 25440 20260 25492
rect 20312 25480 20318 25492
rect 20441 25483 20499 25489
rect 20441 25480 20453 25483
rect 20312 25452 20453 25480
rect 20312 25440 20318 25452
rect 20441 25449 20453 25452
rect 20487 25449 20499 25483
rect 20441 25443 20499 25449
rect 21266 25440 21272 25492
rect 21324 25480 21330 25492
rect 21729 25483 21787 25489
rect 21729 25480 21741 25483
rect 21324 25452 21741 25480
rect 21324 25440 21330 25452
rect 21729 25449 21741 25452
rect 21775 25449 21787 25483
rect 21729 25443 21787 25449
rect 22370 25440 22376 25492
rect 22428 25440 22434 25492
rect 23109 25483 23167 25489
rect 23109 25449 23121 25483
rect 23155 25480 23167 25483
rect 23382 25480 23388 25492
rect 23155 25452 23388 25480
rect 23155 25449 23167 25452
rect 23109 25443 23167 25449
rect 23382 25440 23388 25452
rect 23440 25440 23446 25492
rect 26421 25483 26479 25489
rect 26421 25449 26433 25483
rect 26467 25480 26479 25483
rect 26878 25480 26884 25492
rect 26467 25452 26884 25480
rect 26467 25449 26479 25452
rect 26421 25443 26479 25449
rect 5534 25372 5540 25424
rect 5592 25372 5598 25424
rect 10704 25412 10732 25440
rect 14737 25415 14795 25421
rect 14737 25412 14749 25415
rect 10704 25384 14749 25412
rect 14737 25381 14749 25384
rect 14783 25412 14795 25415
rect 15654 25412 15660 25424
rect 14783 25384 15660 25412
rect 14783 25381 14795 25384
rect 14737 25375 14795 25381
rect 15654 25372 15660 25384
rect 15712 25372 15718 25424
rect 16132 25412 16160 25440
rect 16393 25415 16451 25421
rect 16393 25412 16405 25415
rect 16132 25384 16405 25412
rect 16393 25381 16405 25384
rect 16439 25381 16451 25415
rect 16393 25375 16451 25381
rect 5353 25347 5411 25353
rect 5353 25344 5365 25347
rect 5184 25316 5365 25344
rect 2133 25143 2191 25149
rect 2133 25109 2145 25143
rect 2179 25140 2191 25143
rect 2866 25140 2872 25152
rect 2179 25112 2872 25140
rect 2179 25109 2191 25112
rect 2133 25103 2191 25109
rect 2866 25100 2872 25112
rect 2924 25100 2930 25152
rect 3602 25100 3608 25152
rect 3660 25140 3666 25152
rect 3973 25143 4031 25149
rect 3973 25140 3985 25143
rect 3660 25112 3985 25140
rect 3660 25100 3666 25112
rect 3973 25109 3985 25112
rect 4019 25109 4031 25143
rect 3973 25103 4031 25109
rect 4154 25100 4160 25152
rect 4212 25140 4218 25152
rect 5074 25140 5080 25152
rect 4212 25112 5080 25140
rect 4212 25100 4218 25112
rect 5074 25100 5080 25112
rect 5132 25140 5138 25152
rect 5184 25149 5212 25316
rect 5353 25313 5365 25316
rect 5399 25313 5411 25347
rect 5552 25344 5580 25372
rect 11057 25347 11115 25353
rect 5552 25316 5672 25344
rect 5353 25307 5411 25313
rect 5644 25285 5672 25316
rect 11057 25313 11069 25347
rect 11103 25344 11115 25347
rect 11238 25344 11244 25356
rect 11103 25316 11244 25344
rect 11103 25313 11115 25316
rect 11057 25307 11115 25313
rect 11238 25304 11244 25316
rect 11296 25304 11302 25356
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25344 11943 25347
rect 12894 25344 12900 25356
rect 11931 25316 12900 25344
rect 11931 25313 11943 25316
rect 11885 25307 11943 25313
rect 12894 25304 12900 25316
rect 12952 25304 12958 25356
rect 12986 25304 12992 25356
rect 13044 25304 13050 25356
rect 16574 25304 16580 25356
rect 16632 25344 16638 25356
rect 18248 25344 18276 25440
rect 20809 25415 20867 25421
rect 20809 25381 20821 25415
rect 20855 25412 20867 25415
rect 22186 25412 22192 25424
rect 20855 25384 22192 25412
rect 20855 25381 20867 25384
rect 20809 25375 20867 25381
rect 22186 25372 22192 25384
rect 22244 25372 22250 25424
rect 24949 25415 25007 25421
rect 24949 25381 24961 25415
rect 24995 25381 25007 25415
rect 24949 25375 25007 25381
rect 16632 25316 18276 25344
rect 16632 25304 16638 25316
rect 20070 25304 20076 25356
rect 20128 25304 20134 25356
rect 20901 25347 20959 25353
rect 20901 25344 20913 25347
rect 20272 25316 20913 25344
rect 5537 25279 5595 25285
rect 5537 25245 5549 25279
rect 5583 25245 5595 25279
rect 5537 25239 5595 25245
rect 5629 25279 5687 25285
rect 5629 25245 5641 25279
rect 5675 25245 5687 25279
rect 5629 25239 5687 25245
rect 5169 25143 5227 25149
rect 5169 25140 5181 25143
rect 5132 25112 5181 25140
rect 5132 25100 5138 25112
rect 5169 25109 5181 25112
rect 5215 25109 5227 25143
rect 5552 25140 5580 25239
rect 11146 25236 11152 25288
rect 11204 25236 11210 25288
rect 12069 25279 12127 25285
rect 12069 25245 12081 25279
rect 12115 25245 12127 25279
rect 12069 25239 12127 25245
rect 10321 25211 10379 25217
rect 10321 25177 10333 25211
rect 10367 25208 10379 25211
rect 11054 25208 11060 25220
rect 10367 25180 11060 25208
rect 10367 25177 10379 25180
rect 10321 25171 10379 25177
rect 11054 25168 11060 25180
rect 11112 25168 11118 25220
rect 12084 25208 12112 25239
rect 12434 25236 12440 25288
rect 12492 25236 12498 25288
rect 14550 25236 14556 25288
rect 14608 25276 14614 25288
rect 15565 25279 15623 25285
rect 15565 25276 15577 25279
rect 14608 25248 15577 25276
rect 14608 25236 14614 25248
rect 15565 25245 15577 25248
rect 15611 25276 15623 25279
rect 16022 25276 16028 25288
rect 15611 25248 16028 25276
rect 15611 25245 15623 25248
rect 15565 25239 15623 25245
rect 16022 25236 16028 25248
rect 16080 25236 16086 25288
rect 16298 25236 16304 25288
rect 16356 25236 16362 25288
rect 18785 25279 18843 25285
rect 18785 25245 18797 25279
rect 18831 25276 18843 25279
rect 18874 25276 18880 25288
rect 18831 25248 18880 25276
rect 18831 25245 18843 25248
rect 18785 25239 18843 25245
rect 18874 25236 18880 25248
rect 18932 25236 18938 25288
rect 18969 25279 19027 25285
rect 18969 25245 18981 25279
rect 19015 25276 19027 25279
rect 19334 25276 19340 25288
rect 19015 25248 19340 25276
rect 19015 25245 19027 25248
rect 18969 25239 19027 25245
rect 19334 25236 19340 25248
rect 19392 25236 19398 25288
rect 12526 25208 12532 25220
rect 12084 25180 12532 25208
rect 12526 25168 12532 25180
rect 12584 25168 12590 25220
rect 15194 25168 15200 25220
rect 15252 25208 15258 25220
rect 16316 25208 16344 25236
rect 15252 25180 16344 25208
rect 20088 25208 20116 25304
rect 20272 25288 20300 25316
rect 20901 25313 20913 25316
rect 20947 25313 20959 25347
rect 20901 25307 20959 25313
rect 22204 25316 22784 25344
rect 20254 25236 20260 25288
rect 20312 25236 20318 25288
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 20714 25276 20720 25288
rect 20671 25248 20720 25276
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 20714 25236 20720 25248
rect 20772 25236 20778 25288
rect 21910 25236 21916 25288
rect 21968 25276 21974 25288
rect 22204 25285 22232 25316
rect 22756 25285 22784 25316
rect 23382 25304 23388 25356
rect 23440 25344 23446 25356
rect 24489 25347 24547 25353
rect 24489 25344 24501 25347
rect 23440 25316 24501 25344
rect 23440 25304 23446 25316
rect 24489 25313 24501 25316
rect 24535 25313 24547 25347
rect 24964 25344 24992 25375
rect 25317 25347 25375 25353
rect 25317 25344 25329 25347
rect 24964 25316 25329 25344
rect 24489 25307 24547 25313
rect 25317 25313 25329 25316
rect 25363 25313 25375 25347
rect 25317 25307 25375 25313
rect 25777 25347 25835 25353
rect 25777 25313 25789 25347
rect 25823 25313 25835 25347
rect 25777 25307 25835 25313
rect 22189 25279 22247 25285
rect 21968 25248 21993 25276
rect 21968 25236 21974 25248
rect 22189 25245 22201 25279
rect 22235 25245 22247 25279
rect 22189 25239 22247 25245
rect 22281 25279 22339 25285
rect 22281 25245 22293 25279
rect 22327 25245 22339 25279
rect 22281 25239 22339 25245
rect 22649 25279 22707 25285
rect 22649 25245 22661 25279
rect 22695 25245 22707 25279
rect 22649 25239 22707 25245
rect 22741 25279 22799 25285
rect 22741 25245 22753 25279
rect 22787 25276 22799 25279
rect 23198 25276 23204 25288
rect 22787 25248 23204 25276
rect 22787 25245 22799 25248
rect 22741 25239 22799 25245
rect 21928 25208 21956 25236
rect 22296 25208 22324 25239
rect 20088 25180 22324 25208
rect 22664 25208 22692 25239
rect 23198 25236 23204 25248
rect 23256 25276 23262 25288
rect 23293 25279 23351 25285
rect 23293 25276 23305 25279
rect 23256 25248 23305 25276
rect 23256 25236 23262 25248
rect 23293 25245 23305 25248
rect 23339 25245 23351 25279
rect 23293 25239 23351 25245
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25276 23535 25279
rect 23934 25276 23940 25288
rect 23523 25248 23940 25276
rect 23523 25245 23535 25248
rect 23477 25239 23535 25245
rect 23492 25208 23520 25239
rect 23934 25236 23940 25248
rect 23992 25236 23998 25288
rect 24578 25236 24584 25288
rect 24636 25236 24642 25288
rect 25406 25236 25412 25288
rect 25464 25236 25470 25288
rect 22664 25180 23520 25208
rect 25792 25208 25820 25307
rect 26528 25285 26556 25452
rect 26878 25440 26884 25452
rect 26936 25440 26942 25492
rect 32398 25480 32404 25492
rect 31726 25452 32404 25480
rect 31205 25415 31263 25421
rect 31205 25381 31217 25415
rect 31251 25412 31263 25415
rect 31726 25412 31754 25452
rect 32398 25440 32404 25452
rect 32456 25440 32462 25492
rect 31251 25384 31754 25412
rect 31251 25381 31263 25384
rect 31205 25375 31263 25381
rect 28261 25347 28319 25353
rect 28261 25313 28273 25347
rect 28307 25344 28319 25347
rect 28307 25316 30880 25344
rect 28307 25313 28319 25316
rect 28261 25307 28319 25313
rect 30852 25288 30880 25316
rect 30926 25304 30932 25356
rect 30984 25304 30990 25356
rect 34057 25347 34115 25353
rect 34057 25313 34069 25347
rect 34103 25313 34115 25347
rect 34057 25307 34115 25313
rect 26513 25279 26571 25285
rect 26513 25245 26525 25279
rect 26559 25245 26571 25279
rect 26513 25239 26571 25245
rect 30834 25236 30840 25288
rect 30892 25236 30898 25288
rect 34072 25220 34100 25307
rect 34330 25236 34336 25288
rect 34388 25236 34394 25288
rect 26789 25211 26847 25217
rect 26789 25208 26801 25211
rect 25792 25180 26801 25208
rect 15252 25168 15258 25180
rect 5626 25140 5632 25152
rect 5552 25112 5632 25140
rect 5169 25103 5227 25109
rect 5626 25100 5632 25112
rect 5684 25100 5690 25152
rect 14366 25100 14372 25152
rect 14424 25100 14430 25152
rect 15105 25143 15163 25149
rect 15105 25109 15117 25143
rect 15151 25140 15163 25143
rect 16114 25140 16120 25152
rect 15151 25112 16120 25140
rect 15151 25109 15163 25112
rect 15105 25103 15163 25109
rect 16114 25100 16120 25112
rect 16172 25100 16178 25152
rect 16209 25143 16267 25149
rect 16209 25109 16221 25143
rect 16255 25140 16267 25143
rect 16758 25140 16764 25152
rect 16255 25112 16764 25140
rect 16255 25109 16267 25112
rect 16209 25103 16267 25109
rect 16758 25100 16764 25112
rect 16816 25100 16822 25152
rect 17497 25143 17555 25149
rect 17497 25109 17509 25143
rect 17543 25140 17555 25143
rect 17678 25140 17684 25152
rect 17543 25112 17684 25140
rect 17543 25109 17555 25112
rect 17497 25103 17555 25109
rect 17678 25100 17684 25112
rect 17736 25140 17742 25152
rect 17954 25140 17960 25152
rect 17736 25112 17960 25140
rect 17736 25100 17742 25112
rect 17954 25100 17960 25112
rect 18012 25100 18018 25152
rect 22097 25143 22155 25149
rect 22097 25109 22109 25143
rect 22143 25140 22155 25143
rect 22664 25140 22692 25180
rect 26789 25177 26801 25180
rect 26835 25177 26847 25211
rect 26789 25171 26847 25177
rect 27798 25168 27804 25220
rect 27856 25168 27862 25220
rect 34054 25168 34060 25220
rect 34112 25168 34118 25220
rect 22143 25112 22692 25140
rect 32033 25143 32091 25149
rect 22143 25109 22155 25112
rect 22097 25103 22155 25109
rect 32033 25109 32045 25143
rect 32079 25140 32091 25143
rect 32122 25140 32128 25152
rect 32079 25112 32128 25140
rect 32079 25109 32091 25112
rect 32033 25103 32091 25109
rect 32122 25100 32128 25112
rect 32180 25140 32186 25152
rect 32398 25140 32404 25152
rect 32180 25112 32404 25140
rect 32180 25100 32186 25112
rect 32398 25100 32404 25112
rect 32456 25100 32462 25152
rect 1104 25050 35236 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 35236 25050
rect 1104 24976 35236 24998
rect 11146 24896 11152 24948
rect 11204 24896 11210 24948
rect 11238 24896 11244 24948
rect 11296 24936 11302 24948
rect 11517 24939 11575 24945
rect 11517 24936 11529 24939
rect 11296 24908 11529 24936
rect 11296 24896 11302 24908
rect 11517 24905 11529 24908
rect 11563 24905 11575 24939
rect 11517 24899 11575 24905
rect 12345 24939 12403 24945
rect 12345 24905 12357 24939
rect 12391 24936 12403 24939
rect 12434 24936 12440 24948
rect 12391 24908 12440 24936
rect 12391 24905 12403 24908
rect 12345 24899 12403 24905
rect 12434 24896 12440 24908
rect 12492 24896 12498 24948
rect 12526 24896 12532 24948
rect 12584 24896 12590 24948
rect 14550 24896 14556 24948
rect 14608 24896 14614 24948
rect 14918 24896 14924 24948
rect 14976 24896 14982 24948
rect 15378 24896 15384 24948
rect 15436 24896 15442 24948
rect 16574 24896 16580 24948
rect 16632 24936 16638 24948
rect 16669 24939 16727 24945
rect 16669 24936 16681 24939
rect 16632 24908 16681 24936
rect 16632 24896 16638 24908
rect 16669 24905 16681 24908
rect 16715 24905 16727 24939
rect 16669 24899 16727 24905
rect 17126 24896 17132 24948
rect 17184 24936 17190 24948
rect 17184 24908 22094 24936
rect 17184 24896 17190 24908
rect 3970 24828 3976 24880
rect 4028 24868 4034 24880
rect 5994 24868 6000 24880
rect 4028 24840 4936 24868
rect 4028 24828 4034 24840
rect 934 24760 940 24812
rect 992 24800 998 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 992 24772 1409 24800
rect 992 24760 998 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 3881 24803 3939 24809
rect 3881 24769 3893 24803
rect 3927 24800 3939 24803
rect 3988 24800 4016 24828
rect 3927 24772 4016 24800
rect 3927 24769 3939 24772
rect 3881 24763 3939 24769
rect 4062 24760 4068 24812
rect 4120 24760 4126 24812
rect 4157 24803 4215 24809
rect 4157 24769 4169 24803
rect 4203 24769 4215 24803
rect 4157 24763 4215 24769
rect 4080 24732 4108 24760
rect 3436 24704 4108 24732
rect 3436 24673 3464 24704
rect 3421 24667 3479 24673
rect 3421 24633 3433 24667
rect 3467 24633 3479 24667
rect 4172 24664 4200 24763
rect 4246 24760 4252 24812
rect 4304 24760 4310 24812
rect 4614 24760 4620 24812
rect 4672 24800 4678 24812
rect 4801 24803 4859 24809
rect 4801 24800 4813 24803
rect 4672 24772 4813 24800
rect 4672 24760 4678 24772
rect 4801 24769 4813 24772
rect 4847 24769 4859 24803
rect 4908 24800 4936 24840
rect 5460 24840 6000 24868
rect 5350 24800 5356 24812
rect 4908 24772 5356 24800
rect 4801 24763 4859 24769
rect 5350 24760 5356 24772
rect 5408 24800 5414 24812
rect 5460 24800 5488 24840
rect 5994 24828 6000 24840
rect 6052 24828 6058 24880
rect 9398 24828 9404 24880
rect 9456 24828 9462 24880
rect 10686 24828 10692 24880
rect 10744 24868 10750 24880
rect 10744 24840 11560 24868
rect 10744 24828 10750 24840
rect 5408 24772 5488 24800
rect 5408 24760 5414 24772
rect 5534 24760 5540 24812
rect 5592 24800 5598 24812
rect 5813 24803 5871 24809
rect 5813 24800 5825 24803
rect 5592 24772 5825 24800
rect 5592 24760 5598 24772
rect 5813 24769 5825 24772
rect 5859 24769 5871 24803
rect 5813 24763 5871 24769
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6549 24803 6607 24809
rect 6549 24800 6561 24803
rect 5960 24772 6561 24800
rect 5960 24760 5966 24772
rect 6549 24769 6561 24772
rect 6595 24769 6607 24803
rect 6549 24763 6607 24769
rect 7926 24760 7932 24812
rect 7984 24760 7990 24812
rect 8294 24760 8300 24812
rect 8352 24800 8358 24812
rect 8389 24803 8447 24809
rect 8389 24800 8401 24803
rect 8352 24772 8401 24800
rect 8352 24760 8358 24772
rect 8389 24769 8401 24772
rect 8435 24769 8447 24803
rect 10321 24803 10379 24809
rect 10321 24800 10333 24803
rect 8389 24763 8447 24769
rect 9876 24772 10333 24800
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24732 4583 24735
rect 4709 24735 4767 24741
rect 4709 24732 4721 24735
rect 4571 24704 4721 24732
rect 4571 24701 4583 24704
rect 4525 24695 4583 24701
rect 4709 24701 4721 24704
rect 4755 24701 4767 24735
rect 4709 24695 4767 24701
rect 5718 24692 5724 24744
rect 5776 24692 5782 24744
rect 6181 24735 6239 24741
rect 6181 24701 6193 24735
rect 6227 24732 6239 24735
rect 6825 24735 6883 24741
rect 6825 24732 6837 24735
rect 6227 24704 6500 24732
rect 6227 24701 6239 24704
rect 6181 24695 6239 24701
rect 6472 24664 6500 24704
rect 6656 24704 6837 24732
rect 6656 24664 6684 24704
rect 6825 24701 6837 24704
rect 6871 24701 6883 24735
rect 8665 24735 8723 24741
rect 8665 24732 8677 24735
rect 6825 24695 6883 24701
rect 8496 24704 8677 24732
rect 8496 24664 8524 24704
rect 8665 24701 8677 24704
rect 8711 24701 8723 24735
rect 8665 24695 8723 24701
rect 4172 24636 4752 24664
rect 3421 24627 3479 24633
rect 4724 24608 4752 24636
rect 5184 24636 6316 24664
rect 6472 24636 6684 24664
rect 7852 24636 8524 24664
rect 1578 24556 1584 24608
rect 1636 24556 1642 24608
rect 3602 24556 3608 24608
rect 3660 24596 3666 24608
rect 3697 24599 3755 24605
rect 3697 24596 3709 24599
rect 3660 24568 3709 24596
rect 3660 24556 3666 24568
rect 3697 24565 3709 24568
rect 3743 24565 3755 24599
rect 3697 24559 3755 24565
rect 4706 24556 4712 24608
rect 4764 24556 4770 24608
rect 5184 24605 5212 24636
rect 5169 24599 5227 24605
rect 5169 24565 5181 24599
rect 5215 24565 5227 24599
rect 6288 24596 6316 24636
rect 7852 24596 7880 24636
rect 6288 24568 7880 24596
rect 8297 24599 8355 24605
rect 5169 24559 5227 24565
rect 8297 24565 8309 24599
rect 8343 24596 8355 24599
rect 9876 24596 9904 24772
rect 10321 24769 10333 24772
rect 10367 24769 10379 24803
rect 10321 24763 10379 24769
rect 11057 24803 11115 24809
rect 11057 24769 11069 24803
rect 11103 24800 11115 24803
rect 11146 24800 11152 24812
rect 11103 24772 11152 24800
rect 11103 24769 11115 24772
rect 11057 24763 11115 24769
rect 11146 24760 11152 24772
rect 11204 24760 11210 24812
rect 11241 24803 11299 24809
rect 11241 24769 11253 24803
rect 11287 24800 11299 24803
rect 11422 24800 11428 24812
rect 11287 24772 11428 24800
rect 11287 24769 11299 24772
rect 11241 24763 11299 24769
rect 10873 24735 10931 24741
rect 10873 24701 10885 24735
rect 10919 24732 10931 24735
rect 11256 24732 11284 24763
rect 11422 24760 11428 24772
rect 11480 24760 11486 24812
rect 11532 24809 11560 24840
rect 11992 24840 12664 24868
rect 11517 24803 11575 24809
rect 11517 24769 11529 24803
rect 11563 24769 11575 24803
rect 11517 24763 11575 24769
rect 11698 24760 11704 24812
rect 11756 24760 11762 24812
rect 10919 24704 11284 24732
rect 10919 24701 10931 24704
rect 10873 24695 10931 24701
rect 11992 24608 12020 24840
rect 12158 24760 12164 24812
rect 12216 24760 12222 24812
rect 12342 24760 12348 24812
rect 12400 24760 12406 24812
rect 12434 24760 12440 24812
rect 12492 24800 12498 24812
rect 12636 24809 12664 24840
rect 15010 24828 15016 24880
rect 15068 24868 15074 24880
rect 15562 24877 15568 24880
rect 15289 24871 15347 24877
rect 15068 24837 15132 24868
rect 15068 24828 15071 24837
rect 12621 24803 12679 24809
rect 12492 24772 12572 24800
rect 12492 24760 12498 24772
rect 12544 24732 12572 24772
rect 12621 24769 12633 24803
rect 12667 24800 12679 24803
rect 13725 24803 13783 24809
rect 13725 24800 13737 24803
rect 12667 24772 13737 24800
rect 12667 24769 12679 24772
rect 12621 24763 12679 24769
rect 13725 24769 13737 24772
rect 13771 24769 13783 24803
rect 13725 24763 13783 24769
rect 14182 24760 14188 24812
rect 14240 24800 14246 24812
rect 14645 24803 14703 24809
rect 14645 24800 14657 24803
rect 14240 24772 14657 24800
rect 14240 24760 14246 24772
rect 14645 24769 14657 24772
rect 14691 24769 14703 24803
rect 14645 24763 14703 24769
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 15059 24803 15071 24828
rect 15105 24806 15132 24837
rect 15289 24837 15301 24871
rect 15335 24837 15347 24871
rect 15289 24831 15347 24837
rect 15549 24871 15568 24877
rect 15549 24837 15561 24871
rect 15549 24831 15568 24837
rect 15105 24803 15117 24806
rect 15059 24797 15117 24803
rect 15304 24732 15332 24831
rect 15562 24828 15568 24831
rect 15620 24828 15626 24880
rect 15654 24828 15660 24880
rect 15712 24868 15718 24880
rect 15749 24871 15807 24877
rect 15749 24868 15761 24871
rect 15712 24840 15761 24868
rect 15712 24828 15718 24840
rect 15749 24837 15761 24840
rect 15795 24837 15807 24871
rect 17218 24868 17224 24880
rect 15749 24831 15807 24837
rect 16868 24840 17224 24868
rect 16390 24760 16396 24812
rect 16448 24800 16454 24812
rect 16868 24809 16896 24840
rect 17218 24828 17224 24840
rect 17276 24868 17282 24880
rect 17497 24871 17555 24877
rect 17497 24868 17509 24871
rect 17276 24840 17509 24868
rect 17276 24828 17282 24840
rect 17497 24837 17509 24840
rect 17543 24837 17555 24871
rect 17497 24831 17555 24837
rect 18616 24840 19104 24868
rect 16853 24803 16911 24809
rect 16853 24800 16865 24803
rect 16448 24772 16865 24800
rect 16448 24760 16454 24772
rect 16853 24769 16865 24772
rect 16899 24769 16911 24803
rect 16853 24763 16911 24769
rect 16945 24803 17003 24809
rect 16945 24769 16957 24803
rect 16991 24769 17003 24803
rect 16945 24763 17003 24769
rect 16758 24732 16764 24744
rect 12544 24704 12940 24732
rect 12912 24673 12940 24704
rect 14476 24704 15332 24732
rect 15396 24704 16764 24732
rect 14476 24676 14504 24704
rect 12897 24667 12955 24673
rect 12897 24633 12909 24667
rect 12943 24664 12955 24667
rect 13357 24667 13415 24673
rect 13357 24664 13369 24667
rect 12943 24636 13369 24664
rect 12943 24633 12955 24636
rect 12897 24627 12955 24633
rect 13357 24633 13369 24636
rect 13403 24664 13415 24667
rect 14458 24664 14464 24676
rect 13403 24636 14464 24664
rect 13403 24633 13415 24636
rect 13357 24627 13415 24633
rect 14458 24624 14464 24636
rect 14516 24624 14522 24676
rect 14829 24667 14887 24673
rect 14829 24633 14841 24667
rect 14875 24664 14887 24667
rect 15194 24664 15200 24676
rect 14875 24636 15200 24664
rect 14875 24633 14887 24636
rect 14829 24627 14887 24633
rect 15194 24624 15200 24636
rect 15252 24624 15258 24676
rect 8343 24568 9904 24596
rect 8343 24565 8355 24568
rect 8297 24559 8355 24565
rect 10134 24556 10140 24608
rect 10192 24556 10198 24608
rect 11974 24556 11980 24608
rect 12032 24556 12038 24608
rect 13538 24556 13544 24608
rect 13596 24596 13602 24608
rect 14090 24596 14096 24608
rect 13596 24568 14096 24596
rect 13596 24556 13602 24568
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14642 24556 14648 24608
rect 14700 24596 14706 24608
rect 15105 24599 15163 24605
rect 15105 24596 15117 24599
rect 14700 24568 15117 24596
rect 14700 24556 14706 24568
rect 15105 24565 15117 24568
rect 15151 24596 15163 24599
rect 15396 24596 15424 24704
rect 16758 24692 16764 24704
rect 16816 24732 16822 24744
rect 16960 24732 16988 24763
rect 17034 24760 17040 24812
rect 17092 24760 17098 24812
rect 18230 24760 18236 24812
rect 18288 24800 18294 24812
rect 18616 24809 18644 24840
rect 18601 24803 18659 24809
rect 18601 24800 18613 24803
rect 18288 24772 18613 24800
rect 18288 24760 18294 24772
rect 18601 24769 18613 24772
rect 18647 24769 18659 24803
rect 18601 24763 18659 24769
rect 18782 24760 18788 24812
rect 18840 24760 18846 24812
rect 19076 24809 19104 24840
rect 18877 24803 18935 24809
rect 18877 24769 18889 24803
rect 18923 24769 18935 24803
rect 18877 24763 18935 24769
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24800 19119 24803
rect 19337 24803 19395 24809
rect 19337 24800 19349 24803
rect 19107 24772 19349 24800
rect 19107 24769 19119 24772
rect 19061 24763 19119 24769
rect 19337 24769 19349 24772
rect 19383 24769 19395 24803
rect 22066 24800 22094 24908
rect 23198 24896 23204 24948
rect 23256 24896 23262 24948
rect 23934 24896 23940 24948
rect 23992 24896 23998 24948
rect 24578 24896 24584 24948
rect 24636 24896 24642 24948
rect 25317 24939 25375 24945
rect 25317 24905 25329 24939
rect 25363 24936 25375 24939
rect 25406 24936 25412 24948
rect 25363 24908 25412 24936
rect 25363 24905 25375 24908
rect 25317 24899 25375 24905
rect 25406 24896 25412 24908
rect 25464 24896 25470 24948
rect 30466 24896 30472 24948
rect 30524 24896 30530 24948
rect 30926 24896 30932 24948
rect 30984 24936 30990 24948
rect 31205 24939 31263 24945
rect 31205 24936 31217 24939
rect 30984 24908 31217 24936
rect 30984 24896 30990 24908
rect 31205 24905 31217 24908
rect 31251 24905 31263 24939
rect 31205 24899 31263 24905
rect 34149 24939 34207 24945
rect 34149 24905 34161 24939
rect 34195 24936 34207 24939
rect 34330 24936 34336 24948
rect 34195 24908 34336 24936
rect 34195 24905 34207 24908
rect 34149 24899 34207 24905
rect 34330 24896 34336 24908
rect 34388 24896 34394 24948
rect 23492 24840 24624 24868
rect 23382 24800 23388 24812
rect 22066 24772 23388 24800
rect 19337 24763 19395 24769
rect 18417 24735 18475 24741
rect 18417 24732 18429 24735
rect 16816 24704 16988 24732
rect 18340 24704 18429 24732
rect 16816 24692 16822 24704
rect 16114 24624 16120 24676
rect 16172 24624 16178 24676
rect 17221 24667 17279 24673
rect 17221 24664 17233 24667
rect 16408 24636 17233 24664
rect 15151 24568 15424 24596
rect 15151 24565 15163 24568
rect 15105 24559 15163 24565
rect 15470 24556 15476 24608
rect 15528 24596 15534 24608
rect 16408 24605 16436 24636
rect 17221 24633 17233 24636
rect 17267 24633 17279 24667
rect 17221 24627 17279 24633
rect 18340 24608 18368 24704
rect 18417 24701 18429 24704
rect 18463 24732 18475 24735
rect 18892 24732 18920 24763
rect 23382 24760 23388 24772
rect 23440 24760 23446 24812
rect 23492 24741 23520 24840
rect 23615 24803 23673 24809
rect 23615 24769 23627 24803
rect 23661 24800 23673 24803
rect 23934 24800 23940 24812
rect 23661 24772 23940 24800
rect 23661 24769 23673 24772
rect 23615 24763 23673 24769
rect 23934 24760 23940 24772
rect 23992 24800 23998 24812
rect 24228 24809 24256 24840
rect 24121 24803 24179 24809
rect 24121 24800 24133 24803
rect 23992 24772 24133 24800
rect 23992 24760 23998 24772
rect 24121 24769 24133 24772
rect 24167 24769 24179 24803
rect 24121 24763 24179 24769
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 24305 24803 24363 24809
rect 24305 24769 24317 24803
rect 24351 24800 24363 24803
rect 24351 24772 24440 24800
rect 24351 24769 24363 24772
rect 24305 24763 24363 24769
rect 18463 24704 18552 24732
rect 18463 24701 18475 24704
rect 18417 24695 18475 24701
rect 18524 24664 18552 24704
rect 18800 24704 18920 24732
rect 23477 24735 23535 24741
rect 18800 24664 18828 24704
rect 23477 24701 23489 24735
rect 23523 24701 23535 24735
rect 23477 24695 23535 24701
rect 23753 24735 23811 24741
rect 23753 24701 23765 24735
rect 23799 24701 23811 24735
rect 23753 24695 23811 24701
rect 23845 24735 23903 24741
rect 23845 24701 23857 24735
rect 23891 24732 23903 24735
rect 24026 24732 24032 24744
rect 23891 24704 24032 24732
rect 23891 24701 23903 24704
rect 23845 24695 23903 24701
rect 18524 24636 18828 24664
rect 18874 24624 18880 24676
rect 18932 24664 18938 24676
rect 18969 24667 19027 24673
rect 18969 24664 18981 24667
rect 18932 24636 18981 24664
rect 18932 24624 18938 24636
rect 18969 24633 18981 24636
rect 19015 24633 19027 24667
rect 18969 24627 19027 24633
rect 19242 24624 19248 24676
rect 19300 24664 19306 24676
rect 21542 24664 21548 24676
rect 19300 24636 21548 24664
rect 19300 24624 19306 24636
rect 21542 24624 21548 24636
rect 21600 24624 21606 24676
rect 23492 24664 23520 24695
rect 23216 24636 23520 24664
rect 23768 24664 23796 24695
rect 24026 24692 24032 24704
rect 24084 24692 24090 24744
rect 24412 24732 24440 24772
rect 24486 24760 24492 24812
rect 24544 24760 24550 24812
rect 24596 24809 24624 24840
rect 24688 24840 25268 24868
rect 24581 24803 24639 24809
rect 24581 24769 24593 24803
rect 24627 24769 24639 24803
rect 24581 24763 24639 24769
rect 24688 24732 24716 24840
rect 25240 24812 25268 24840
rect 30852 24840 31064 24868
rect 24765 24803 24823 24809
rect 24765 24769 24777 24803
rect 24811 24769 24823 24803
rect 24765 24763 24823 24769
rect 25133 24803 25191 24809
rect 25133 24769 25145 24803
rect 25179 24769 25191 24803
rect 25133 24763 25191 24769
rect 24412 24704 24716 24732
rect 24504 24664 24532 24704
rect 23768 24636 24532 24664
rect 23216 24608 23244 24636
rect 15565 24599 15623 24605
rect 15565 24596 15577 24599
rect 15528 24568 15577 24596
rect 15528 24556 15534 24568
rect 15565 24565 15577 24568
rect 15611 24596 15623 24599
rect 16393 24599 16451 24605
rect 16393 24596 16405 24599
rect 15611 24568 16405 24596
rect 15611 24565 15623 24568
rect 15565 24559 15623 24565
rect 16393 24565 16405 24568
rect 16439 24565 16451 24599
rect 16393 24559 16451 24565
rect 18230 24556 18236 24608
rect 18288 24556 18294 24608
rect 18322 24556 18328 24608
rect 18380 24556 18386 24608
rect 19610 24556 19616 24608
rect 19668 24596 19674 24608
rect 23106 24596 23112 24608
rect 19668 24568 23112 24596
rect 19668 24556 19674 24568
rect 23106 24556 23112 24568
rect 23164 24556 23170 24608
rect 23198 24556 23204 24608
rect 23256 24556 23262 24608
rect 23934 24556 23940 24608
rect 23992 24596 23998 24608
rect 24780 24596 24808 24763
rect 24854 24692 24860 24744
rect 24912 24732 24918 24744
rect 25148 24732 25176 24763
rect 25222 24760 25228 24812
rect 25280 24800 25286 24812
rect 25317 24803 25375 24809
rect 25317 24800 25329 24803
rect 25280 24772 25329 24800
rect 25280 24760 25286 24772
rect 25317 24769 25329 24772
rect 25363 24769 25375 24803
rect 25317 24763 25375 24769
rect 26602 24760 26608 24812
rect 26660 24800 26666 24812
rect 30852 24809 30880 24840
rect 26973 24803 27031 24809
rect 26973 24800 26985 24803
rect 26660 24772 26985 24800
rect 26660 24760 26666 24772
rect 26973 24769 26985 24772
rect 27019 24800 27031 24803
rect 28997 24803 29055 24809
rect 28997 24800 29009 24803
rect 27019 24772 29009 24800
rect 27019 24769 27031 24772
rect 26973 24763 27031 24769
rect 28997 24769 29009 24772
rect 29043 24769 29055 24803
rect 28997 24763 29055 24769
rect 30837 24803 30895 24809
rect 30837 24769 30849 24803
rect 30883 24769 30895 24803
rect 30837 24763 30895 24769
rect 30929 24803 30987 24809
rect 30929 24769 30941 24803
rect 30975 24769 30987 24803
rect 30929 24763 30987 24769
rect 24912 24704 25176 24732
rect 30745 24735 30803 24741
rect 24912 24692 24918 24704
rect 30745 24701 30757 24735
rect 30791 24732 30803 24735
rect 30944 24732 30972 24763
rect 30791 24704 30972 24732
rect 30791 24701 30803 24704
rect 30745 24695 30803 24701
rect 23992 24568 24808 24596
rect 23992 24556 23998 24568
rect 27338 24556 27344 24608
rect 27396 24596 27402 24608
rect 28261 24599 28319 24605
rect 28261 24596 28273 24599
rect 27396 24568 28273 24596
rect 27396 24556 27402 24568
rect 28261 24565 28273 24568
rect 28307 24565 28319 24599
rect 28261 24559 28319 24565
rect 30650 24556 30656 24608
rect 30708 24596 30714 24608
rect 30760 24596 30788 24695
rect 31036 24673 31064 24840
rect 33778 24760 33784 24812
rect 33836 24760 33842 24812
rect 31205 24735 31263 24741
rect 31205 24701 31217 24735
rect 31251 24732 31263 24735
rect 31570 24732 31576 24744
rect 31251 24704 31576 24732
rect 31251 24701 31263 24704
rect 31205 24695 31263 24701
rect 31570 24692 31576 24704
rect 31628 24692 31634 24744
rect 32401 24735 32459 24741
rect 32401 24701 32413 24735
rect 32447 24701 32459 24735
rect 32401 24695 32459 24701
rect 31021 24667 31079 24673
rect 31021 24633 31033 24667
rect 31067 24664 31079 24667
rect 31067 24636 31708 24664
rect 31067 24633 31079 24636
rect 31021 24627 31079 24633
rect 31680 24608 31708 24636
rect 32416 24608 32444 24695
rect 32674 24692 32680 24744
rect 32732 24692 32738 24744
rect 30708 24568 30788 24596
rect 30708 24556 30714 24568
rect 30834 24556 30840 24608
rect 30892 24556 30898 24608
rect 31570 24556 31576 24608
rect 31628 24556 31634 24608
rect 31662 24556 31668 24608
rect 31720 24556 31726 24608
rect 31941 24599 31999 24605
rect 31941 24565 31953 24599
rect 31987 24596 31999 24599
rect 32398 24596 32404 24608
rect 31987 24568 32404 24596
rect 31987 24565 31999 24568
rect 31941 24559 31999 24565
rect 32398 24556 32404 24568
rect 32456 24556 32462 24608
rect 33318 24556 33324 24608
rect 33376 24596 33382 24608
rect 34146 24596 34152 24608
rect 33376 24568 34152 24596
rect 33376 24556 33382 24568
rect 34146 24556 34152 24568
rect 34204 24596 34210 24608
rect 34425 24599 34483 24605
rect 34425 24596 34437 24599
rect 34204 24568 34437 24596
rect 34204 24556 34210 24568
rect 34425 24565 34437 24568
rect 34471 24565 34483 24599
rect 34425 24559 34483 24565
rect 1104 24506 35248 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 35248 24506
rect 1104 24432 35248 24454
rect 2038 24392 2044 24404
rect 1596 24364 2044 24392
rect 1394 24216 1400 24268
rect 1452 24256 1458 24268
rect 1596 24265 1624 24364
rect 2038 24352 2044 24364
rect 2096 24392 2102 24404
rect 3602 24392 3608 24404
rect 2096 24364 3608 24392
rect 2096 24352 2102 24364
rect 3602 24352 3608 24364
rect 3660 24352 3666 24404
rect 4525 24395 4583 24401
rect 4525 24361 4537 24395
rect 4571 24392 4583 24395
rect 4614 24392 4620 24404
rect 4571 24364 4620 24392
rect 4571 24361 4583 24364
rect 4525 24355 4583 24361
rect 4614 24352 4620 24364
rect 4672 24352 4678 24404
rect 5350 24352 5356 24404
rect 5408 24392 5414 24404
rect 5537 24395 5595 24401
rect 5537 24392 5549 24395
rect 5408 24364 5549 24392
rect 5408 24352 5414 24364
rect 5537 24361 5549 24364
rect 5583 24361 5595 24395
rect 5537 24355 5595 24361
rect 5718 24352 5724 24404
rect 5776 24352 5782 24404
rect 7926 24352 7932 24404
rect 7984 24392 7990 24404
rect 9033 24395 9091 24401
rect 9033 24392 9045 24395
rect 7984 24364 9045 24392
rect 7984 24352 7990 24364
rect 9033 24361 9045 24364
rect 9079 24361 9091 24395
rect 9033 24355 9091 24361
rect 9398 24352 9404 24404
rect 9456 24392 9462 24404
rect 9493 24395 9551 24401
rect 9493 24392 9505 24395
rect 9456 24364 9505 24392
rect 9456 24352 9462 24364
rect 9493 24361 9505 24364
rect 9539 24361 9551 24395
rect 9493 24355 9551 24361
rect 9582 24352 9588 24404
rect 9640 24392 9646 24404
rect 10045 24395 10103 24401
rect 10045 24392 10057 24395
rect 9640 24364 10057 24392
rect 9640 24352 9646 24364
rect 10045 24361 10057 24364
rect 10091 24361 10103 24395
rect 10045 24355 10103 24361
rect 10134 24352 10140 24404
rect 10192 24352 10198 24404
rect 14737 24395 14795 24401
rect 14737 24361 14749 24395
rect 14783 24392 14795 24395
rect 14826 24392 14832 24404
rect 14783 24364 14832 24392
rect 14783 24361 14795 24364
rect 14737 24355 14795 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 15010 24352 15016 24404
rect 15068 24392 15074 24404
rect 15197 24395 15255 24401
rect 15197 24392 15209 24395
rect 15068 24364 15209 24392
rect 15068 24352 15074 24364
rect 15197 24361 15209 24364
rect 15243 24361 15255 24395
rect 15197 24355 15255 24361
rect 15473 24395 15531 24401
rect 15473 24361 15485 24395
rect 15519 24392 15531 24395
rect 15562 24392 15568 24404
rect 15519 24364 15568 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 3620 24296 4936 24324
rect 1581 24259 1639 24265
rect 1581 24256 1593 24259
rect 1452 24228 1593 24256
rect 1452 24216 1458 24228
rect 1581 24225 1593 24228
rect 1627 24225 1639 24259
rect 1581 24219 1639 24225
rect 1854 24216 1860 24268
rect 1912 24216 1918 24268
rect 3620 24265 3648 24296
rect 3605 24259 3663 24265
rect 3605 24225 3617 24259
rect 3651 24225 3663 24259
rect 4433 24259 4491 24265
rect 4433 24256 4445 24259
rect 3605 24219 3663 24225
rect 4172 24228 4445 24256
rect 4172 24200 4200 24228
rect 4433 24225 4445 24228
rect 4479 24225 4491 24259
rect 4433 24219 4491 24225
rect 4908 24200 4936 24296
rect 3973 24191 4031 24197
rect 2990 24160 3924 24188
rect 3896 24129 3924 24160
rect 3973 24157 3985 24191
rect 4019 24188 4031 24191
rect 4019 24160 4108 24188
rect 4019 24157 4031 24160
rect 3973 24151 4031 24157
rect 3881 24123 3939 24129
rect 3881 24089 3893 24123
rect 3927 24089 3939 24123
rect 3881 24083 3939 24089
rect 4080 24064 4108 24160
rect 4154 24148 4160 24200
rect 4212 24148 4218 24200
rect 4341 24191 4399 24197
rect 4341 24157 4353 24191
rect 4387 24157 4399 24191
rect 4341 24151 4399 24157
rect 4356 24120 4384 24151
rect 4890 24148 4896 24200
rect 4948 24148 4954 24200
rect 5074 24148 5080 24200
rect 5132 24188 5138 24200
rect 5132 24160 5396 24188
rect 5132 24148 5138 24160
rect 5368 24129 5396 24160
rect 5626 24148 5632 24200
rect 5684 24148 5690 24200
rect 8757 24191 8815 24197
rect 8757 24157 8769 24191
rect 8803 24188 8815 24191
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 8803 24160 9137 24188
rect 8803 24157 8815 24160
rect 8757 24151 8815 24157
rect 9125 24157 9137 24160
rect 9171 24188 9183 24191
rect 9401 24191 9459 24197
rect 9401 24188 9413 24191
rect 9171 24160 9413 24188
rect 9171 24157 9183 24160
rect 9125 24151 9183 24157
rect 9401 24157 9413 24160
rect 9447 24188 9459 24191
rect 10152 24188 10180 24352
rect 14642 24324 14648 24336
rect 13740 24296 14648 24324
rect 10597 24191 10655 24197
rect 10597 24188 10609 24191
rect 9447 24160 9904 24188
rect 10152 24160 10609 24188
rect 9447 24157 9459 24160
rect 9401 24151 9459 24157
rect 5353 24123 5411 24129
rect 4356 24092 4660 24120
rect 4632 24064 4660 24092
rect 4724 24092 5304 24120
rect 4062 24012 4068 24064
rect 4120 24012 4126 24064
rect 4614 24012 4620 24064
rect 4672 24012 4678 24064
rect 4724 24061 4752 24092
rect 4709 24055 4767 24061
rect 4709 24021 4721 24055
rect 4755 24021 4767 24055
rect 4709 24015 4767 24021
rect 5074 24012 5080 24064
rect 5132 24052 5138 24064
rect 5169 24055 5227 24061
rect 5169 24052 5181 24055
rect 5132 24024 5181 24052
rect 5132 24012 5138 24024
rect 5169 24021 5181 24024
rect 5215 24021 5227 24055
rect 5276 24052 5304 24092
rect 5353 24089 5365 24123
rect 5399 24089 5411 24123
rect 5353 24083 5411 24089
rect 5558 24055 5616 24061
rect 5558 24052 5570 24055
rect 5276 24024 5570 24052
rect 5169 24015 5227 24021
rect 5558 24021 5570 24024
rect 5604 24052 5616 24055
rect 5644 24052 5672 24148
rect 9876 24064 9904 24160
rect 10597 24157 10609 24160
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 11425 24191 11483 24197
rect 11425 24157 11437 24191
rect 11471 24188 11483 24191
rect 12069 24191 12127 24197
rect 12069 24188 12081 24191
rect 11471 24160 12081 24188
rect 11471 24157 11483 24160
rect 11425 24151 11483 24157
rect 12069 24157 12081 24160
rect 12115 24188 12127 24191
rect 12158 24188 12164 24200
rect 12115 24160 12164 24188
rect 12115 24157 12127 24160
rect 12069 24151 12127 24157
rect 12158 24148 12164 24160
rect 12216 24188 12222 24200
rect 13740 24197 13768 24296
rect 14642 24284 14648 24296
rect 14700 24284 14706 24336
rect 15488 24324 15516 24355
rect 15562 24352 15568 24364
rect 15620 24352 15626 24404
rect 16022 24352 16028 24404
rect 16080 24392 16086 24404
rect 18230 24392 18236 24404
rect 16080 24364 18236 24392
rect 16080 24352 16086 24364
rect 18230 24352 18236 24364
rect 18288 24352 18294 24404
rect 18417 24395 18475 24401
rect 18417 24361 18429 24395
rect 18463 24392 18475 24395
rect 18598 24392 18604 24404
rect 18463 24364 18604 24392
rect 18463 24361 18475 24364
rect 18417 24355 18475 24361
rect 18598 24352 18604 24364
rect 18656 24352 18662 24404
rect 19334 24352 19340 24404
rect 19392 24392 19398 24404
rect 19610 24392 19616 24404
rect 19392 24364 19616 24392
rect 19392 24352 19398 24364
rect 19610 24352 19616 24364
rect 19668 24352 19674 24404
rect 27338 24392 27344 24404
rect 19720 24364 27344 24392
rect 14936 24296 15516 24324
rect 14369 24259 14427 24265
rect 14369 24225 14381 24259
rect 14415 24256 14427 24259
rect 14415 24228 14688 24256
rect 14415 24225 14427 24228
rect 14369 24219 14427 24225
rect 12529 24191 12587 24197
rect 12529 24188 12541 24191
rect 12216 24160 12541 24188
rect 12216 24148 12222 24160
rect 12529 24157 12541 24160
rect 12575 24188 12587 24191
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 12575 24160 13737 24188
rect 12575 24157 12587 24160
rect 12529 24151 12587 24157
rect 13725 24157 13737 24160
rect 13771 24157 13783 24191
rect 13725 24151 13783 24157
rect 13906 24148 13912 24200
rect 13964 24148 13970 24200
rect 14090 24188 14096 24200
rect 14052 24160 14096 24188
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 14182 24148 14188 24200
rect 14240 24148 14246 24200
rect 14274 24148 14280 24200
rect 14332 24188 14338 24200
rect 14660 24197 14688 24228
rect 14936 24197 14964 24296
rect 15654 24284 15660 24336
rect 15712 24324 15718 24336
rect 15841 24327 15899 24333
rect 15841 24324 15853 24327
rect 15712 24296 15853 24324
rect 15712 24284 15718 24296
rect 15841 24293 15853 24296
rect 15887 24293 15899 24327
rect 15841 24287 15899 24293
rect 17037 24327 17095 24333
rect 17037 24293 17049 24327
rect 17083 24324 17095 24327
rect 17310 24324 17316 24336
rect 17083 24296 17316 24324
rect 17083 24293 17095 24296
rect 17037 24287 17095 24293
rect 17310 24284 17316 24296
rect 17368 24284 17374 24336
rect 17402 24284 17408 24336
rect 17460 24324 17466 24336
rect 19720 24324 19748 24364
rect 27338 24352 27344 24364
rect 27396 24352 27402 24404
rect 27617 24395 27675 24401
rect 27617 24361 27629 24395
rect 27663 24392 27675 24395
rect 27798 24392 27804 24404
rect 27663 24364 27804 24392
rect 27663 24361 27675 24364
rect 27617 24355 27675 24361
rect 27798 24352 27804 24364
rect 27856 24352 27862 24404
rect 31205 24395 31263 24401
rect 31205 24361 31217 24395
rect 31251 24392 31263 24395
rect 32674 24392 32680 24404
rect 31251 24364 32680 24392
rect 31251 24361 31263 24364
rect 31205 24355 31263 24361
rect 32674 24352 32680 24364
rect 32732 24352 32738 24404
rect 33505 24395 33563 24401
rect 33505 24361 33517 24395
rect 33551 24392 33563 24395
rect 33778 24392 33784 24404
rect 33551 24364 33784 24392
rect 33551 24361 33563 24364
rect 33505 24355 33563 24361
rect 33778 24352 33784 24364
rect 33836 24352 33842 24404
rect 17460 24296 19748 24324
rect 17460 24284 17466 24296
rect 20990 24284 20996 24336
rect 21048 24284 21054 24336
rect 27356 24324 27384 24352
rect 33134 24324 33140 24336
rect 27356 24296 33140 24324
rect 33134 24284 33140 24296
rect 33192 24324 33198 24336
rect 33318 24324 33324 24336
rect 33192 24296 33324 24324
rect 33192 24284 33198 24296
rect 33318 24284 33324 24296
rect 33376 24284 33382 24336
rect 16761 24259 16819 24265
rect 15396 24228 16252 24256
rect 15102 24197 15108 24200
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14332 24160 14473 24188
rect 14332 24148 14338 24160
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24188 14703 24191
rect 14921 24191 14979 24197
rect 14921 24188 14933 24191
rect 14691 24160 14933 24188
rect 14691 24157 14703 24160
rect 14645 24151 14703 24157
rect 14921 24157 14933 24160
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 15073 24191 15108 24197
rect 15073 24157 15085 24191
rect 15073 24151 15108 24157
rect 12986 24080 12992 24132
rect 13044 24120 13050 24132
rect 13173 24123 13231 24129
rect 13173 24120 13185 24123
rect 13044 24092 13185 24120
rect 13044 24080 13050 24092
rect 13173 24089 13185 24092
rect 13219 24120 13231 24123
rect 13538 24120 13544 24132
rect 13219 24092 13544 24120
rect 13219 24089 13231 24092
rect 13173 24083 13231 24089
rect 13538 24080 13544 24092
rect 13596 24080 13602 24132
rect 13817 24123 13875 24129
rect 13817 24089 13829 24123
rect 13863 24120 13875 24123
rect 14200 24120 14228 24148
rect 13863 24092 14228 24120
rect 14476 24120 14504 24151
rect 15102 24148 15108 24151
rect 15160 24148 15166 24200
rect 15396 24197 15424 24228
rect 15289 24191 15347 24197
rect 15289 24157 15301 24191
rect 15335 24188 15347 24191
rect 15381 24191 15439 24197
rect 15381 24188 15393 24191
rect 15335 24160 15393 24188
rect 15335 24157 15347 24160
rect 15289 24151 15347 24157
rect 15381 24157 15393 24160
rect 15427 24157 15439 24191
rect 15381 24151 15439 24157
rect 15562 24148 15568 24200
rect 15620 24188 15626 24200
rect 16022 24188 16028 24200
rect 15620 24160 16028 24188
rect 15620 24148 15626 24160
rect 16022 24148 16028 24160
rect 16080 24148 16086 24200
rect 16117 24123 16175 24129
rect 14476 24092 14780 24120
rect 13863 24089 13875 24092
rect 13817 24083 13875 24089
rect 5604 24024 5672 24052
rect 5604 24021 5616 24024
rect 5558 24015 5616 24021
rect 9858 24012 9864 24064
rect 9916 24012 9922 24064
rect 10505 24055 10563 24061
rect 10505 24021 10517 24055
rect 10551 24052 10563 24055
rect 11422 24052 11428 24064
rect 10551 24024 11428 24052
rect 10551 24021 10563 24024
rect 10505 24015 10563 24021
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 12526 24012 12532 24064
rect 12584 24052 12590 24064
rect 12805 24055 12863 24061
rect 12805 24052 12817 24055
rect 12584 24024 12817 24052
rect 12584 24012 12590 24024
rect 12805 24021 12817 24024
rect 12851 24052 12863 24055
rect 13906 24052 13912 24064
rect 12851 24024 13912 24052
rect 12851 24021 12863 24024
rect 12805 24015 12863 24021
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 14366 24012 14372 24064
rect 14424 24012 14430 24064
rect 14550 24012 14556 24064
rect 14608 24012 14614 24064
rect 14752 24052 14780 24092
rect 16117 24089 16129 24123
rect 16163 24089 16175 24123
rect 16117 24083 16175 24089
rect 15102 24052 15108 24064
rect 14752 24024 15108 24052
rect 15102 24012 15108 24024
rect 15160 24012 15166 24064
rect 15470 24012 15476 24064
rect 15528 24052 15534 24064
rect 16132 24052 16160 24083
rect 16224 24064 16252 24228
rect 16761 24225 16773 24259
rect 16807 24256 16819 24259
rect 17129 24259 17187 24265
rect 17129 24256 17141 24259
rect 16807 24228 17141 24256
rect 16807 24225 16819 24228
rect 16761 24219 16819 24225
rect 17129 24225 17141 24228
rect 17175 24225 17187 24259
rect 21082 24256 21088 24268
rect 17129 24219 17187 24225
rect 17236 24228 19932 24256
rect 16393 24191 16451 24197
rect 16393 24157 16405 24191
rect 16439 24188 16451 24191
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16439 24160 16681 24188
rect 16439 24157 16451 24160
rect 16393 24151 16451 24157
rect 16669 24157 16681 24160
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 17034 24148 17040 24200
rect 17092 24188 17098 24200
rect 17236 24188 17264 24228
rect 17092 24160 17264 24188
rect 17092 24148 17098 24160
rect 17310 24148 17316 24200
rect 17368 24188 17374 24200
rect 17405 24191 17463 24197
rect 17405 24188 17417 24191
rect 17368 24160 17417 24188
rect 17368 24148 17374 24160
rect 17405 24157 17417 24160
rect 17451 24157 17463 24191
rect 17405 24151 17463 24157
rect 17862 24148 17868 24200
rect 17920 24188 17926 24200
rect 18141 24191 18199 24197
rect 18141 24188 18153 24191
rect 17920 24160 18153 24188
rect 17920 24148 17926 24160
rect 18141 24157 18153 24160
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 15528 24024 16160 24052
rect 15528 24012 15534 24024
rect 16206 24012 16212 24064
rect 16264 24052 16270 24064
rect 17052 24052 17080 24148
rect 17497 24123 17555 24129
rect 17497 24120 17509 24123
rect 17144 24092 17509 24120
rect 17144 24064 17172 24092
rect 17497 24089 17509 24092
rect 17543 24089 17555 24123
rect 17497 24083 17555 24089
rect 17678 24080 17684 24132
rect 17736 24080 17742 24132
rect 18156 24120 18184 24151
rect 18322 24148 18328 24200
rect 18380 24148 18386 24200
rect 18601 24191 18659 24197
rect 18601 24157 18613 24191
rect 18647 24188 18659 24191
rect 19242 24188 19248 24200
rect 18647 24160 18828 24188
rect 18647 24157 18659 24160
rect 18601 24151 18659 24157
rect 18800 24120 18828 24160
rect 18156 24092 18828 24120
rect 18984 24160 19248 24188
rect 16264 24024 17080 24052
rect 16264 24012 16270 24024
rect 17126 24012 17132 24064
rect 17184 24012 17190 24064
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 18984 24061 19012 24160
rect 19242 24148 19248 24160
rect 19300 24148 19306 24200
rect 19444 24197 19472 24228
rect 19904 24197 19932 24228
rect 19996 24228 20392 24256
rect 19996 24200 20024 24228
rect 19429 24191 19487 24197
rect 19429 24157 19441 24191
rect 19475 24157 19487 24191
rect 19429 24151 19487 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 19978 24148 19984 24200
rect 20036 24148 20042 24200
rect 20364 24197 20392 24228
rect 20640 24228 21088 24256
rect 20640 24197 20668 24228
rect 21082 24216 21088 24228
rect 21140 24216 21146 24268
rect 23106 24216 23112 24268
rect 23164 24256 23170 24268
rect 25038 24256 25044 24268
rect 23164 24228 25044 24256
rect 23164 24216 23170 24228
rect 25038 24216 25044 24228
rect 25096 24216 25102 24268
rect 27062 24216 27068 24268
rect 27120 24256 27126 24268
rect 27433 24259 27491 24265
rect 27433 24256 27445 24259
rect 27120 24228 27445 24256
rect 27120 24216 27126 24228
rect 27433 24225 27445 24228
rect 27479 24256 27491 24259
rect 30098 24256 30104 24268
rect 27479 24228 30104 24256
rect 27479 24225 27491 24228
rect 27433 24219 27491 24225
rect 27540 24197 27568 24228
rect 30098 24216 30104 24228
rect 30156 24216 30162 24268
rect 31021 24259 31079 24265
rect 31021 24225 31033 24259
rect 31067 24256 31079 24259
rect 31481 24259 31539 24265
rect 31481 24256 31493 24259
rect 31067 24228 31493 24256
rect 31067 24225 31079 24228
rect 31021 24219 31079 24225
rect 31481 24225 31493 24228
rect 31527 24225 31539 24259
rect 31481 24219 31539 24225
rect 20349 24191 20407 24197
rect 20349 24157 20361 24191
rect 20395 24157 20407 24191
rect 20349 24151 20407 24157
rect 20625 24191 20683 24197
rect 20625 24157 20637 24191
rect 20671 24157 20683 24191
rect 20625 24151 20683 24157
rect 20717 24191 20775 24197
rect 20717 24157 20729 24191
rect 20763 24157 20775 24191
rect 20717 24151 20775 24157
rect 27525 24191 27583 24197
rect 27525 24157 27537 24191
rect 27571 24157 27583 24191
rect 30650 24188 30656 24200
rect 27525 24151 27583 24157
rect 29564 24160 30656 24188
rect 20165 24123 20223 24129
rect 20165 24089 20177 24123
rect 20211 24120 20223 24123
rect 20732 24120 20760 24151
rect 20211 24092 20760 24120
rect 20211 24089 20223 24092
rect 20165 24083 20223 24089
rect 20806 24080 20812 24132
rect 20864 24080 20870 24132
rect 20898 24080 20904 24132
rect 20956 24120 20962 24132
rect 20993 24123 21051 24129
rect 20993 24120 21005 24123
rect 20956 24092 21005 24120
rect 20956 24080 20962 24092
rect 20993 24089 21005 24092
rect 21039 24089 21051 24123
rect 20993 24083 21051 24089
rect 29564 24064 29592 24160
rect 30650 24148 30656 24160
rect 30708 24188 30714 24200
rect 30929 24191 30987 24197
rect 30929 24188 30941 24191
rect 30708 24160 30941 24188
rect 30708 24148 30714 24160
rect 30929 24157 30941 24160
rect 30975 24157 30987 24191
rect 30929 24151 30987 24157
rect 31389 24191 31447 24197
rect 31389 24157 31401 24191
rect 31435 24157 31447 24191
rect 31389 24151 31447 24157
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24188 31631 24191
rect 33336 24188 33364 24284
rect 33413 24191 33471 24197
rect 33413 24188 33425 24191
rect 31619 24160 31708 24188
rect 33336 24160 33425 24188
rect 31619 24157 31631 24160
rect 31573 24151 31631 24157
rect 31404 24120 31432 24151
rect 31680 24132 31708 24160
rect 33413 24157 33425 24160
rect 33459 24157 33471 24191
rect 33413 24151 33471 24157
rect 31404 24092 31616 24120
rect 31588 24064 31616 24092
rect 31662 24080 31668 24132
rect 31720 24080 31726 24132
rect 17313 24055 17371 24061
rect 17313 24052 17325 24055
rect 17276 24024 17325 24052
rect 17276 24012 17282 24024
rect 17313 24021 17325 24024
rect 17359 24052 17371 24055
rect 18969 24055 19027 24061
rect 18969 24052 18981 24055
rect 17359 24024 18981 24052
rect 17359 24021 17371 24024
rect 17313 24015 17371 24021
rect 18969 24021 18981 24024
rect 19015 24021 19027 24055
rect 18969 24015 19027 24021
rect 20533 24055 20591 24061
rect 20533 24021 20545 24055
rect 20579 24052 20591 24055
rect 21174 24052 21180 24064
rect 20579 24024 21180 24052
rect 20579 24021 20591 24024
rect 20533 24015 20591 24021
rect 21174 24012 21180 24024
rect 21232 24012 21238 24064
rect 29546 24012 29552 24064
rect 29604 24012 29610 24064
rect 31570 24012 31576 24064
rect 31628 24052 31634 24064
rect 31941 24055 31999 24061
rect 31941 24052 31953 24055
rect 31628 24024 31953 24052
rect 31628 24012 31634 24024
rect 31941 24021 31953 24024
rect 31987 24021 31999 24055
rect 31941 24015 31999 24021
rect 1104 23962 35236 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 35236 23962
rect 1104 23888 35236 23910
rect 1578 23808 1584 23860
rect 1636 23808 1642 23860
rect 3786 23808 3792 23860
rect 3844 23848 3850 23860
rect 4062 23848 4068 23860
rect 3844 23820 4068 23848
rect 3844 23808 3850 23820
rect 4062 23808 4068 23820
rect 4120 23848 4126 23860
rect 4982 23848 4988 23860
rect 4120 23820 4988 23848
rect 4120 23808 4126 23820
rect 4982 23808 4988 23820
rect 5040 23848 5046 23860
rect 5040 23820 6914 23848
rect 5040 23808 5046 23820
rect 1596 23780 1624 23808
rect 1673 23783 1731 23789
rect 1673 23780 1685 23783
rect 1596 23752 1685 23780
rect 1673 23749 1685 23752
rect 1719 23749 1731 23783
rect 1673 23743 1731 23749
rect 2774 23672 2780 23724
rect 2832 23672 2838 23724
rect 6362 23672 6368 23724
rect 6420 23672 6426 23724
rect 1394 23604 1400 23656
rect 1452 23604 1458 23656
rect 6886 23644 6914 23820
rect 11422 23808 11428 23860
rect 11480 23848 11486 23860
rect 12710 23848 12716 23860
rect 11480 23820 12716 23848
rect 11480 23808 11486 23820
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 14366 23848 14372 23860
rect 13188 23820 14372 23848
rect 8294 23740 8300 23792
rect 8352 23780 8358 23792
rect 8481 23783 8539 23789
rect 8481 23780 8493 23783
rect 8352 23752 8493 23780
rect 8352 23740 8358 23752
rect 8481 23749 8493 23752
rect 8527 23780 8539 23783
rect 8846 23780 8852 23792
rect 8527 23752 8852 23780
rect 8527 23749 8539 23752
rect 8481 23743 8539 23749
rect 8846 23740 8852 23752
rect 8904 23740 8910 23792
rect 9309 23783 9367 23789
rect 9309 23749 9321 23783
rect 9355 23780 9367 23783
rect 12434 23780 12440 23792
rect 9355 23752 12440 23780
rect 9355 23749 9367 23752
rect 9309 23743 9367 23749
rect 12434 23740 12440 23752
rect 12492 23740 12498 23792
rect 12621 23783 12679 23789
rect 12621 23749 12633 23783
rect 12667 23780 12679 23783
rect 12989 23783 13047 23789
rect 12989 23780 13001 23783
rect 12667 23752 13001 23780
rect 12667 23749 12679 23752
rect 12621 23743 12679 23749
rect 12989 23749 13001 23752
rect 13035 23749 13047 23783
rect 12989 23743 13047 23749
rect 9030 23672 9036 23724
rect 9088 23672 9094 23724
rect 9766 23672 9772 23724
rect 9824 23712 9830 23724
rect 12342 23712 12348 23724
rect 9824 23684 12348 23712
rect 9824 23672 9830 23684
rect 12342 23672 12348 23684
rect 12400 23712 12406 23724
rect 12529 23715 12587 23721
rect 12529 23712 12541 23715
rect 12400 23684 12541 23712
rect 12400 23672 12406 23684
rect 12529 23681 12541 23684
rect 12575 23681 12587 23715
rect 12529 23675 12587 23681
rect 12544 23644 12572 23675
rect 12710 23672 12716 23724
rect 12768 23672 12774 23724
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23712 12863 23715
rect 12894 23712 12900 23724
rect 12851 23684 12900 23712
rect 12851 23681 12863 23684
rect 12805 23675 12863 23681
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 13188 23721 13216 23820
rect 14366 23808 14372 23820
rect 14424 23808 14430 23860
rect 14550 23808 14556 23860
rect 14608 23848 14614 23860
rect 15013 23851 15071 23857
rect 15013 23848 15025 23851
rect 14608 23820 15025 23848
rect 14608 23808 14614 23820
rect 15013 23817 15025 23820
rect 15059 23817 15071 23851
rect 15013 23811 15071 23817
rect 15102 23808 15108 23860
rect 15160 23848 15166 23860
rect 15933 23851 15991 23857
rect 15933 23848 15945 23851
rect 15160 23820 15945 23848
rect 15160 23808 15166 23820
rect 13464 23752 15516 23780
rect 13081 23715 13139 23721
rect 13081 23681 13093 23715
rect 13127 23681 13139 23715
rect 13081 23675 13139 23681
rect 13173 23715 13231 23721
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13096 23644 13124 23675
rect 13464 23644 13492 23752
rect 13814 23672 13820 23724
rect 13872 23712 13878 23724
rect 14274 23712 14280 23724
rect 13872 23684 14280 23712
rect 13872 23672 13878 23684
rect 14274 23672 14280 23684
rect 14332 23672 14338 23724
rect 14550 23672 14556 23724
rect 14608 23672 14614 23724
rect 15488 23721 15516 23752
rect 15473 23715 15531 23721
rect 15473 23681 15485 23715
rect 15519 23681 15531 23715
rect 15580 23712 15608 23820
rect 15933 23817 15945 23820
rect 15979 23848 15991 23851
rect 16390 23848 16396 23860
rect 15979 23820 16396 23848
rect 15979 23817 15991 23820
rect 15933 23811 15991 23817
rect 16390 23808 16396 23820
rect 16448 23808 16454 23860
rect 20990 23808 20996 23860
rect 21048 23808 21054 23860
rect 21269 23851 21327 23857
rect 21269 23817 21281 23851
rect 21315 23848 21327 23851
rect 21634 23848 21640 23860
rect 21315 23820 21640 23848
rect 21315 23817 21327 23820
rect 21269 23811 21327 23817
rect 21634 23808 21640 23820
rect 21692 23808 21698 23860
rect 23845 23851 23903 23857
rect 22572 23820 23704 23848
rect 17126 23780 17132 23792
rect 15764 23752 17132 23780
rect 15657 23715 15715 23721
rect 15657 23712 15669 23715
rect 15580 23684 15669 23712
rect 15473 23675 15531 23681
rect 15657 23681 15669 23684
rect 15703 23681 15715 23715
rect 15657 23675 15715 23681
rect 6886 23616 12480 23644
rect 12544 23616 13492 23644
rect 13541 23647 13599 23653
rect 3145 23579 3203 23585
rect 3145 23545 3157 23579
rect 3191 23576 3203 23579
rect 4062 23576 4068 23588
rect 3191 23548 4068 23576
rect 3191 23545 3203 23548
rect 3145 23539 3203 23545
rect 4062 23536 4068 23548
rect 4120 23536 4126 23588
rect 11698 23576 11704 23588
rect 11256 23548 11704 23576
rect 11256 23520 11284 23548
rect 11698 23536 11704 23548
rect 11756 23576 11762 23588
rect 11885 23579 11943 23585
rect 11885 23576 11897 23579
rect 11756 23548 11897 23576
rect 11756 23536 11762 23548
rect 11885 23545 11897 23548
rect 11931 23545 11943 23579
rect 12452 23576 12480 23616
rect 13541 23613 13553 23647
rect 13587 23613 13599 23647
rect 13541 23607 13599 23613
rect 12618 23576 12624 23588
rect 12452 23548 12624 23576
rect 11885 23539 11943 23545
rect 12618 23536 12624 23548
rect 12676 23536 12682 23588
rect 13357 23579 13415 23585
rect 13357 23545 13369 23579
rect 13403 23576 13415 23579
rect 13556 23576 13584 23607
rect 15102 23604 15108 23656
rect 15160 23604 15166 23656
rect 15194 23604 15200 23656
rect 15252 23604 15258 23656
rect 15488 23644 15516 23675
rect 15764 23656 15792 23752
rect 17126 23740 17132 23752
rect 17184 23780 17190 23792
rect 18322 23780 18328 23792
rect 17184 23752 18328 23780
rect 17184 23740 17190 23752
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 20254 23780 20260 23792
rect 19550 23752 20260 23780
rect 20254 23740 20260 23752
rect 20312 23740 20318 23792
rect 18414 23672 18420 23724
rect 18472 23672 18478 23724
rect 18598 23672 18604 23724
rect 18656 23672 18662 23724
rect 20165 23715 20223 23721
rect 20165 23681 20177 23715
rect 20211 23712 20223 23715
rect 20438 23712 20444 23724
rect 20211 23684 20444 23712
rect 20211 23681 20223 23684
rect 20165 23675 20223 23681
rect 20438 23672 20444 23684
rect 20496 23672 20502 23724
rect 21008 23721 21036 23808
rect 21174 23740 21180 23792
rect 21232 23780 21238 23792
rect 21232 23752 21680 23780
rect 21232 23740 21238 23752
rect 20717 23715 20775 23721
rect 20717 23681 20729 23715
rect 20763 23712 20775 23715
rect 20993 23715 21051 23721
rect 20763 23684 20944 23712
rect 20763 23681 20775 23684
rect 20717 23675 20775 23681
rect 15746 23644 15752 23656
rect 15488 23616 15752 23644
rect 15746 23604 15752 23616
rect 15804 23604 15810 23656
rect 16758 23604 16764 23656
rect 16816 23644 16822 23656
rect 17310 23644 17316 23656
rect 16816 23616 17316 23644
rect 16816 23604 16822 23616
rect 17310 23604 17316 23616
rect 17368 23604 17374 23656
rect 19978 23604 19984 23656
rect 20036 23644 20042 23656
rect 20073 23647 20131 23653
rect 20073 23644 20085 23647
rect 20036 23616 20085 23644
rect 20036 23604 20042 23616
rect 20073 23613 20085 23616
rect 20119 23613 20131 23647
rect 20073 23607 20131 23613
rect 20533 23647 20591 23653
rect 20533 23613 20545 23647
rect 20579 23644 20591 23647
rect 20622 23644 20628 23656
rect 20579 23616 20628 23644
rect 20579 23613 20591 23616
rect 20533 23607 20591 23613
rect 20622 23604 20628 23616
rect 20680 23604 20686 23656
rect 20806 23604 20812 23656
rect 20864 23604 20870 23656
rect 20916 23644 20944 23684
rect 20993 23681 21005 23715
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 21085 23715 21143 23721
rect 21085 23681 21097 23715
rect 21131 23712 21143 23715
rect 21266 23712 21272 23724
rect 21131 23684 21272 23712
rect 21131 23681 21143 23684
rect 21085 23675 21143 23681
rect 21266 23672 21272 23684
rect 21324 23672 21330 23724
rect 21450 23721 21456 23724
rect 21441 23715 21456 23721
rect 21441 23681 21453 23715
rect 21441 23675 21456 23681
rect 21450 23672 21456 23675
rect 21508 23672 21514 23724
rect 21652 23721 21680 23752
rect 22572 23724 22600 23820
rect 22646 23740 22652 23792
rect 22704 23780 22710 23792
rect 23293 23783 23351 23789
rect 23293 23780 23305 23783
rect 22704 23752 23305 23780
rect 22704 23740 22710 23752
rect 23293 23749 23305 23752
rect 23339 23780 23351 23783
rect 23385 23783 23443 23789
rect 23385 23780 23397 23783
rect 23339 23752 23397 23780
rect 23339 23749 23351 23752
rect 23293 23743 23351 23749
rect 23385 23749 23397 23752
rect 23431 23749 23443 23783
rect 23385 23743 23443 23749
rect 21637 23715 21695 23721
rect 21637 23681 21649 23715
rect 21683 23712 21695 23715
rect 21821 23715 21879 23721
rect 21821 23712 21833 23715
rect 21683 23684 21833 23712
rect 21683 23681 21695 23684
rect 21637 23675 21695 23681
rect 21821 23681 21833 23684
rect 21867 23681 21879 23715
rect 21821 23675 21879 23681
rect 21910 23672 21916 23724
rect 21968 23712 21974 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21968 23684 22017 23712
rect 21968 23672 21974 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22005 23675 22063 23681
rect 22554 23672 22560 23724
rect 22612 23672 22618 23724
rect 22830 23672 22836 23724
rect 22888 23672 22894 23724
rect 22925 23715 22983 23721
rect 22925 23681 22937 23715
rect 22971 23681 22983 23715
rect 22925 23675 22983 23681
rect 20916 23616 21128 23644
rect 13403 23548 13584 23576
rect 14461 23579 14519 23585
rect 13403 23545 13415 23548
rect 13357 23539 13415 23545
rect 14461 23545 14473 23579
rect 14507 23545 14519 23579
rect 14461 23539 14519 23545
rect 3513 23511 3571 23517
rect 3513 23477 3525 23511
rect 3559 23508 3571 23511
rect 3602 23508 3608 23520
rect 3559 23480 3608 23508
rect 3559 23477 3571 23480
rect 3513 23471 3571 23477
rect 3602 23468 3608 23480
rect 3660 23468 3666 23520
rect 4617 23511 4675 23517
rect 4617 23477 4629 23511
rect 4663 23508 4675 23511
rect 5074 23508 5080 23520
rect 4663 23480 5080 23508
rect 4663 23477 4675 23480
rect 4617 23471 4675 23477
rect 5074 23468 5080 23480
rect 5132 23468 5138 23520
rect 6549 23511 6607 23517
rect 6549 23477 6561 23511
rect 6595 23508 6607 23511
rect 7006 23508 7012 23520
rect 6595 23480 7012 23508
rect 6595 23477 6607 23480
rect 6549 23471 6607 23477
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 8754 23468 8760 23520
rect 8812 23508 8818 23520
rect 8849 23511 8907 23517
rect 8849 23508 8861 23511
rect 8812 23480 8861 23508
rect 8812 23468 8818 23480
rect 8849 23477 8861 23480
rect 8895 23477 8907 23511
rect 8849 23471 8907 23477
rect 9858 23468 9864 23520
rect 9916 23508 9922 23520
rect 10594 23508 10600 23520
rect 9916 23480 10600 23508
rect 9916 23468 9922 23480
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 11238 23468 11244 23520
rect 11296 23468 11302 23520
rect 11974 23468 11980 23520
rect 12032 23508 12038 23520
rect 12345 23511 12403 23517
rect 12345 23508 12357 23511
rect 12032 23480 12357 23508
rect 12032 23468 12038 23480
rect 12345 23477 12357 23480
rect 12391 23477 12403 23511
rect 14476 23508 14504 23539
rect 14550 23536 14556 23588
rect 14608 23576 14614 23588
rect 14645 23579 14703 23585
rect 14645 23576 14657 23579
rect 14608 23548 14657 23576
rect 14608 23536 14614 23548
rect 14645 23545 14657 23548
rect 14691 23545 14703 23579
rect 14645 23539 14703 23545
rect 15010 23536 15016 23588
rect 15068 23576 15074 23588
rect 15565 23579 15623 23585
rect 15565 23576 15577 23579
rect 15068 23548 15577 23576
rect 15068 23536 15074 23548
rect 15565 23545 15577 23548
rect 15611 23545 15623 23579
rect 21100 23576 21128 23616
rect 21453 23579 21511 23585
rect 21453 23576 21465 23579
rect 15565 23539 15623 23545
rect 15672 23548 18184 23576
rect 21100 23548 21465 23576
rect 15672 23508 15700 23548
rect 14476 23480 15700 23508
rect 12345 23471 12403 23477
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 16945 23511 17003 23517
rect 16945 23508 16957 23511
rect 16908 23480 16957 23508
rect 16908 23468 16914 23480
rect 16945 23477 16957 23480
rect 16991 23508 17003 23511
rect 17678 23508 17684 23520
rect 16991 23480 17684 23508
rect 16991 23477 17003 23480
rect 16945 23471 17003 23477
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 18156 23508 18184 23548
rect 21453 23545 21465 23548
rect 21499 23545 21511 23579
rect 21453 23539 21511 23545
rect 22189 23579 22247 23585
rect 22189 23545 22201 23579
rect 22235 23576 22247 23579
rect 22848 23576 22876 23672
rect 22940 23644 22968 23675
rect 23198 23672 23204 23724
rect 23256 23672 23262 23724
rect 23676 23721 23704 23820
rect 23845 23817 23857 23851
rect 23891 23848 23903 23851
rect 23934 23848 23940 23860
rect 23891 23820 23940 23848
rect 23891 23817 23903 23820
rect 23845 23811 23903 23817
rect 23934 23808 23940 23820
rect 23992 23808 23998 23860
rect 25685 23851 25743 23857
rect 25685 23817 25697 23851
rect 25731 23848 25743 23851
rect 26878 23848 26884 23860
rect 25731 23820 26884 23848
rect 25731 23817 25743 23820
rect 25685 23811 25743 23817
rect 26878 23808 26884 23820
rect 26936 23808 26942 23860
rect 27525 23851 27583 23857
rect 27525 23817 27537 23851
rect 27571 23817 27583 23851
rect 27525 23811 27583 23817
rect 27540 23780 27568 23811
rect 29546 23808 29552 23860
rect 29604 23808 29610 23860
rect 28077 23783 28135 23789
rect 28077 23780 28089 23783
rect 27540 23752 28089 23780
rect 28077 23749 28089 23752
rect 28123 23749 28135 23783
rect 29733 23783 29791 23789
rect 29733 23780 29745 23783
rect 29302 23752 29745 23780
rect 28077 23743 28135 23749
rect 29733 23749 29745 23752
rect 29779 23749 29791 23783
rect 29733 23743 29791 23749
rect 23661 23715 23719 23721
rect 23661 23681 23673 23715
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 25317 23715 25375 23721
rect 25317 23712 25329 23715
rect 24544 23684 25329 23712
rect 24544 23672 24550 23684
rect 25317 23681 25329 23684
rect 25363 23681 25375 23715
rect 25317 23675 25375 23681
rect 26234 23672 26240 23724
rect 26292 23712 26298 23724
rect 27157 23715 27215 23721
rect 27157 23712 27169 23715
rect 26292 23684 27169 23712
rect 26292 23672 26298 23684
rect 27157 23681 27169 23684
rect 27203 23681 27215 23715
rect 27157 23675 27215 23681
rect 27706 23672 27712 23724
rect 27764 23712 27770 23724
rect 27801 23715 27859 23721
rect 27801 23712 27813 23715
rect 27764 23684 27813 23712
rect 27764 23672 27770 23684
rect 27801 23681 27813 23684
rect 27847 23681 27859 23715
rect 27801 23675 27859 23681
rect 29825 23715 29883 23721
rect 29825 23681 29837 23715
rect 29871 23712 29883 23715
rect 29871 23684 30144 23712
rect 29871 23681 29883 23684
rect 29825 23675 29883 23681
rect 23014 23644 23020 23656
rect 22940 23616 23020 23644
rect 23014 23604 23020 23616
rect 23072 23604 23078 23656
rect 23566 23604 23572 23656
rect 23624 23604 23630 23656
rect 25409 23647 25467 23653
rect 25409 23613 25421 23647
rect 25455 23644 25467 23647
rect 26142 23644 26148 23656
rect 25455 23616 26148 23644
rect 25455 23613 25467 23616
rect 25409 23607 25467 23613
rect 26142 23604 26148 23616
rect 26200 23604 26206 23656
rect 26694 23604 26700 23656
rect 26752 23604 26758 23656
rect 27065 23647 27123 23653
rect 27065 23613 27077 23647
rect 27111 23613 27123 23647
rect 27065 23607 27123 23613
rect 22235 23548 22876 23576
rect 22235 23545 22247 23548
rect 22189 23539 22247 23545
rect 24762 23536 24768 23588
rect 24820 23576 24826 23588
rect 26329 23579 26387 23585
rect 26329 23576 26341 23579
rect 24820 23548 26341 23576
rect 24820 23536 24826 23548
rect 26329 23545 26341 23548
rect 26375 23545 26387 23579
rect 26329 23539 26387 23545
rect 22922 23508 22928 23520
rect 18156 23480 22928 23508
rect 22922 23468 22928 23480
rect 22980 23468 22986 23520
rect 23106 23468 23112 23520
rect 23164 23508 23170 23520
rect 23385 23511 23443 23517
rect 23385 23508 23397 23511
rect 23164 23480 23397 23508
rect 23164 23468 23170 23480
rect 23385 23477 23397 23480
rect 23431 23477 23443 23511
rect 23385 23471 23443 23477
rect 26237 23511 26295 23517
rect 26237 23477 26249 23511
rect 26283 23508 26295 23511
rect 27080 23508 27108 23607
rect 30116 23520 30144 23684
rect 26283 23480 27108 23508
rect 26283 23477 26295 23480
rect 26237 23471 26295 23477
rect 30098 23468 30104 23520
rect 30156 23468 30162 23520
rect 1104 23418 35248 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 35248 23418
rect 1104 23344 35248 23366
rect 2317 23307 2375 23313
rect 2317 23273 2329 23307
rect 2363 23304 2375 23307
rect 2774 23304 2780 23316
rect 2363 23276 2780 23304
rect 2363 23273 2375 23276
rect 2317 23267 2375 23273
rect 2774 23264 2780 23276
rect 2832 23264 2838 23316
rect 4890 23264 4896 23316
rect 4948 23264 4954 23316
rect 6181 23307 6239 23313
rect 5000 23276 5764 23304
rect 4525 23239 4583 23245
rect 4525 23205 4537 23239
rect 4571 23236 4583 23239
rect 5000 23236 5028 23276
rect 4571 23208 5028 23236
rect 5077 23239 5135 23245
rect 4571 23205 4583 23208
rect 4525 23199 4583 23205
rect 5077 23205 5089 23239
rect 5123 23205 5135 23239
rect 5736 23236 5764 23276
rect 6181 23273 6193 23307
rect 6227 23304 6239 23307
rect 6362 23304 6368 23316
rect 6227 23276 6368 23304
rect 6227 23273 6239 23276
rect 6181 23267 6239 23273
rect 6362 23264 6368 23276
rect 6420 23264 6426 23316
rect 8481 23307 8539 23313
rect 6472 23276 8064 23304
rect 6472 23236 6500 23276
rect 5736 23208 6500 23236
rect 5077 23199 5135 23205
rect 4249 23171 4307 23177
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 4338 23168 4344 23180
rect 4295 23140 4344 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 4338 23128 4344 23140
rect 4396 23128 4402 23180
rect 5092 23168 5120 23199
rect 5261 23171 5319 23177
rect 5261 23168 5273 23171
rect 5092 23140 5273 23168
rect 5261 23137 5273 23140
rect 5307 23137 5319 23171
rect 5261 23131 5319 23137
rect 5718 23128 5724 23180
rect 5776 23128 5782 23180
rect 7006 23128 7012 23180
rect 7064 23128 7070 23180
rect 8036 23168 8064 23276
rect 8481 23273 8493 23307
rect 8527 23304 8539 23307
rect 9030 23304 9036 23316
rect 8527 23276 9036 23304
rect 8527 23273 8539 23276
rect 8481 23267 8539 23273
rect 9030 23264 9036 23276
rect 9088 23264 9094 23316
rect 11974 23264 11980 23316
rect 12032 23304 12038 23316
rect 13449 23307 13507 23313
rect 13449 23304 13461 23307
rect 12032 23276 13461 23304
rect 12032 23264 12038 23276
rect 13449 23273 13461 23276
rect 13495 23304 13507 23307
rect 13814 23304 13820 23316
rect 13495 23276 13820 23304
rect 13495 23273 13507 23276
rect 13449 23267 13507 23273
rect 13814 23264 13820 23276
rect 13872 23264 13878 23316
rect 14090 23264 14096 23316
rect 14148 23264 14154 23316
rect 14829 23307 14887 23313
rect 14829 23273 14841 23307
rect 14875 23304 14887 23307
rect 15102 23304 15108 23316
rect 14875 23276 15108 23304
rect 14875 23273 14887 23276
rect 14829 23267 14887 23273
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15654 23264 15660 23316
rect 15712 23304 15718 23316
rect 16022 23304 16028 23316
rect 15712 23276 16028 23304
rect 15712 23264 15718 23276
rect 16022 23264 16028 23276
rect 16080 23264 16086 23316
rect 18414 23264 18420 23316
rect 18472 23304 18478 23316
rect 18509 23307 18567 23313
rect 18509 23304 18521 23307
rect 18472 23276 18521 23304
rect 18472 23264 18478 23276
rect 18509 23273 18521 23276
rect 18555 23273 18567 23307
rect 18509 23267 18567 23273
rect 20165 23307 20223 23313
rect 20165 23273 20177 23307
rect 20211 23304 20223 23307
rect 20806 23304 20812 23316
rect 20211 23276 20812 23304
rect 20211 23273 20223 23276
rect 20165 23267 20223 23273
rect 20806 23264 20812 23276
rect 20864 23264 20870 23316
rect 20993 23307 21051 23313
rect 20993 23273 21005 23307
rect 21039 23304 21051 23307
rect 21082 23304 21088 23316
rect 21039 23276 21088 23304
rect 21039 23273 21051 23276
rect 20993 23267 21051 23273
rect 21082 23264 21088 23276
rect 21140 23304 21146 23316
rect 21450 23304 21456 23316
rect 21140 23276 21456 23304
rect 21140 23264 21146 23276
rect 21450 23264 21456 23276
rect 21508 23264 21514 23316
rect 22925 23307 22983 23313
rect 22925 23273 22937 23307
rect 22971 23304 22983 23307
rect 23014 23304 23020 23316
rect 22971 23276 23020 23304
rect 22971 23273 22983 23276
rect 22925 23267 22983 23273
rect 23014 23264 23020 23276
rect 23072 23304 23078 23316
rect 23566 23304 23572 23316
rect 23072 23276 23572 23304
rect 23072 23264 23078 23276
rect 23566 23264 23572 23276
rect 23624 23264 23630 23316
rect 24673 23307 24731 23313
rect 24673 23273 24685 23307
rect 24719 23304 24731 23307
rect 26234 23304 26240 23316
rect 24719 23276 26240 23304
rect 24719 23273 24731 23276
rect 24673 23267 24731 23273
rect 26234 23264 26240 23276
rect 26292 23264 26298 23316
rect 26694 23264 26700 23316
rect 26752 23304 26758 23316
rect 26789 23307 26847 23313
rect 26789 23304 26801 23307
rect 26752 23276 26801 23304
rect 26752 23264 26758 23276
rect 26789 23273 26801 23276
rect 26835 23273 26847 23307
rect 26789 23267 26847 23273
rect 27706 23264 27712 23316
rect 27764 23304 27770 23316
rect 28350 23304 28356 23316
rect 27764 23276 28356 23304
rect 27764 23264 27770 23276
rect 28350 23264 28356 23276
rect 28408 23264 28414 23316
rect 14108 23236 14136 23264
rect 15289 23239 15347 23245
rect 15289 23236 15301 23239
rect 14108 23208 15301 23236
rect 15289 23205 15301 23208
rect 15335 23236 15347 23239
rect 15470 23236 15476 23248
rect 15335 23208 15476 23236
rect 15335 23205 15347 23208
rect 15289 23199 15347 23205
rect 15470 23196 15476 23208
rect 15528 23196 15534 23248
rect 21174 23196 21180 23248
rect 21232 23236 21238 23248
rect 21361 23239 21419 23245
rect 21361 23236 21373 23239
rect 21232 23208 21373 23236
rect 21232 23196 21238 23208
rect 21361 23205 21373 23208
rect 21407 23205 21419 23239
rect 21468 23236 21496 23264
rect 24121 23239 24179 23245
rect 21468 23208 23520 23236
rect 21361 23199 21419 23205
rect 9217 23171 9275 23177
rect 9217 23168 9229 23171
rect 8036 23140 9229 23168
rect 9217 23137 9229 23140
rect 9263 23137 9275 23171
rect 9217 23131 9275 23137
rect 10689 23171 10747 23177
rect 10689 23137 10701 23171
rect 10735 23137 10747 23171
rect 10689 23131 10747 23137
rect 14185 23171 14243 23177
rect 14185 23137 14197 23171
rect 14231 23168 14243 23171
rect 15010 23168 15016 23180
rect 14231 23140 15016 23168
rect 14231 23137 14243 23140
rect 14185 23131 14243 23137
rect 2225 23103 2283 23109
rect 2225 23069 2237 23103
rect 2271 23100 2283 23103
rect 2866 23100 2872 23112
rect 2271 23072 2872 23100
rect 2271 23069 2283 23072
rect 2225 23063 2283 23069
rect 2792 22973 2820 23072
rect 2866 23060 2872 23072
rect 2924 23060 2930 23112
rect 4154 23060 4160 23112
rect 4212 23060 4218 23112
rect 5353 23103 5411 23109
rect 5353 23069 5365 23103
rect 5399 23100 5411 23103
rect 5626 23100 5632 23112
rect 5399 23072 5632 23100
rect 5399 23069 5411 23072
rect 5353 23063 5411 23069
rect 5626 23060 5632 23072
rect 5684 23060 5690 23112
rect 5810 23060 5816 23112
rect 5868 23060 5874 23112
rect 5997 23103 6055 23109
rect 5997 23069 6009 23103
rect 6043 23069 6055 23103
rect 5997 23063 6055 23069
rect 4709 23035 4767 23041
rect 4709 23001 4721 23035
rect 4755 23032 4767 23035
rect 5074 23032 5080 23044
rect 4755 23004 5080 23032
rect 4755 23001 4767 23004
rect 4709 22995 4767 23001
rect 5074 22992 5080 23004
rect 5132 22992 5138 23044
rect 5166 22992 5172 23044
rect 5224 23032 5230 23044
rect 6012 23032 6040 23063
rect 6362 23060 6368 23112
rect 6420 23100 6426 23112
rect 6733 23103 6791 23109
rect 6733 23100 6745 23103
rect 6420 23072 6745 23100
rect 6420 23060 6426 23072
rect 6733 23069 6745 23072
rect 6779 23069 6791 23103
rect 6733 23063 6791 23069
rect 8754 23060 8760 23112
rect 8812 23060 8818 23112
rect 8846 23060 8852 23112
rect 8904 23100 8910 23112
rect 8941 23103 8999 23109
rect 8941 23100 8953 23103
rect 8904 23072 8953 23100
rect 8904 23060 8910 23072
rect 8941 23069 8953 23072
rect 8987 23069 8999 23103
rect 10704 23100 10732 23131
rect 15010 23128 15016 23140
rect 15068 23128 15074 23180
rect 15562 23128 15568 23180
rect 15620 23128 15626 23180
rect 17957 23171 18015 23177
rect 17957 23137 17969 23171
rect 18003 23168 18015 23171
rect 18230 23168 18236 23180
rect 18003 23140 18236 23168
rect 18003 23137 18015 23140
rect 17957 23131 18015 23137
rect 18230 23128 18236 23140
rect 18288 23168 18294 23180
rect 18288 23140 18828 23168
rect 18288 23128 18294 23140
rect 10965 23103 11023 23109
rect 10965 23100 10977 23103
rect 10704 23072 10977 23100
rect 8941 23063 8999 23069
rect 10965 23069 10977 23072
rect 11011 23069 11023 23103
rect 10965 23063 11023 23069
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 12069 23103 12127 23109
rect 12069 23100 12081 23103
rect 11296 23072 12081 23100
rect 11296 23060 11302 23072
rect 12069 23069 12081 23072
rect 12115 23100 12127 23103
rect 12713 23103 12771 23109
rect 12713 23100 12725 23103
rect 12115 23072 12725 23100
rect 12115 23069 12127 23072
rect 12069 23063 12127 23069
rect 12713 23069 12725 23072
rect 12759 23100 12771 23103
rect 12986 23100 12992 23112
rect 12759 23072 12992 23100
rect 12759 23069 12771 23072
rect 12713 23063 12771 23069
rect 12986 23060 12992 23072
rect 13044 23060 13050 23112
rect 13372 23072 14320 23100
rect 8665 23035 8723 23041
rect 8665 23032 8677 23035
rect 5224 23004 6040 23032
rect 8234 23004 8677 23032
rect 5224 22992 5230 23004
rect 8665 23001 8677 23004
rect 8711 23001 8723 23035
rect 8665 22995 8723 23001
rect 2777 22967 2835 22973
rect 2777 22933 2789 22967
rect 2823 22964 2835 22967
rect 3418 22964 3424 22976
rect 2823 22936 3424 22964
rect 2823 22933 2835 22936
rect 2777 22927 2835 22933
rect 3418 22924 3424 22936
rect 3476 22924 3482 22976
rect 3602 22924 3608 22976
rect 3660 22964 3666 22976
rect 4062 22964 4068 22976
rect 3660 22936 4068 22964
rect 3660 22924 3666 22936
rect 4062 22924 4068 22936
rect 4120 22924 4126 22976
rect 4919 22967 4977 22973
rect 4919 22933 4931 22967
rect 4965 22964 4977 22967
rect 5258 22964 5264 22976
rect 4965 22936 5264 22964
rect 4965 22933 4977 22936
rect 4919 22927 4977 22933
rect 5258 22924 5264 22936
rect 5316 22924 5322 22976
rect 8386 22924 8392 22976
rect 8444 22964 8450 22976
rect 8772 22964 8800 23060
rect 9950 22992 9956 23044
rect 10008 22992 10014 23044
rect 11793 23035 11851 23041
rect 11793 23001 11805 23035
rect 11839 23032 11851 23035
rect 11882 23032 11888 23044
rect 11839 23004 11888 23032
rect 11839 23001 11851 23004
rect 11793 22995 11851 23001
rect 11882 22992 11888 23004
rect 11940 22992 11946 23044
rect 12253 23035 12311 23041
rect 12253 23001 12265 23035
rect 12299 23032 12311 23035
rect 12342 23032 12348 23044
rect 12299 23004 12348 23032
rect 12299 23001 12311 23004
rect 12253 22995 12311 23001
rect 12342 22992 12348 23004
rect 12400 23032 12406 23044
rect 13372 23032 13400 23072
rect 14292 23041 14320 23072
rect 14366 23060 14372 23112
rect 14424 23100 14430 23112
rect 14553 23103 14611 23109
rect 14553 23100 14565 23103
rect 14424 23072 14565 23100
rect 14424 23060 14430 23072
rect 14553 23069 14565 23072
rect 14599 23069 14611 23103
rect 14553 23063 14611 23069
rect 14645 23103 14703 23109
rect 14645 23069 14657 23103
rect 14691 23100 14703 23103
rect 15580 23100 15608 23128
rect 18524 23109 18552 23140
rect 18800 23112 18828 23140
rect 19904 23140 20668 23168
rect 14691 23072 15608 23100
rect 18509 23103 18567 23109
rect 14691 23069 14703 23072
rect 14645 23063 14703 23069
rect 18509 23069 18521 23103
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23069 18659 23103
rect 18601 23063 18659 23069
rect 12400 23004 13400 23032
rect 14277 23035 14335 23041
rect 12400 22992 12406 23004
rect 14277 23001 14289 23035
rect 14323 23001 14335 23035
rect 14277 22995 14335 23001
rect 8444 22936 8800 22964
rect 8444 22924 8450 22936
rect 12710 22924 12716 22976
rect 12768 22964 12774 22976
rect 13081 22967 13139 22973
rect 13081 22964 13093 22967
rect 12768 22936 13093 22964
rect 12768 22924 12774 22936
rect 13081 22933 13093 22936
rect 13127 22964 13139 22967
rect 13909 22967 13967 22973
rect 13909 22964 13921 22967
rect 13127 22936 13921 22964
rect 13127 22933 13139 22936
rect 13081 22927 13139 22933
rect 13909 22933 13921 22936
rect 13955 22964 13967 22967
rect 14660 22964 14688 23063
rect 18230 22992 18236 23044
rect 18288 23032 18294 23044
rect 18616 23032 18644 23063
rect 18782 23060 18788 23112
rect 18840 23060 18846 23112
rect 19904 23109 19932 23140
rect 20640 23112 20668 23140
rect 20732 23140 21036 23168
rect 19889 23103 19947 23109
rect 19889 23069 19901 23103
rect 19935 23069 19947 23103
rect 19889 23063 19947 23069
rect 20438 23060 20444 23112
rect 20496 23060 20502 23112
rect 20622 23060 20628 23112
rect 20680 23060 20686 23112
rect 20732 23109 20760 23140
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 18288 23004 18644 23032
rect 20165 23035 20223 23041
rect 18288 22992 18294 23004
rect 20165 23001 20177 23035
rect 20211 23032 20223 23035
rect 20257 23035 20315 23041
rect 20257 23032 20269 23035
rect 20211 23004 20269 23032
rect 20211 23001 20223 23004
rect 20165 22995 20223 23001
rect 20257 23001 20269 23004
rect 20303 23001 20315 23035
rect 20257 22995 20315 23001
rect 13955 22936 14688 22964
rect 17405 22967 17463 22973
rect 13955 22933 13967 22936
rect 13909 22927 13967 22933
rect 17405 22933 17417 22967
rect 17451 22964 17463 22967
rect 18506 22964 18512 22976
rect 17451 22936 18512 22964
rect 17451 22933 17463 22936
rect 17405 22927 17463 22933
rect 18506 22924 18512 22936
rect 18564 22924 18570 22976
rect 19978 22924 19984 22976
rect 20036 22964 20042 22976
rect 20732 22964 20760 23063
rect 20898 23060 20904 23112
rect 20956 23060 20962 23112
rect 20036 22936 20760 22964
rect 20809 22967 20867 22973
rect 20036 22924 20042 22936
rect 20809 22933 20821 22967
rect 20855 22964 20867 22967
rect 20916 22964 20944 23060
rect 21008 22973 21036 23140
rect 21192 23041 21220 23196
rect 22922 23128 22928 23180
rect 22980 23168 22986 23180
rect 23382 23168 23388 23180
rect 22980 23140 23388 23168
rect 22980 23128 22986 23140
rect 23382 23128 23388 23140
rect 23440 23128 23446 23180
rect 21269 23103 21327 23109
rect 21269 23069 21281 23103
rect 21315 23100 21327 23103
rect 22741 23103 22799 23109
rect 22741 23100 22753 23103
rect 21315 23072 22140 23100
rect 21315 23069 21327 23072
rect 21269 23063 21327 23069
rect 21177 23035 21235 23041
rect 21177 23001 21189 23035
rect 21223 23001 21235 23035
rect 21177 22995 21235 23001
rect 22002 22992 22008 23044
rect 22060 23032 22066 23044
rect 22112 23032 22140 23072
rect 22480 23072 22753 23100
rect 22373 23035 22431 23041
rect 22373 23032 22385 23035
rect 22060 23004 22385 23032
rect 22060 22992 22066 23004
rect 22373 23001 22385 23004
rect 22419 23001 22431 23035
rect 22373 22995 22431 23001
rect 20855 22936 20944 22964
rect 20977 22967 21036 22973
rect 20855 22933 20867 22936
rect 20809 22927 20867 22933
rect 20977 22933 20989 22967
rect 21023 22936 21036 22967
rect 21023 22933 21035 22936
rect 20977 22927 21035 22933
rect 21358 22924 21364 22976
rect 21416 22964 21422 22976
rect 22480 22964 22508 23072
rect 22741 23069 22753 23072
rect 22787 23069 22799 23103
rect 23492 23100 23520 23208
rect 24121 23205 24133 23239
rect 24167 23236 24179 23239
rect 24762 23236 24768 23248
rect 24167 23208 24768 23236
rect 24167 23205 24179 23208
rect 24121 23199 24179 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 24857 23239 24915 23245
rect 24857 23205 24869 23239
rect 24903 23236 24915 23239
rect 25222 23236 25228 23248
rect 24903 23208 25228 23236
rect 24903 23205 24915 23208
rect 24857 23199 24915 23205
rect 25222 23196 25228 23208
rect 25280 23196 25286 23248
rect 23661 23171 23719 23177
rect 23661 23137 23673 23171
rect 23707 23168 23719 23171
rect 34057 23171 34115 23177
rect 23707 23140 26188 23168
rect 23707 23137 23719 23140
rect 23661 23131 23719 23137
rect 26160 23112 26188 23140
rect 34057 23137 34069 23171
rect 34103 23168 34115 23171
rect 34103 23140 34652 23168
rect 34103 23137 34115 23140
rect 34057 23131 34115 23137
rect 23753 23103 23811 23109
rect 23753 23100 23765 23103
rect 23492 23072 23765 23100
rect 22741 23063 22799 23069
rect 23753 23069 23765 23072
rect 23799 23069 23811 23103
rect 23753 23063 23811 23069
rect 24121 23103 24179 23109
rect 24121 23069 24133 23103
rect 24167 23100 24179 23103
rect 24167 23072 24256 23100
rect 24167 23069 24179 23072
rect 24121 23063 24179 23069
rect 22557 23035 22615 23041
rect 22557 23001 22569 23035
rect 22603 23032 22615 23035
rect 23290 23032 23296 23044
rect 22603 23004 23296 23032
rect 22603 23001 22615 23004
rect 22557 22995 22615 23001
rect 23290 22992 23296 23004
rect 23348 22992 23354 23044
rect 21416 22936 22508 22964
rect 21416 22924 21422 22936
rect 22646 22924 22652 22976
rect 22704 22924 22710 22976
rect 23768 22964 23796 23063
rect 24228 23032 24256 23072
rect 24486 23060 24492 23112
rect 24544 23060 24550 23112
rect 24765 23103 24823 23109
rect 24765 23069 24777 23103
rect 24811 23100 24823 23103
rect 25130 23100 25136 23112
rect 24811 23072 25136 23100
rect 24811 23069 24823 23072
rect 24765 23063 24823 23069
rect 25130 23060 25136 23072
rect 25188 23060 25194 23112
rect 25225 23103 25283 23109
rect 25225 23069 25237 23103
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 25593 23103 25651 23109
rect 25593 23069 25605 23103
rect 25639 23069 25651 23103
rect 25593 23063 25651 23069
rect 24394 23032 24400 23044
rect 24228 23004 24400 23032
rect 24394 22992 24400 23004
rect 24452 22992 24458 23044
rect 24504 22964 24532 23060
rect 24578 22992 24584 23044
rect 24636 23032 24642 23044
rect 25240 23032 25268 23063
rect 24636 23004 25268 23032
rect 24636 22992 24642 23004
rect 25314 22964 25320 22976
rect 23768 22936 25320 22964
rect 25314 22924 25320 22936
rect 25372 22964 25378 22976
rect 25608 22964 25636 23063
rect 26050 23060 26056 23112
rect 26108 23060 26114 23112
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26421 23103 26479 23109
rect 26421 23100 26433 23103
rect 26200 23072 26433 23100
rect 26200 23060 26206 23072
rect 26421 23069 26433 23072
rect 26467 23069 26479 23103
rect 26421 23063 26479 23069
rect 26789 23103 26847 23109
rect 26789 23069 26801 23103
rect 26835 23069 26847 23103
rect 26789 23063 26847 23069
rect 26068 23032 26096 23060
rect 26804 23032 26832 23063
rect 26878 23060 26884 23112
rect 26936 23100 26942 23112
rect 26973 23103 27031 23109
rect 26973 23100 26985 23103
rect 26936 23072 26985 23100
rect 26936 23060 26942 23072
rect 26973 23069 26985 23072
rect 27019 23069 27031 23103
rect 26973 23063 27031 23069
rect 34330 23060 34336 23112
rect 34388 23060 34394 23112
rect 34624 23044 34652 23140
rect 26068 23004 26832 23032
rect 34606 22992 34612 23044
rect 34664 22992 34670 23044
rect 25372 22936 25636 22964
rect 25372 22924 25378 22936
rect 1104 22874 35236 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 35236 22874
rect 1104 22800 35236 22822
rect 4338 22720 4344 22772
rect 4396 22720 4402 22772
rect 5077 22763 5135 22769
rect 5077 22729 5089 22763
rect 5123 22760 5135 22763
rect 5166 22760 5172 22772
rect 5123 22732 5172 22760
rect 5123 22729 5135 22732
rect 5077 22723 5135 22729
rect 5166 22720 5172 22732
rect 5224 22720 5230 22772
rect 5626 22720 5632 22772
rect 5684 22720 5690 22772
rect 5718 22720 5724 22772
rect 5776 22760 5782 22772
rect 5776 22732 6684 22760
rect 5776 22720 5782 22732
rect 1762 22652 1768 22704
rect 1820 22692 1826 22704
rect 2133 22695 2191 22701
rect 2133 22692 2145 22695
rect 1820 22664 2145 22692
rect 1820 22652 1826 22664
rect 2133 22661 2145 22664
rect 2179 22661 2191 22695
rect 2133 22655 2191 22661
rect 2866 22652 2872 22704
rect 2924 22652 2930 22704
rect 3973 22695 4031 22701
rect 3973 22661 3985 22695
rect 4019 22661 4031 22695
rect 3973 22655 4031 22661
rect 4189 22695 4247 22701
rect 4189 22661 4201 22695
rect 4235 22692 4247 22695
rect 4235 22664 4660 22692
rect 4235 22661 4247 22664
rect 4189 22655 4247 22661
rect 3988 22568 4016 22655
rect 4632 22636 4660 22664
rect 4614 22584 4620 22636
rect 4672 22584 4678 22636
rect 5258 22584 5264 22636
rect 5316 22584 5322 22636
rect 5353 22627 5411 22633
rect 5353 22593 5365 22627
rect 5399 22624 5411 22627
rect 5644 22624 5672 22720
rect 6656 22701 6684 22732
rect 9950 22720 9956 22772
rect 10008 22720 10014 22772
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 21910 22760 21916 22772
rect 20772 22732 21916 22760
rect 20772 22720 20778 22732
rect 21910 22720 21916 22732
rect 21968 22720 21974 22772
rect 23290 22720 23296 22772
rect 23348 22720 23354 22772
rect 23382 22720 23388 22772
rect 23440 22760 23446 22772
rect 24121 22763 24179 22769
rect 24121 22760 24133 22763
rect 23440 22732 24133 22760
rect 23440 22720 23446 22732
rect 24121 22729 24133 22732
rect 24167 22760 24179 22763
rect 24302 22760 24308 22772
rect 24167 22732 24308 22760
rect 24167 22729 24179 22732
rect 24121 22723 24179 22729
rect 24302 22720 24308 22732
rect 24360 22720 24366 22772
rect 6641 22695 6699 22701
rect 6641 22661 6653 22695
rect 6687 22661 6699 22695
rect 8297 22695 8355 22701
rect 8297 22692 8309 22695
rect 7866 22664 8309 22692
rect 6641 22655 6699 22661
rect 8297 22661 8309 22664
rect 8343 22661 8355 22695
rect 16393 22695 16451 22701
rect 8297 22655 8355 22661
rect 8404 22664 9904 22692
rect 8404 22636 8432 22664
rect 5399 22596 5672 22624
rect 5399 22593 5411 22596
rect 5353 22587 5411 22593
rect 8386 22584 8392 22636
rect 8444 22584 8450 22636
rect 9876 22633 9904 22664
rect 16393 22661 16405 22695
rect 16439 22692 16451 22695
rect 18417 22695 18475 22701
rect 16439 22664 17908 22692
rect 16439 22661 16451 22664
rect 16393 22655 16451 22661
rect 8849 22627 8907 22633
rect 8849 22593 8861 22627
rect 8895 22593 8907 22627
rect 8849 22587 8907 22593
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 10321 22627 10379 22633
rect 10321 22624 10333 22627
rect 9907 22596 10333 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 10321 22593 10333 22596
rect 10367 22593 10379 22627
rect 10321 22587 10379 22593
rect 1857 22559 1915 22565
rect 1857 22525 1869 22559
rect 1903 22525 1915 22559
rect 1857 22519 1915 22525
rect 1872 22420 1900 22519
rect 3970 22516 3976 22568
rect 4028 22556 4034 22568
rect 5074 22556 5080 22568
rect 4028 22528 5080 22556
rect 4028 22516 4034 22528
rect 5074 22516 5080 22528
rect 5132 22516 5138 22568
rect 6362 22516 6368 22568
rect 6420 22516 6426 22568
rect 8113 22559 8171 22565
rect 8113 22525 8125 22559
rect 8159 22556 8171 22559
rect 8864 22556 8892 22587
rect 11146 22584 11152 22636
rect 11204 22624 11210 22636
rect 12069 22627 12127 22633
rect 12069 22624 12081 22627
rect 11204 22596 12081 22624
rect 11204 22584 11210 22596
rect 12069 22593 12081 22596
rect 12115 22624 12127 22627
rect 12345 22627 12403 22633
rect 12345 22624 12357 22627
rect 12115 22596 12357 22624
rect 12115 22593 12127 22596
rect 12069 22587 12127 22593
rect 12345 22593 12357 22596
rect 12391 22624 12403 22627
rect 12526 22624 12532 22636
rect 12391 22596 12532 22624
rect 12391 22593 12403 22596
rect 12345 22587 12403 22593
rect 12526 22584 12532 22596
rect 12584 22584 12590 22636
rect 15378 22584 15384 22636
rect 15436 22584 15442 22636
rect 15654 22584 15660 22636
rect 15712 22584 15718 22636
rect 16942 22584 16948 22636
rect 17000 22584 17006 22636
rect 17144 22633 17172 22664
rect 17880 22636 17908 22664
rect 18417 22661 18429 22695
rect 18463 22692 18475 22695
rect 20438 22692 20444 22704
rect 18463 22664 20444 22692
rect 18463 22661 18475 22664
rect 18417 22655 18475 22661
rect 20438 22652 20444 22664
rect 20496 22652 20502 22704
rect 22002 22652 22008 22704
rect 22060 22692 22066 22704
rect 22557 22695 22615 22701
rect 22557 22692 22569 22695
rect 22060 22664 22569 22692
rect 22060 22652 22066 22664
rect 22557 22661 22569 22664
rect 22603 22661 22615 22695
rect 23308 22692 23336 22720
rect 23308 22664 24348 22692
rect 22557 22655 22615 22661
rect 17129 22627 17187 22633
rect 17129 22593 17141 22627
rect 17175 22593 17187 22627
rect 17129 22587 17187 22593
rect 17678 22584 17684 22636
rect 17736 22584 17742 22636
rect 17862 22584 17868 22636
rect 17920 22584 17926 22636
rect 18046 22584 18052 22636
rect 18104 22584 18110 22636
rect 18230 22584 18236 22636
rect 18288 22584 18294 22636
rect 21266 22584 21272 22636
rect 21324 22624 21330 22636
rect 24320 22633 24348 22664
rect 24394 22652 24400 22704
rect 24452 22692 24458 22704
rect 24581 22695 24639 22701
rect 24581 22692 24593 22695
rect 24452 22664 24593 22692
rect 24452 22652 24458 22664
rect 24581 22661 24593 22664
rect 24627 22661 24639 22695
rect 24581 22655 24639 22661
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 21324 22596 22385 22624
rect 21324 22584 21330 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 24213 22627 24271 22633
rect 24213 22593 24225 22627
rect 24259 22593 24271 22627
rect 24213 22587 24271 22593
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22624 24363 22627
rect 24946 22624 24952 22636
rect 24351 22596 24952 22624
rect 24351 22593 24363 22596
rect 24305 22587 24363 22593
rect 8159 22528 8892 22556
rect 9401 22559 9459 22565
rect 8159 22525 8171 22528
rect 8113 22519 8171 22525
rect 9401 22525 9413 22559
rect 9447 22556 9459 22559
rect 9766 22556 9772 22568
rect 9447 22528 9772 22556
rect 9447 22525 9459 22528
rect 9401 22519 9459 22525
rect 9766 22516 9772 22528
rect 9824 22516 9830 22568
rect 12437 22559 12495 22565
rect 12437 22525 12449 22559
rect 12483 22556 12495 22559
rect 13262 22556 13268 22568
rect 12483 22528 13268 22556
rect 12483 22525 12495 22528
rect 12437 22519 12495 22525
rect 13262 22516 13268 22528
rect 13320 22516 13326 22568
rect 18248 22556 18276 22584
rect 17512 22528 18276 22556
rect 3605 22491 3663 22497
rect 3605 22457 3617 22491
rect 3651 22488 3663 22491
rect 4706 22488 4712 22500
rect 3651 22460 4712 22488
rect 3651 22457 3663 22460
rect 3605 22451 3663 22457
rect 4706 22448 4712 22460
rect 4764 22448 4770 22500
rect 5350 22488 5356 22500
rect 4816 22460 5356 22488
rect 2314 22420 2320 22432
rect 1872 22392 2320 22420
rect 2314 22380 2320 22392
rect 2372 22380 2378 22432
rect 4157 22423 4215 22429
rect 4157 22389 4169 22423
rect 4203 22420 4215 22423
rect 4816 22420 4844 22460
rect 5184 22432 5212 22460
rect 5350 22448 5356 22460
rect 5408 22448 5414 22500
rect 8846 22448 8852 22500
rect 8904 22488 8910 22500
rect 10781 22491 10839 22497
rect 10781 22488 10793 22491
rect 8904 22460 10793 22488
rect 8904 22448 8910 22460
rect 10781 22457 10793 22460
rect 10827 22457 10839 22491
rect 10781 22451 10839 22457
rect 12713 22491 12771 22497
rect 12713 22457 12725 22491
rect 12759 22488 12771 22491
rect 13814 22488 13820 22500
rect 12759 22460 13820 22488
rect 12759 22457 12771 22460
rect 12713 22451 12771 22457
rect 13814 22448 13820 22460
rect 13872 22448 13878 22500
rect 14458 22448 14464 22500
rect 14516 22488 14522 22500
rect 16850 22488 16856 22500
rect 14516 22460 16856 22488
rect 14516 22448 14522 22460
rect 15580 22432 15608 22460
rect 16850 22448 16856 22460
rect 16908 22488 16914 22500
rect 17512 22497 17540 22528
rect 22646 22516 22652 22568
rect 22704 22516 22710 22568
rect 23842 22516 23848 22568
rect 23900 22516 23906 22568
rect 24228 22556 24256 22587
rect 24946 22584 24952 22596
rect 25004 22584 25010 22636
rect 25314 22584 25320 22636
rect 25372 22584 25378 22636
rect 25409 22627 25467 22633
rect 25409 22593 25421 22627
rect 25455 22593 25467 22627
rect 25409 22587 25467 22593
rect 25424 22556 25452 22587
rect 25866 22556 25872 22568
rect 24228 22528 25872 22556
rect 17497 22491 17555 22497
rect 17497 22488 17509 22491
rect 16908 22460 17509 22488
rect 16908 22448 16914 22460
rect 17497 22457 17509 22460
rect 17543 22457 17555 22491
rect 17497 22451 17555 22457
rect 18506 22448 18512 22500
rect 18564 22448 18570 22500
rect 22664 22488 22692 22516
rect 23382 22488 23388 22500
rect 22664 22460 23388 22488
rect 23382 22448 23388 22460
rect 23440 22488 23446 22500
rect 24228 22488 24256 22528
rect 25866 22516 25872 22528
rect 25924 22516 25930 22568
rect 23440 22460 24256 22488
rect 23440 22448 23446 22460
rect 24302 22448 24308 22500
rect 24360 22488 24366 22500
rect 26050 22488 26056 22500
rect 24360 22460 26056 22488
rect 24360 22448 24366 22460
rect 26050 22448 26056 22460
rect 26108 22448 26114 22500
rect 4203 22392 4844 22420
rect 4985 22423 5043 22429
rect 4203 22389 4215 22392
rect 4157 22383 4215 22389
rect 4985 22389 4997 22423
rect 5031 22420 5043 22423
rect 5074 22420 5080 22432
rect 5031 22392 5080 22420
rect 5031 22389 5043 22392
rect 4985 22383 5043 22389
rect 5074 22380 5080 22392
rect 5132 22380 5138 22432
rect 5166 22380 5172 22432
rect 5224 22380 5230 22432
rect 14918 22380 14924 22432
rect 14976 22380 14982 22432
rect 15562 22380 15568 22432
rect 15620 22380 15626 22432
rect 17034 22380 17040 22432
rect 17092 22380 17098 22432
rect 22738 22380 22744 22432
rect 22796 22380 22802 22432
rect 23934 22380 23940 22432
rect 23992 22380 23998 22432
rect 1104 22330 35248 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 35248 22330
rect 1104 22256 35248 22278
rect 2866 22176 2872 22228
rect 2924 22216 2930 22228
rect 2961 22219 3019 22225
rect 2961 22216 2973 22219
rect 2924 22188 2973 22216
rect 2924 22176 2930 22188
rect 2961 22185 2973 22188
rect 3007 22185 3019 22219
rect 2961 22179 3019 22185
rect 3605 22219 3663 22225
rect 3605 22185 3617 22219
rect 3651 22216 3663 22219
rect 3970 22216 3976 22228
rect 3651 22188 3976 22216
rect 3651 22185 3663 22188
rect 3605 22179 3663 22185
rect 3970 22176 3976 22188
rect 4028 22216 4034 22228
rect 4522 22216 4528 22228
rect 4028 22188 4528 22216
rect 4028 22176 4034 22188
rect 4522 22176 4528 22188
rect 4580 22176 4586 22228
rect 4706 22176 4712 22228
rect 4764 22176 4770 22228
rect 4985 22219 5043 22225
rect 4985 22185 4997 22219
rect 5031 22216 5043 22219
rect 5258 22216 5264 22228
rect 5031 22188 5264 22216
rect 5031 22185 5043 22188
rect 4985 22179 5043 22185
rect 5258 22176 5264 22188
rect 5316 22176 5322 22228
rect 8297 22219 8355 22225
rect 8297 22185 8309 22219
rect 8343 22216 8355 22219
rect 8846 22216 8852 22228
rect 8343 22188 8852 22216
rect 8343 22185 8355 22188
rect 8297 22179 8355 22185
rect 4724 22148 4752 22176
rect 5350 22148 5356 22160
rect 4724 22120 5356 22148
rect 5350 22108 5356 22120
rect 5408 22108 5414 22160
rect 3142 22080 3148 22092
rect 2884 22052 3148 22080
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 2884 22021 2912 22052
rect 3142 22040 3148 22052
rect 3200 22080 3206 22092
rect 3786 22080 3792 22092
rect 3200 22052 3792 22080
rect 3200 22040 3206 22052
rect 3786 22040 3792 22052
rect 3844 22040 3850 22092
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 992 21984 1409 22012
rect 992 21972 998 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 2777 22015 2835 22021
rect 2777 21981 2789 22015
rect 2823 22012 2835 22015
rect 2869 22015 2927 22021
rect 2869 22012 2881 22015
rect 2823 21984 2881 22012
rect 2823 21981 2835 21984
rect 2777 21975 2835 21981
rect 2869 21981 2881 21984
rect 2915 21981 2927 22015
rect 2869 21975 2927 21981
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 21981 4675 22015
rect 4617 21975 4675 21981
rect 4801 22015 4859 22021
rect 4801 21981 4813 22015
rect 4847 22012 4859 22015
rect 4847 21984 5028 22012
rect 4847 21981 4859 21984
rect 4801 21975 4859 21981
rect 4632 21944 4660 21975
rect 4632 21916 4844 21944
rect 4816 21888 4844 21916
rect 5000 21888 5028 21984
rect 8312 21956 8340 22179
rect 8846 22176 8852 22188
rect 8904 22176 8910 22228
rect 14553 22219 14611 22225
rect 14553 22185 14565 22219
rect 14599 22216 14611 22219
rect 14599 22188 15240 22216
rect 14599 22185 14611 22188
rect 14553 22179 14611 22185
rect 15212 22089 15240 22188
rect 15378 22176 15384 22228
rect 15436 22176 15442 22228
rect 15654 22176 15660 22228
rect 15712 22176 15718 22228
rect 16942 22216 16948 22228
rect 16684 22188 16948 22216
rect 16393 22151 16451 22157
rect 16393 22117 16405 22151
rect 16439 22148 16451 22151
rect 16684 22148 16712 22188
rect 16942 22176 16948 22188
rect 17000 22176 17006 22228
rect 20714 22176 20720 22228
rect 20772 22176 20778 22228
rect 21269 22219 21327 22225
rect 21269 22185 21281 22219
rect 21315 22185 21327 22219
rect 21269 22179 21327 22185
rect 16439 22120 16712 22148
rect 16761 22151 16819 22157
rect 16439 22117 16451 22120
rect 16393 22111 16451 22117
rect 16761 22117 16773 22151
rect 16807 22148 16819 22151
rect 16807 22120 16896 22148
rect 16807 22117 16819 22120
rect 16761 22111 16819 22117
rect 15197 22083 15255 22089
rect 15197 22049 15209 22083
rect 15243 22080 15255 22083
rect 16868 22080 16896 22120
rect 17770 22108 17776 22160
rect 17828 22108 17834 22160
rect 18601 22151 18659 22157
rect 18601 22117 18613 22151
rect 18647 22148 18659 22151
rect 18647 22120 19472 22148
rect 18647 22117 18659 22120
rect 18601 22111 18659 22117
rect 15243 22052 15608 22080
rect 15243 22049 15255 22052
rect 15197 22043 15255 22049
rect 15580 22024 15608 22052
rect 16684 22052 16896 22080
rect 13817 22015 13875 22021
rect 13817 21981 13829 22015
rect 13863 22012 13875 22015
rect 13998 22012 14004 22024
rect 13863 21984 14004 22012
rect 13863 21981 13875 21984
rect 13817 21975 13875 21981
rect 13998 21972 14004 21984
rect 14056 22012 14062 22024
rect 14277 22015 14335 22021
rect 14277 22012 14289 22015
rect 14056 21984 14289 22012
rect 14056 21972 14062 21984
rect 14277 21981 14289 21984
rect 14323 21981 14335 22015
rect 14277 21975 14335 21981
rect 14550 21972 14556 22024
rect 14608 22012 14614 22024
rect 14645 22015 14703 22021
rect 14645 22012 14657 22015
rect 14608 21984 14657 22012
rect 14608 21972 14614 21984
rect 14645 21981 14657 21984
rect 14691 22012 14703 22015
rect 14918 22012 14924 22024
rect 14691 21984 14924 22012
rect 14691 21981 14703 21984
rect 14645 21975 14703 21981
rect 14918 21972 14924 21984
rect 14976 22012 14982 22024
rect 15289 22015 15347 22021
rect 15289 22012 15301 22015
rect 14976 21984 15301 22012
rect 14976 21972 14982 21984
rect 15289 21981 15301 21984
rect 15335 21981 15347 22015
rect 15289 21975 15347 21981
rect 15470 21972 15476 22024
rect 15528 21972 15534 22024
rect 15562 21972 15568 22024
rect 15620 21972 15626 22024
rect 15746 21972 15752 22024
rect 15804 21972 15810 22024
rect 16206 21972 16212 22024
rect 16264 21972 16270 22024
rect 16298 21972 16304 22024
rect 16356 21972 16362 22024
rect 16482 21972 16488 22024
rect 16540 21972 16546 22024
rect 16684 22021 16712 22052
rect 17034 22040 17040 22092
rect 17092 22080 17098 22092
rect 17221 22083 17279 22089
rect 17221 22080 17233 22083
rect 17092 22052 17233 22080
rect 17092 22040 17098 22052
rect 17221 22049 17233 22052
rect 17267 22049 17279 22083
rect 17221 22043 17279 22049
rect 17313 22083 17371 22089
rect 17313 22049 17325 22083
rect 17359 22080 17371 22083
rect 17788 22080 17816 22108
rect 19444 22089 19472 22120
rect 20732 22120 21128 22148
rect 18141 22083 18199 22089
rect 18141 22080 18153 22083
rect 17359 22052 18153 22080
rect 17359 22049 17371 22052
rect 17313 22043 17371 22049
rect 18141 22049 18153 22052
rect 18187 22049 18199 22083
rect 18141 22043 18199 22049
rect 19429 22083 19487 22089
rect 19429 22049 19441 22083
rect 19475 22049 19487 22083
rect 19429 22043 19487 22049
rect 16669 22015 16727 22021
rect 16669 21981 16681 22015
rect 16715 21981 16727 22015
rect 16669 21975 16727 21981
rect 16850 21972 16856 22024
rect 16908 22012 16914 22024
rect 17328 22012 17356 22043
rect 17773 22015 17831 22021
rect 16908 21984 17356 22012
rect 17512 21984 17724 22012
rect 16908 21972 16914 21984
rect 8294 21944 8300 21956
rect 7852 21916 8300 21944
rect 1578 21836 1584 21888
rect 1636 21836 1642 21888
rect 3970 21836 3976 21888
rect 4028 21876 4034 21888
rect 4157 21879 4215 21885
rect 4157 21876 4169 21879
rect 4028 21848 4169 21876
rect 4028 21836 4034 21848
rect 4157 21845 4169 21848
rect 4203 21845 4215 21879
rect 4157 21839 4215 21845
rect 4798 21836 4804 21888
rect 4856 21836 4862 21888
rect 4982 21836 4988 21888
rect 5040 21836 5046 21888
rect 6362 21836 6368 21888
rect 6420 21876 6426 21888
rect 7852 21885 7880 21916
rect 8294 21904 8300 21916
rect 8352 21904 8358 21956
rect 16025 21947 16083 21953
rect 16025 21913 16037 21947
rect 16071 21944 16083 21947
rect 17512 21944 17540 21984
rect 16071 21916 17540 21944
rect 16071 21913 16083 21916
rect 16025 21907 16083 21913
rect 17586 21904 17592 21956
rect 17644 21904 17650 21956
rect 17696 21944 17724 21984
rect 17773 21981 17785 22015
rect 17819 22012 17831 22015
rect 17862 22012 17868 22024
rect 17819 21984 17868 22012
rect 17819 21981 17831 21984
rect 17773 21975 17831 21981
rect 17862 21972 17868 21984
rect 17920 22012 17926 22024
rect 18233 22015 18291 22021
rect 18233 22012 18245 22015
rect 17920 21984 18245 22012
rect 17920 21972 17926 21984
rect 18233 21981 18245 21984
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 18690 21972 18696 22024
rect 18748 22012 18754 22024
rect 19521 22015 19579 22021
rect 19521 22012 19533 22015
rect 18748 21984 19533 22012
rect 18748 21972 18754 21984
rect 19521 21981 19533 21984
rect 19567 21981 19579 22015
rect 19521 21975 19579 21981
rect 20732 21953 20760 22120
rect 21100 22080 21128 22120
rect 21174 22108 21180 22160
rect 21232 22148 21238 22160
rect 21284 22148 21312 22179
rect 21358 22176 21364 22228
rect 21416 22216 21422 22228
rect 21453 22219 21511 22225
rect 21453 22216 21465 22219
rect 21416 22188 21465 22216
rect 21416 22176 21422 22188
rect 21453 22185 21465 22188
rect 21499 22185 21511 22219
rect 21453 22179 21511 22185
rect 22554 22176 22560 22228
rect 22612 22176 22618 22228
rect 23658 22176 23664 22228
rect 23716 22176 23722 22228
rect 23845 22219 23903 22225
rect 23845 22185 23857 22219
rect 23891 22216 23903 22219
rect 23934 22216 23940 22228
rect 23891 22188 23940 22216
rect 23891 22185 23903 22188
rect 23845 22179 23903 22185
rect 23934 22176 23940 22188
rect 23992 22176 23998 22228
rect 32566 22219 32624 22225
rect 32566 22216 32578 22219
rect 31726 22188 32578 22216
rect 21232 22120 22324 22148
rect 21232 22108 21238 22120
rect 21266 22080 21272 22092
rect 21100 22052 21272 22080
rect 21266 22040 21272 22052
rect 21324 22040 21330 22092
rect 22296 22080 22324 22120
rect 23676 22080 23704 22176
rect 22296 22052 23704 22080
rect 23952 22080 23980 22176
rect 24673 22151 24731 22157
rect 24673 22117 24685 22151
rect 24719 22148 24731 22151
rect 26142 22148 26148 22160
rect 24719 22120 26148 22148
rect 24719 22117 24731 22120
rect 24673 22111 24731 22117
rect 26142 22108 26148 22120
rect 26200 22108 26206 22160
rect 31573 22151 31631 22157
rect 31573 22117 31585 22151
rect 31619 22148 31631 22151
rect 31726 22148 31754 22188
rect 32566 22185 32578 22188
rect 32612 22185 32624 22219
rect 32566 22179 32624 22185
rect 34057 22219 34115 22225
rect 34057 22185 34069 22219
rect 34103 22216 34115 22219
rect 34330 22216 34336 22228
rect 34103 22188 34336 22216
rect 34103 22185 34115 22188
rect 34057 22179 34115 22185
rect 34330 22176 34336 22188
rect 34388 22176 34394 22228
rect 31619 22120 31754 22148
rect 31619 22117 31631 22120
rect 31573 22111 31631 22117
rect 23952 22052 24624 22080
rect 21008 22021 21128 22022
rect 20993 22015 21128 22021
rect 20993 21981 21005 22015
rect 21039 22012 21128 22015
rect 21174 22012 21180 22024
rect 21039 21994 21180 22012
rect 21039 21981 21051 21994
rect 21100 21984 21180 21994
rect 20993 21975 21051 21981
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 21284 22012 21312 22040
rect 21284 21987 21328 22012
rect 21284 21984 21373 21987
rect 21300 21981 21373 21984
rect 20717 21947 20775 21953
rect 20717 21944 20729 21947
rect 17696 21916 20729 21944
rect 20717 21913 20729 21916
rect 20763 21913 20775 21947
rect 20717 21907 20775 21913
rect 21085 21947 21143 21953
rect 21085 21913 21097 21947
rect 21131 21913 21143 21947
rect 21300 21947 21327 21981
rect 21361 21947 21373 21981
rect 21910 21972 21916 22024
rect 21968 21972 21974 22024
rect 22296 22021 22324 22052
rect 22051 22015 22109 22021
rect 22051 21990 22063 22015
rect 22020 21981 22063 21990
rect 22097 21981 22109 22015
rect 22020 21975 22109 21981
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 21981 22339 22015
rect 22281 21975 22339 21981
rect 22557 22015 22615 22021
rect 22557 21981 22569 22015
rect 22603 21981 22615 22015
rect 22557 21975 22615 21981
rect 21300 21944 21373 21947
rect 22020 21962 22094 21975
rect 22020 21944 22048 21962
rect 22186 21953 22192 21956
rect 21300 21916 22048 21944
rect 21085 21907 21143 21913
rect 22185 21907 22192 21953
rect 22244 21944 22250 21956
rect 22244 21916 22285 21944
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 6420 21848 7849 21876
rect 6420 21836 6426 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 7837 21839 7895 21845
rect 8386 21836 8392 21888
rect 8444 21876 8450 21888
rect 8573 21879 8631 21885
rect 8573 21876 8585 21879
rect 8444 21848 8585 21876
rect 8444 21836 8450 21848
rect 8573 21845 8585 21848
rect 8619 21845 8631 21879
rect 8573 21839 8631 21845
rect 9398 21836 9404 21888
rect 9456 21876 9462 21888
rect 9585 21879 9643 21885
rect 9585 21876 9597 21879
rect 9456 21848 9597 21876
rect 9456 21836 9462 21848
rect 9585 21845 9597 21848
rect 9631 21845 9643 21879
rect 9585 21839 9643 21845
rect 11606 21836 11612 21888
rect 11664 21876 11670 21888
rect 11885 21879 11943 21885
rect 11885 21876 11897 21879
rect 11664 21848 11897 21876
rect 11664 21836 11670 21848
rect 11885 21845 11897 21848
rect 11931 21876 11943 21879
rect 13173 21879 13231 21885
rect 13173 21876 13185 21879
rect 11931 21848 13185 21876
rect 11931 21845 11943 21848
rect 11885 21839 11943 21845
rect 13173 21845 13185 21848
rect 13219 21876 13231 21879
rect 13262 21876 13268 21888
rect 13219 21848 13268 21876
rect 13219 21845 13231 21848
rect 13173 21839 13231 21845
rect 13262 21836 13268 21848
rect 13320 21836 13326 21888
rect 13541 21879 13599 21885
rect 13541 21845 13553 21879
rect 13587 21876 13599 21879
rect 13630 21876 13636 21888
rect 13587 21848 13636 21876
rect 13587 21845 13599 21848
rect 13541 21839 13599 21845
rect 13630 21836 13636 21848
rect 13688 21836 13694 21888
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14093 21879 14151 21885
rect 14093 21876 14105 21879
rect 13964 21848 14105 21876
rect 13964 21836 13970 21848
rect 14093 21845 14105 21848
rect 14139 21845 14151 21879
rect 14093 21839 14151 21845
rect 16298 21836 16304 21888
rect 16356 21876 16362 21888
rect 16850 21876 16856 21888
rect 16356 21848 16856 21876
rect 16356 21836 16362 21848
rect 16850 21836 16856 21848
rect 16908 21836 16914 21888
rect 17129 21879 17187 21885
rect 17129 21845 17141 21879
rect 17175 21876 17187 21879
rect 17218 21876 17224 21888
rect 17175 21848 17224 21876
rect 17175 21845 17187 21848
rect 17129 21839 17187 21845
rect 17218 21836 17224 21848
rect 17276 21876 17282 21888
rect 17957 21879 18015 21885
rect 17957 21876 17969 21879
rect 17276 21848 17969 21876
rect 17276 21836 17282 21848
rect 17957 21845 17969 21848
rect 18003 21845 18015 21879
rect 17957 21839 18015 21845
rect 20346 21836 20352 21888
rect 20404 21836 20410 21888
rect 20898 21836 20904 21888
rect 20956 21876 20962 21888
rect 21100 21876 21128 21907
rect 22186 21904 22192 21907
rect 22244 21904 22250 21916
rect 20956 21848 21128 21876
rect 22465 21879 22523 21885
rect 20956 21836 20962 21848
rect 22465 21845 22477 21879
rect 22511 21876 22523 21879
rect 22572 21876 22600 21975
rect 22738 21972 22744 22024
rect 22796 21972 22802 22024
rect 23014 21972 23020 22024
rect 23072 21972 23078 22024
rect 23382 21972 23388 22024
rect 23440 21972 23446 22024
rect 23750 21972 23756 22024
rect 23808 22012 23814 22024
rect 24596 22021 24624 22052
rect 31110 22040 31116 22092
rect 31168 22040 31174 22092
rect 31662 22040 31668 22092
rect 31720 22040 31726 22092
rect 32306 22040 32312 22092
rect 32364 22040 32370 22092
rect 24397 22015 24455 22021
rect 24397 22012 24409 22015
rect 23808 21984 24409 22012
rect 23808 21972 23814 21984
rect 24397 21981 24409 21984
rect 24443 21981 24455 22015
rect 24397 21975 24455 21981
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 31205 22015 31263 22021
rect 31205 22012 31217 22015
rect 24581 21975 24639 21981
rect 30300 21984 31217 22012
rect 23477 21947 23535 21953
rect 23477 21913 23489 21947
rect 23523 21913 23535 21947
rect 23477 21907 23535 21913
rect 22511 21848 22600 21876
rect 22511 21845 22523 21848
rect 22465 21839 22523 21845
rect 23198 21836 23204 21888
rect 23256 21876 23262 21888
rect 23492 21876 23520 21907
rect 30300 21888 30328 21984
rect 31205 21981 31217 21984
rect 31251 22012 31263 22015
rect 31849 22015 31907 22021
rect 31849 22012 31861 22015
rect 31251 21984 31861 22012
rect 31251 21981 31263 21984
rect 31205 21975 31263 21981
rect 31849 21981 31861 21984
rect 31895 21981 31907 22015
rect 31849 21975 31907 21981
rect 32030 21904 32036 21956
rect 32088 21904 32094 21956
rect 33318 21904 33324 21956
rect 33376 21904 33382 21956
rect 23256 21848 23520 21876
rect 23256 21836 23262 21848
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 23677 21879 23735 21885
rect 23677 21876 23689 21879
rect 23624 21848 23689 21876
rect 23624 21836 23630 21848
rect 23677 21845 23689 21848
rect 23723 21845 23735 21879
rect 23677 21839 23735 21845
rect 30282 21836 30288 21888
rect 30340 21836 30346 21888
rect 1104 21786 35236 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 35236 21786
rect 1104 21712 35236 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 1636 21644 2636 21672
rect 1636 21632 1642 21644
rect 2608 21613 2636 21644
rect 4798 21632 4804 21684
rect 4856 21632 4862 21684
rect 9861 21675 9919 21681
rect 9861 21641 9873 21675
rect 9907 21672 9919 21675
rect 11146 21672 11152 21684
rect 9907 21644 11152 21672
rect 9907 21641 9919 21644
rect 9861 21635 9919 21641
rect 2593 21607 2651 21613
rect 2593 21573 2605 21607
rect 2639 21573 2651 21607
rect 2593 21567 2651 21573
rect 3326 21564 3332 21616
rect 3384 21564 3390 21616
rect 4816 21604 4844 21632
rect 4724 21576 4844 21604
rect 2314 21496 2320 21548
rect 2372 21496 2378 21548
rect 4430 21496 4436 21548
rect 4488 21496 4494 21548
rect 4614 21496 4620 21548
rect 4672 21496 4678 21548
rect 4724 21545 4752 21576
rect 7374 21564 7380 21616
rect 7432 21564 7438 21616
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21505 4767 21539
rect 4709 21499 4767 21505
rect 4801 21539 4859 21545
rect 4801 21505 4813 21539
rect 4847 21536 4859 21539
rect 4847 21508 5028 21536
rect 4847 21505 4859 21508
rect 4801 21499 4859 21505
rect 2332 21468 2360 21496
rect 5000 21480 5028 21508
rect 5350 21496 5356 21548
rect 5408 21496 5414 21548
rect 8389 21539 8447 21545
rect 8389 21505 8401 21539
rect 8435 21505 8447 21539
rect 8389 21499 8447 21505
rect 9217 21539 9275 21545
rect 9217 21505 9229 21539
rect 9263 21536 9275 21539
rect 9674 21536 9680 21548
rect 9263 21508 9680 21536
rect 9263 21505 9275 21508
rect 9217 21499 9275 21505
rect 3970 21468 3976 21480
rect 2332 21440 3976 21468
rect 3970 21428 3976 21440
rect 4028 21428 4034 21480
rect 4065 21471 4123 21477
rect 4065 21437 4077 21471
rect 4111 21468 4123 21471
rect 4982 21468 4988 21480
rect 4111 21440 4988 21468
rect 4111 21437 4123 21440
rect 4065 21431 4123 21437
rect 4982 21428 4988 21440
rect 5040 21428 5046 21480
rect 5077 21471 5135 21477
rect 5077 21437 5089 21471
rect 5123 21468 5135 21471
rect 5261 21471 5319 21477
rect 5261 21468 5273 21471
rect 5123 21440 5273 21468
rect 5123 21437 5135 21440
rect 5077 21431 5135 21437
rect 5261 21437 5273 21440
rect 5307 21437 5319 21471
rect 6362 21468 6368 21480
rect 5261 21431 5319 21437
rect 5644 21440 6368 21468
rect 3988 21400 4016 21428
rect 5644 21400 5672 21440
rect 6362 21428 6368 21440
rect 6420 21428 6426 21480
rect 6641 21471 6699 21477
rect 6641 21468 6653 21471
rect 6472 21440 6653 21468
rect 3988 21372 5672 21400
rect 5721 21403 5779 21409
rect 5721 21369 5733 21403
rect 5767 21400 5779 21403
rect 6472 21400 6500 21440
rect 6641 21437 6653 21440
rect 6687 21437 6699 21471
rect 6641 21431 6699 21437
rect 8113 21471 8171 21477
rect 8113 21437 8125 21471
rect 8159 21468 8171 21471
rect 8404 21468 8432 21499
rect 9674 21496 9680 21508
rect 9732 21536 9738 21548
rect 9968 21545 9996 21644
rect 11146 21632 11152 21644
rect 11204 21632 11210 21684
rect 11333 21675 11391 21681
rect 11333 21641 11345 21675
rect 11379 21672 11391 21675
rect 11606 21672 11612 21684
rect 11379 21644 11612 21672
rect 11379 21641 11391 21644
rect 11333 21635 11391 21641
rect 10045 21607 10103 21613
rect 10045 21573 10057 21607
rect 10091 21604 10103 21607
rect 10965 21607 11023 21613
rect 10965 21604 10977 21607
rect 10091 21576 10364 21604
rect 10091 21573 10103 21576
rect 10045 21567 10103 21573
rect 10336 21545 10364 21576
rect 10428 21576 10977 21604
rect 9953 21539 10011 21545
rect 9953 21536 9965 21539
rect 9732 21508 9965 21536
rect 9732 21496 9738 21508
rect 9953 21505 9965 21508
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21505 10195 21539
rect 10137 21499 10195 21505
rect 10321 21539 10379 21545
rect 10321 21505 10333 21539
rect 10367 21505 10379 21539
rect 10321 21499 10379 21505
rect 10152 21468 10180 21499
rect 10428 21468 10456 21576
rect 10965 21573 10977 21576
rect 11011 21604 11023 21607
rect 11238 21604 11244 21616
rect 11011 21576 11244 21604
rect 11011 21573 11023 21576
rect 10965 21567 11023 21573
rect 11238 21564 11244 21576
rect 11296 21604 11302 21616
rect 11348 21604 11376 21635
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 11974 21632 11980 21684
rect 12032 21632 12038 21684
rect 13262 21632 13268 21684
rect 13320 21672 13326 21684
rect 13446 21672 13452 21684
rect 13320 21644 13452 21672
rect 13320 21632 13326 21644
rect 13446 21632 13452 21644
rect 13504 21672 13510 21684
rect 13504 21644 14228 21672
rect 13504 21632 13510 21644
rect 14093 21607 14151 21613
rect 14093 21604 14105 21607
rect 11296 21576 11376 21604
rect 13648 21576 14105 21604
rect 11296 21564 11302 21576
rect 11514 21496 11520 21548
rect 11572 21496 11578 21548
rect 11793 21539 11851 21545
rect 11793 21505 11805 21539
rect 11839 21505 11851 21539
rect 11793 21499 11851 21505
rect 8159 21440 8432 21468
rect 9416 21440 10456 21468
rect 10597 21471 10655 21477
rect 8159 21437 8171 21440
rect 8113 21431 8171 21437
rect 5767 21372 6500 21400
rect 5767 21369 5779 21372
rect 5721 21363 5779 21369
rect 9416 21344 9444 21440
rect 10597 21437 10609 21471
rect 10643 21468 10655 21471
rect 10778 21468 10784 21480
rect 10643 21440 10784 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 10778 21428 10784 21440
rect 10836 21428 10842 21480
rect 10962 21428 10968 21480
rect 11020 21468 11026 21480
rect 11808 21468 11836 21499
rect 13262 21496 13268 21548
rect 13320 21536 13326 21548
rect 13357 21539 13415 21545
rect 13357 21536 13369 21539
rect 13320 21508 13369 21536
rect 13320 21496 13326 21508
rect 13357 21505 13369 21508
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 13449 21539 13507 21545
rect 13449 21505 13461 21539
rect 13495 21505 13507 21539
rect 13449 21499 13507 21505
rect 11020 21440 11836 21468
rect 11020 21428 11026 21440
rect 12342 21428 12348 21480
rect 12400 21468 12406 21480
rect 13464 21468 13492 21499
rect 13538 21496 13544 21548
rect 13596 21536 13602 21548
rect 13648 21545 13676 21576
rect 14093 21573 14105 21576
rect 14139 21573 14151 21607
rect 14093 21567 14151 21573
rect 13633 21539 13691 21545
rect 13633 21536 13645 21539
rect 13596 21508 13645 21536
rect 13596 21496 13602 21508
rect 13633 21505 13645 21508
rect 13679 21505 13691 21539
rect 13633 21499 13691 21505
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 13906 21536 13912 21548
rect 13771 21508 13912 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 13906 21496 13912 21508
rect 13964 21496 13970 21548
rect 13998 21496 14004 21548
rect 14056 21496 14062 21548
rect 14200 21545 14228 21644
rect 16206 21632 16212 21684
rect 16264 21632 16270 21684
rect 16482 21632 16488 21684
rect 16540 21672 16546 21684
rect 17037 21675 17095 21681
rect 17037 21672 17049 21675
rect 16540 21644 17049 21672
rect 16540 21632 16546 21644
rect 17037 21641 17049 21644
rect 17083 21641 17095 21675
rect 17037 21635 17095 21641
rect 17218 21632 17224 21684
rect 17276 21632 17282 21684
rect 17405 21675 17463 21681
rect 17405 21641 17417 21675
rect 17451 21672 17463 21675
rect 17678 21672 17684 21684
rect 17451 21644 17684 21672
rect 17451 21641 17463 21644
rect 17405 21635 17463 21641
rect 17678 21632 17684 21644
rect 17736 21672 17742 21684
rect 17954 21672 17960 21684
rect 17736 21644 17960 21672
rect 17736 21632 17742 21644
rect 17954 21632 17960 21644
rect 18012 21632 18018 21684
rect 18046 21632 18052 21684
rect 18104 21672 18110 21684
rect 18141 21675 18199 21681
rect 18141 21672 18153 21675
rect 18104 21644 18153 21672
rect 18104 21632 18110 21644
rect 18141 21641 18153 21644
rect 18187 21641 18199 21675
rect 18141 21635 18199 21641
rect 20901 21675 20959 21681
rect 20901 21641 20913 21675
rect 20947 21672 20959 21675
rect 21174 21672 21180 21684
rect 20947 21644 21180 21672
rect 20947 21641 20959 21644
rect 20901 21635 20959 21641
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 23198 21632 23204 21684
rect 23256 21672 23262 21684
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 23256 21644 23397 21672
rect 23256 21632 23262 21644
rect 23385 21641 23397 21644
rect 23431 21641 23443 21675
rect 23385 21635 23443 21641
rect 23658 21632 23664 21684
rect 23716 21632 23722 21684
rect 26789 21675 26847 21681
rect 26789 21641 26801 21675
rect 26835 21672 26847 21675
rect 26835 21644 28856 21672
rect 26835 21641 26847 21644
rect 26789 21635 26847 21641
rect 14185 21539 14243 21545
rect 14185 21505 14197 21539
rect 14231 21536 14243 21539
rect 14231 21508 15608 21536
rect 14231 21505 14243 21508
rect 14185 21499 14243 21505
rect 12400 21440 13492 21468
rect 14016 21468 14044 21496
rect 14016 21440 14412 21468
rect 12400 21428 12434 21440
rect 4430 21292 4436 21344
rect 4488 21332 4494 21344
rect 4890 21332 4896 21344
rect 4488 21304 4896 21332
rect 4488 21292 4494 21304
rect 4890 21292 4896 21304
rect 4948 21332 4954 21344
rect 5166 21332 5172 21344
rect 4948 21304 5172 21332
rect 4948 21292 4954 21304
rect 5166 21292 5172 21304
rect 5224 21292 5230 21344
rect 9398 21292 9404 21344
rect 9456 21292 9462 21344
rect 10410 21292 10416 21344
rect 10468 21292 10474 21344
rect 10502 21292 10508 21344
rect 10560 21292 10566 21344
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 12406 21332 12434 21428
rect 14384 21344 14412 21440
rect 11848 21304 12434 21332
rect 11848 21292 11854 21304
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 14366 21292 14372 21344
rect 14424 21332 14430 21344
rect 14461 21335 14519 21341
rect 14461 21332 14473 21335
rect 14424 21304 14473 21332
rect 14424 21292 14430 21304
rect 14461 21301 14473 21304
rect 14507 21301 14519 21335
rect 14461 21295 14519 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 15105 21335 15163 21341
rect 15105 21332 15117 21335
rect 15068 21304 15117 21332
rect 15068 21292 15074 21304
rect 15105 21301 15117 21304
rect 15151 21332 15163 21335
rect 15470 21332 15476 21344
rect 15151 21304 15476 21332
rect 15151 21301 15163 21304
rect 15105 21295 15163 21301
rect 15470 21292 15476 21304
rect 15528 21292 15534 21344
rect 15580 21341 15608 21508
rect 15565 21335 15623 21341
rect 15565 21301 15577 21335
rect 15611 21332 15623 21335
rect 15654 21332 15660 21344
rect 15611 21304 15660 21332
rect 15611 21301 15623 21304
rect 15565 21295 15623 21301
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16224 21332 16252 21632
rect 17236 21545 17264 21632
rect 22186 21604 22192 21616
rect 17512 21576 18552 21604
rect 17512 21548 17540 21576
rect 17221 21539 17279 21545
rect 17221 21505 17233 21539
rect 17267 21505 17279 21539
rect 17221 21499 17279 21505
rect 17494 21496 17500 21548
rect 17552 21496 17558 21548
rect 17770 21496 17776 21548
rect 17828 21496 17834 21548
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 17957 21539 18015 21545
rect 17957 21536 17969 21539
rect 17920 21508 17969 21536
rect 17920 21496 17926 21508
rect 17957 21505 17969 21508
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18046 21496 18052 21548
rect 18104 21536 18110 21548
rect 18524 21545 18552 21576
rect 20916 21576 22192 21604
rect 20916 21548 20944 21576
rect 22186 21564 22192 21576
rect 22244 21604 22250 21616
rect 23216 21604 23244 21632
rect 23676 21604 23704 21632
rect 22244 21576 23244 21604
rect 23308 21576 23704 21604
rect 22244 21564 22250 21576
rect 18233 21539 18291 21545
rect 18233 21536 18245 21539
rect 18104 21508 18245 21536
rect 18104 21496 18110 21508
rect 18233 21505 18245 21508
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 18509 21539 18567 21545
rect 18509 21505 18521 21539
rect 18555 21505 18567 21539
rect 18509 21499 18567 21505
rect 20438 21496 20444 21548
rect 20496 21496 20502 21548
rect 20530 21496 20536 21548
rect 20588 21496 20594 21548
rect 20714 21496 20720 21548
rect 20772 21496 20778 21548
rect 20898 21496 20904 21548
rect 20956 21496 20962 21548
rect 20990 21496 20996 21548
rect 21048 21536 21054 21548
rect 21910 21536 21916 21548
rect 21048 21508 21916 21536
rect 21048 21496 21054 21508
rect 21910 21496 21916 21508
rect 21968 21536 21974 21548
rect 23308 21545 23336 21576
rect 28350 21564 28356 21616
rect 28408 21564 28414 21616
rect 28828 21613 28856 21644
rect 30282 21632 30288 21684
rect 30340 21632 30346 21684
rect 31110 21632 31116 21684
rect 31168 21632 31174 21684
rect 31570 21632 31576 21684
rect 31628 21632 31634 21684
rect 33318 21632 33324 21684
rect 33376 21632 33382 21684
rect 28813 21607 28871 21613
rect 28813 21573 28825 21607
rect 28859 21573 28871 21607
rect 30469 21607 30527 21613
rect 30469 21604 30481 21607
rect 30038 21576 30481 21604
rect 28813 21567 28871 21573
rect 30469 21573 30481 21576
rect 30515 21573 30527 21607
rect 31588 21604 31616 21632
rect 30469 21567 30527 21573
rect 31128 21576 31616 21604
rect 22557 21539 22615 21545
rect 22557 21536 22569 21539
rect 21968 21508 22569 21536
rect 21968 21496 21974 21508
rect 22557 21505 22569 21508
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 23293 21539 23351 21545
rect 23293 21505 23305 21539
rect 23339 21505 23351 21539
rect 23293 21499 23351 21505
rect 23566 21496 23572 21548
rect 23624 21496 23630 21548
rect 24946 21496 24952 21548
rect 25004 21536 25010 21548
rect 25409 21539 25467 21545
rect 25409 21536 25421 21539
rect 25004 21508 25421 21536
rect 25004 21496 25010 21508
rect 25409 21505 25421 21508
rect 25455 21505 25467 21539
rect 25409 21499 25467 21505
rect 26418 21496 26424 21548
rect 26476 21496 26482 21548
rect 28368 21536 28396 21564
rect 28537 21539 28595 21545
rect 28537 21536 28549 21539
rect 28368 21508 28549 21536
rect 28537 21505 28549 21508
rect 28583 21505 28595 21539
rect 28537 21499 28595 21505
rect 30098 21496 30104 21548
rect 30156 21536 30162 21548
rect 30561 21539 30619 21545
rect 30561 21536 30573 21539
rect 30156 21508 30573 21536
rect 30156 21496 30162 21508
rect 30561 21505 30573 21508
rect 30607 21536 30619 21539
rect 30837 21539 30895 21545
rect 30837 21536 30849 21539
rect 30607 21508 30849 21536
rect 30607 21505 30619 21508
rect 30561 21499 30619 21505
rect 30837 21505 30849 21508
rect 30883 21505 30895 21539
rect 30837 21499 30895 21505
rect 31018 21496 31024 21548
rect 31076 21536 31082 21548
rect 31128 21545 31156 21576
rect 31113 21539 31171 21545
rect 31113 21536 31125 21539
rect 31076 21508 31125 21536
rect 31076 21496 31082 21508
rect 31113 21505 31125 21508
rect 31159 21505 31171 21539
rect 31113 21499 31171 21505
rect 31297 21539 31355 21545
rect 31297 21505 31309 21539
rect 31343 21536 31355 21539
rect 32030 21536 32036 21548
rect 31343 21508 32036 21536
rect 31343 21505 31355 21508
rect 31297 21499 31355 21505
rect 32030 21496 32036 21508
rect 32088 21496 32094 21548
rect 33229 21539 33287 21545
rect 33229 21536 33241 21539
rect 33152 21508 33241 21536
rect 17681 21471 17739 21477
rect 17681 21437 17693 21471
rect 17727 21437 17739 21471
rect 17681 21431 17739 21437
rect 17696 21400 17724 21431
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 22465 21471 22523 21477
rect 22465 21468 22477 21471
rect 21324 21440 22477 21468
rect 21324 21428 21330 21440
rect 22465 21437 22477 21440
rect 22511 21437 22523 21471
rect 22465 21431 22523 21437
rect 22925 21471 22983 21477
rect 22925 21437 22937 21471
rect 22971 21468 22983 21471
rect 23584 21468 23612 21496
rect 22971 21440 23612 21468
rect 22971 21437 22983 21440
rect 22925 21431 22983 21437
rect 24854 21428 24860 21480
rect 24912 21468 24918 21480
rect 25317 21471 25375 21477
rect 25317 21468 25329 21471
rect 24912 21440 25329 21468
rect 24912 21428 24918 21440
rect 25317 21437 25329 21440
rect 25363 21437 25375 21471
rect 26329 21471 26387 21477
rect 26329 21468 26341 21471
rect 25317 21431 25375 21437
rect 25792 21440 26341 21468
rect 17862 21400 17868 21412
rect 17696 21372 17868 21400
rect 17862 21360 17868 21372
rect 17920 21400 17926 21412
rect 18325 21403 18383 21409
rect 18325 21400 18337 21403
rect 17920 21372 18337 21400
rect 17920 21360 17926 21372
rect 18325 21369 18337 21372
rect 18371 21369 18383 21403
rect 18325 21363 18383 21369
rect 23569 21403 23627 21409
rect 23569 21369 23581 21403
rect 23615 21400 23627 21403
rect 23750 21400 23756 21412
rect 23615 21372 23756 21400
rect 23615 21369 23627 21372
rect 23569 21363 23627 21369
rect 23750 21360 23756 21372
rect 23808 21360 23814 21412
rect 25792 21409 25820 21440
rect 26329 21437 26341 21440
rect 26375 21437 26387 21471
rect 26329 21431 26387 21437
rect 25777 21403 25835 21409
rect 25777 21369 25789 21403
rect 25823 21369 25835 21403
rect 25777 21363 25835 21369
rect 33152 21344 33180 21508
rect 33229 21505 33241 21508
rect 33275 21505 33287 21539
rect 33229 21499 33287 21505
rect 18690 21332 18696 21344
rect 16224 21304 18696 21332
rect 18690 21292 18696 21304
rect 18748 21292 18754 21344
rect 32398 21292 32404 21344
rect 32456 21332 32462 21344
rect 32674 21332 32680 21344
rect 32456 21304 32680 21332
rect 32456 21292 32462 21304
rect 32674 21292 32680 21304
rect 32732 21292 32738 21344
rect 33134 21292 33140 21344
rect 33192 21292 33198 21344
rect 1104 21242 35248 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 35248 21242
rect 1104 21168 35248 21190
rect 3142 21088 3148 21140
rect 3200 21088 3206 21140
rect 3326 21088 3332 21140
rect 3384 21088 3390 21140
rect 4341 21131 4399 21137
rect 4341 21097 4353 21131
rect 4387 21128 4399 21131
rect 5074 21128 5080 21140
rect 4387 21100 5080 21128
rect 4387 21097 4399 21100
rect 4341 21091 4399 21097
rect 3160 20924 3188 21088
rect 3234 20924 3240 20936
rect 3160 20896 3240 20924
rect 3234 20884 3240 20896
rect 3292 20884 3298 20936
rect 4908 20856 4936 21100
rect 5074 21088 5080 21100
rect 5132 21088 5138 21140
rect 5166 21088 5172 21140
rect 5224 21128 5230 21140
rect 5629 21131 5687 21137
rect 5629 21128 5641 21131
rect 5224 21100 5641 21128
rect 5224 21088 5230 21100
rect 5629 21097 5641 21100
rect 5675 21128 5687 21131
rect 5810 21128 5816 21140
rect 5675 21100 5816 21128
rect 5675 21097 5687 21100
rect 5629 21091 5687 21097
rect 5810 21088 5816 21100
rect 5868 21088 5874 21140
rect 7374 21088 7380 21140
rect 7432 21088 7438 21140
rect 10137 21131 10195 21137
rect 10137 21097 10149 21131
rect 10183 21128 10195 21131
rect 10410 21128 10416 21140
rect 10183 21100 10416 21128
rect 10183 21097 10195 21100
rect 10137 21091 10195 21097
rect 10410 21088 10416 21100
rect 10468 21088 10474 21140
rect 10502 21088 10508 21140
rect 10560 21088 10566 21140
rect 15746 21088 15752 21140
rect 15804 21128 15810 21140
rect 17218 21128 17224 21140
rect 15804 21100 17224 21128
rect 15804 21088 15810 21100
rect 17218 21088 17224 21100
rect 17276 21088 17282 21140
rect 17313 21131 17371 21137
rect 17313 21097 17325 21131
rect 17359 21128 17371 21131
rect 17494 21128 17500 21140
rect 17359 21100 17500 21128
rect 17359 21097 17371 21100
rect 17313 21091 17371 21097
rect 17494 21088 17500 21100
rect 17552 21088 17558 21140
rect 17862 21088 17868 21140
rect 17920 21088 17926 21140
rect 23014 21088 23020 21140
rect 23072 21088 23078 21140
rect 26418 21088 26424 21140
rect 26476 21088 26482 21140
rect 5445 21063 5503 21069
rect 5445 21060 5457 21063
rect 5092 21032 5457 21060
rect 5092 21001 5120 21032
rect 5445 21029 5457 21032
rect 5491 21029 5503 21063
rect 5445 21023 5503 21029
rect 9585 21063 9643 21069
rect 9585 21029 9597 21063
rect 9631 21060 9643 21063
rect 9674 21060 9680 21072
rect 9631 21032 9680 21060
rect 9631 21029 9643 21032
rect 9585 21023 9643 21029
rect 9674 21020 9680 21032
rect 9732 21020 9738 21072
rect 5077 20995 5135 21001
rect 5077 20961 5089 20995
rect 5123 20961 5135 20995
rect 5077 20955 5135 20961
rect 5353 20995 5411 21001
rect 5353 20961 5365 20995
rect 5399 20992 5411 20995
rect 5994 20992 6000 21004
rect 5399 20964 6000 20992
rect 5399 20961 5411 20964
rect 5353 20955 5411 20961
rect 5994 20952 6000 20964
rect 6052 20952 6058 21004
rect 10520 20992 10548 21088
rect 10870 21020 10876 21072
rect 10928 21060 10934 21072
rect 11333 21063 11391 21069
rect 11333 21060 11345 21063
rect 10928 21032 11345 21060
rect 10928 21020 10934 21032
rect 11333 21029 11345 21032
rect 11379 21029 11391 21063
rect 11333 21023 11391 21029
rect 13357 21063 13415 21069
rect 13357 21029 13369 21063
rect 13403 21060 13415 21063
rect 13403 21032 17264 21060
rect 13403 21029 13415 21032
rect 13357 21023 13415 21029
rect 11977 20995 12035 21001
rect 10520 20964 11744 20992
rect 4982 20884 4988 20936
rect 5040 20884 5046 20936
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20924 7343 20927
rect 8386 20924 8392 20936
rect 7331 20896 8392 20924
rect 7331 20893 7343 20896
rect 7285 20887 7343 20893
rect 5813 20859 5871 20865
rect 5813 20856 5825 20859
rect 4908 20828 5825 20856
rect 5813 20825 5825 20828
rect 5859 20856 5871 20859
rect 6086 20856 6092 20868
rect 5859 20828 6092 20856
rect 5859 20825 5871 20828
rect 5813 20819 5871 20825
rect 6086 20816 6092 20828
rect 6144 20816 6150 20868
rect 7576 20800 7604 20896
rect 8386 20884 8392 20896
rect 8444 20884 8450 20936
rect 9861 20927 9919 20933
rect 9861 20924 9873 20927
rect 9416 20896 9873 20924
rect 9416 20868 9444 20896
rect 9861 20893 9873 20896
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 10686 20884 10692 20936
rect 10744 20884 10750 20936
rect 10778 20884 10784 20936
rect 10836 20884 10842 20936
rect 10962 20884 10968 20936
rect 11020 20884 11026 20936
rect 11146 20884 11152 20936
rect 11204 20884 11210 20936
rect 11238 20884 11244 20936
rect 11296 20884 11302 20936
rect 11716 20933 11744 20964
rect 11977 20961 11989 20995
rect 12023 20992 12035 20995
rect 12713 20995 12771 21001
rect 12713 20992 12725 20995
rect 12023 20964 12725 20992
rect 12023 20961 12035 20964
rect 11977 20955 12035 20961
rect 12713 20961 12725 20964
rect 12759 20961 12771 20995
rect 12713 20955 12771 20961
rect 13906 20952 13912 21004
rect 13964 20992 13970 21004
rect 15013 20995 15071 21001
rect 13964 20964 14688 20992
rect 13964 20952 13970 20964
rect 11701 20927 11759 20933
rect 11701 20893 11713 20927
rect 11747 20893 11759 20927
rect 11701 20887 11759 20893
rect 11790 20884 11796 20936
rect 11848 20924 11854 20936
rect 12069 20927 12127 20933
rect 12069 20924 12081 20927
rect 11848 20896 12081 20924
rect 11848 20884 11854 20896
rect 12069 20893 12081 20896
rect 12115 20893 12127 20927
rect 12069 20887 12127 20893
rect 12253 20927 12311 20933
rect 12253 20893 12265 20927
rect 12299 20893 12311 20927
rect 12253 20887 12311 20893
rect 12989 20927 13047 20933
rect 12989 20893 13001 20927
rect 13035 20924 13047 20927
rect 14274 20924 14280 20936
rect 13035 20896 14280 20924
rect 13035 20893 13047 20896
rect 12989 20887 13047 20893
rect 8297 20859 8355 20865
rect 8297 20825 8309 20859
rect 8343 20856 8355 20859
rect 9398 20856 9404 20868
rect 8343 20828 9404 20856
rect 8343 20825 8355 20828
rect 8297 20819 8355 20825
rect 9398 20816 9404 20828
rect 9456 20816 9462 20868
rect 9493 20859 9551 20865
rect 9493 20825 9505 20859
rect 9539 20856 9551 20859
rect 9953 20859 10011 20865
rect 9953 20856 9965 20859
rect 9539 20828 9965 20856
rect 9539 20825 9551 20828
rect 9493 20819 9551 20825
rect 9953 20825 9965 20828
rect 9999 20825 10011 20859
rect 9953 20819 10011 20825
rect 10505 20859 10563 20865
rect 10505 20825 10517 20859
rect 10551 20856 10563 20859
rect 10980 20856 11008 20884
rect 10551 20828 11008 20856
rect 11057 20859 11115 20865
rect 10551 20825 10563 20828
rect 10505 20819 10563 20825
rect 11057 20825 11069 20859
rect 11103 20856 11115 20859
rect 11422 20856 11428 20868
rect 11103 20828 11428 20856
rect 11103 20825 11115 20828
rect 11057 20819 11115 20825
rect 4798 20748 4804 20800
rect 4856 20788 4862 20800
rect 5603 20791 5661 20797
rect 5603 20788 5615 20791
rect 4856 20760 5615 20788
rect 4856 20748 4862 20760
rect 5603 20757 5615 20760
rect 5649 20757 5661 20791
rect 5603 20751 5661 20757
rect 7558 20748 7564 20800
rect 7616 20788 7622 20800
rect 7745 20791 7803 20797
rect 7745 20788 7757 20791
rect 7616 20760 7757 20788
rect 7616 20748 7622 20760
rect 7745 20757 7757 20760
rect 7791 20757 7803 20791
rect 7745 20751 7803 20757
rect 8757 20791 8815 20797
rect 8757 20757 8769 20791
rect 8803 20788 8815 20791
rect 9582 20788 9588 20800
rect 8803 20760 9588 20788
rect 8803 20757 8815 20760
rect 8757 20751 8815 20757
rect 9582 20748 9588 20760
rect 9640 20788 9646 20800
rect 9769 20791 9827 20797
rect 9769 20788 9781 20791
rect 9640 20760 9781 20788
rect 9640 20748 9646 20760
rect 9769 20757 9781 20760
rect 9815 20757 9827 20791
rect 9968 20788 9996 20819
rect 11422 20816 11428 20828
rect 11480 20816 11486 20868
rect 11609 20859 11667 20865
rect 11609 20825 11621 20859
rect 11655 20856 11667 20859
rect 12161 20859 12219 20865
rect 12161 20856 12173 20859
rect 11655 20828 12173 20856
rect 11655 20825 11667 20828
rect 11609 20819 11667 20825
rect 12161 20825 12173 20828
rect 12207 20825 12219 20859
rect 12268 20856 12296 20887
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 14366 20884 14372 20936
rect 14424 20884 14430 20936
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 14660 20933 14688 20964
rect 15013 20961 15025 20995
rect 15059 20992 15071 20995
rect 15565 20995 15623 21001
rect 15565 20992 15577 20995
rect 15059 20964 15577 20992
rect 15059 20961 15071 20964
rect 15013 20955 15071 20961
rect 15565 20961 15577 20964
rect 15611 20961 15623 20995
rect 15565 20955 15623 20961
rect 17236 20992 17264 21032
rect 17236 20964 17908 20992
rect 14645 20927 14703 20933
rect 14645 20893 14657 20927
rect 14691 20893 14703 20927
rect 14645 20887 14703 20893
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 14921 20927 14979 20933
rect 14921 20893 14933 20927
rect 14967 20893 14979 20927
rect 14921 20887 14979 20893
rect 14461 20859 14519 20865
rect 14461 20856 14473 20859
rect 12268 20828 14473 20856
rect 12161 20819 12219 20825
rect 10870 20788 10876 20800
rect 9968 20760 10876 20788
rect 9769 20751 9827 20757
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 10962 20748 10968 20800
rect 11020 20788 11026 20800
rect 11517 20791 11575 20797
rect 11517 20788 11529 20791
rect 11020 20760 11529 20788
rect 11020 20748 11026 20760
rect 11517 20757 11529 20760
rect 11563 20757 11575 20791
rect 11517 20751 11575 20757
rect 11698 20748 11704 20800
rect 11756 20788 11762 20800
rect 12406 20788 12434 20828
rect 14461 20825 14473 20828
rect 14507 20856 14519 20859
rect 14844 20856 14872 20887
rect 14507 20828 14872 20856
rect 14936 20856 14964 20887
rect 15194 20884 15200 20936
rect 15252 20884 15258 20936
rect 15470 20884 15476 20936
rect 15528 20884 15534 20936
rect 15654 20884 15660 20936
rect 15712 20884 15718 20936
rect 17236 20933 17264 20964
rect 17221 20927 17279 20933
rect 17221 20893 17233 20927
rect 17267 20893 17279 20927
rect 17221 20887 17279 20893
rect 17310 20884 17316 20936
rect 17368 20924 17374 20936
rect 17880 20933 17908 20964
rect 20346 20952 20352 21004
rect 20404 20952 20410 21004
rect 25130 20952 25136 21004
rect 25188 20952 25194 21004
rect 25516 20964 26280 20992
rect 25516 20936 25544 20964
rect 17405 20927 17463 20933
rect 17405 20924 17417 20927
rect 17368 20896 17417 20924
rect 17368 20884 17374 20896
rect 17405 20893 17417 20896
rect 17451 20924 17463 20927
rect 17681 20927 17739 20933
rect 17681 20924 17693 20927
rect 17451 20896 17693 20924
rect 17451 20893 17463 20896
rect 17405 20887 17463 20893
rect 17681 20893 17693 20896
rect 17727 20893 17739 20927
rect 17681 20887 17739 20893
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20924 17923 20927
rect 17954 20924 17960 20936
rect 17911 20896 17960 20924
rect 17911 20893 17923 20896
rect 17865 20887 17923 20893
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 20714 20884 20720 20936
rect 20772 20884 20778 20936
rect 21177 20927 21235 20933
rect 21177 20893 21189 20927
rect 21223 20924 21235 20927
rect 21361 20927 21419 20933
rect 21361 20924 21373 20927
rect 21223 20896 21373 20924
rect 21223 20893 21235 20896
rect 21177 20887 21235 20893
rect 21361 20893 21373 20896
rect 21407 20893 21419 20927
rect 21361 20887 21419 20893
rect 21726 20884 21732 20936
rect 21784 20884 21790 20936
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 24949 20927 25007 20933
rect 24949 20924 24961 20927
rect 24912 20896 24961 20924
rect 24912 20884 24918 20896
rect 24949 20893 24961 20896
rect 24995 20893 25007 20927
rect 24949 20887 25007 20893
rect 25038 20884 25044 20936
rect 25096 20884 25102 20936
rect 25498 20884 25504 20936
rect 25556 20884 25562 20936
rect 25593 20927 25651 20933
rect 25593 20893 25605 20927
rect 25639 20893 25651 20927
rect 25593 20887 25651 20893
rect 15562 20856 15568 20868
rect 14936 20828 15568 20856
rect 14507 20825 14519 20828
rect 14461 20819 14519 20825
rect 15562 20816 15568 20828
rect 15620 20816 15626 20868
rect 15672 20856 15700 20884
rect 16298 20856 16304 20868
rect 15672 20828 16304 20856
rect 16298 20816 16304 20828
rect 16356 20816 16362 20868
rect 25056 20856 25084 20884
rect 25608 20856 25636 20887
rect 25774 20884 25780 20936
rect 25832 20884 25838 20936
rect 25866 20884 25872 20936
rect 25924 20924 25930 20936
rect 26252 20933 26280 20964
rect 25961 20927 26019 20933
rect 25961 20924 25973 20927
rect 25924 20896 25973 20924
rect 25924 20884 25930 20896
rect 25961 20893 25973 20896
rect 26007 20893 26019 20927
rect 25961 20887 26019 20893
rect 26237 20927 26295 20933
rect 26237 20893 26249 20927
rect 26283 20893 26295 20927
rect 26237 20887 26295 20893
rect 33318 20884 33324 20936
rect 33376 20884 33382 20936
rect 26326 20856 26332 20868
rect 25056 20828 26332 20856
rect 26326 20816 26332 20828
rect 26384 20816 26390 20868
rect 34330 20816 34336 20868
rect 34388 20816 34394 20868
rect 11756 20760 12434 20788
rect 11756 20748 11762 20760
rect 12894 20748 12900 20800
rect 12952 20748 12958 20800
rect 13909 20791 13967 20797
rect 13909 20757 13921 20791
rect 13955 20788 13967 20791
rect 14366 20788 14372 20800
rect 13955 20760 14372 20788
rect 13955 20757 13967 20760
rect 13909 20751 13967 20757
rect 14366 20748 14372 20760
rect 14424 20748 14430 20800
rect 15378 20748 15384 20800
rect 15436 20748 15442 20800
rect 15470 20748 15476 20800
rect 15528 20788 15534 20800
rect 15746 20788 15752 20800
rect 15528 20760 15752 20788
rect 15528 20748 15534 20760
rect 15746 20748 15752 20760
rect 15804 20788 15810 20800
rect 15933 20791 15991 20797
rect 15933 20788 15945 20791
rect 15804 20760 15945 20788
rect 15804 20748 15810 20760
rect 15933 20757 15945 20760
rect 15979 20788 15991 20791
rect 16114 20788 16120 20800
rect 15979 20760 16120 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 1104 20698 35236 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 35236 20698
rect 1104 20624 35236 20646
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 10870 20544 10876 20596
rect 10928 20584 10934 20596
rect 11054 20584 11060 20596
rect 10928 20556 11060 20584
rect 10928 20544 10934 20556
rect 11054 20544 11060 20556
rect 11112 20544 11118 20596
rect 11146 20544 11152 20596
rect 11204 20584 11210 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 11204 20556 11621 20584
rect 11204 20544 11210 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 11609 20547 11667 20553
rect 12805 20587 12863 20593
rect 12805 20553 12817 20587
rect 12851 20584 12863 20587
rect 12894 20584 12900 20596
rect 12851 20556 12900 20584
rect 12851 20553 12863 20556
rect 12805 20547 12863 20553
rect 12894 20544 12900 20556
rect 12952 20544 12958 20596
rect 13262 20544 13268 20596
rect 13320 20584 13326 20596
rect 13320 20556 13952 20584
rect 13320 20544 13326 20556
rect 5994 20476 6000 20528
rect 6052 20516 6058 20528
rect 6641 20519 6699 20525
rect 6641 20516 6653 20519
rect 6052 20488 6653 20516
rect 6052 20476 6058 20488
rect 6641 20485 6653 20488
rect 6687 20485 6699 20519
rect 6641 20479 6699 20485
rect 7374 20476 7380 20528
rect 7432 20476 7438 20528
rect 11072 20516 11100 20544
rect 12069 20519 12127 20525
rect 12069 20516 12081 20519
rect 11072 20488 12081 20516
rect 12069 20485 12081 20488
rect 12115 20516 12127 20519
rect 12526 20516 12532 20528
rect 12115 20488 12532 20516
rect 12115 20485 12127 20488
rect 12069 20479 12127 20485
rect 12526 20476 12532 20488
rect 12584 20476 12590 20528
rect 12820 20488 13676 20516
rect 6362 20408 6368 20460
rect 6420 20408 6426 20460
rect 8297 20451 8355 20457
rect 8297 20417 8309 20451
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 9953 20451 10011 20457
rect 9953 20417 9965 20451
rect 9999 20448 10011 20451
rect 10410 20448 10416 20460
rect 9999 20420 10416 20448
rect 9999 20417 10011 20420
rect 9953 20411 10011 20417
rect 8113 20383 8171 20389
rect 8113 20349 8125 20383
rect 8159 20380 8171 20383
rect 8312 20380 8340 20411
rect 10410 20408 10416 20420
rect 10468 20408 10474 20460
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20448 11575 20451
rect 11606 20448 11612 20460
rect 11563 20420 11612 20448
rect 11563 20417 11575 20420
rect 11517 20411 11575 20417
rect 11606 20408 11612 20420
rect 11664 20408 11670 20460
rect 11698 20408 11704 20460
rect 11756 20408 11762 20460
rect 12820 20457 12848 20488
rect 12621 20451 12679 20457
rect 12621 20417 12633 20451
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 12805 20451 12863 20457
rect 12805 20417 12817 20451
rect 12851 20417 12863 20451
rect 12805 20411 12863 20417
rect 8159 20352 8340 20380
rect 9125 20383 9183 20389
rect 8159 20349 8171 20352
rect 8113 20343 8171 20349
rect 9125 20349 9137 20383
rect 9171 20380 9183 20383
rect 9171 20352 9628 20380
rect 9171 20349 9183 20352
rect 9125 20343 9183 20349
rect 9600 20324 9628 20352
rect 10042 20340 10048 20392
rect 10100 20340 10106 20392
rect 10321 20383 10379 20389
rect 10321 20349 10333 20383
rect 10367 20380 10379 20383
rect 10686 20380 10692 20392
rect 10367 20352 10692 20380
rect 10367 20349 10379 20352
rect 10321 20343 10379 20349
rect 10686 20340 10692 20352
rect 10744 20340 10750 20392
rect 9582 20272 9588 20324
rect 9640 20312 9646 20324
rect 12437 20315 12495 20321
rect 12437 20312 12449 20315
rect 9640 20284 12449 20312
rect 9640 20272 9646 20284
rect 12437 20281 12449 20284
rect 12483 20312 12495 20315
rect 12526 20312 12532 20324
rect 12483 20284 12532 20312
rect 12483 20281 12495 20284
rect 12437 20275 12495 20281
rect 12526 20272 12532 20284
rect 12584 20272 12590 20324
rect 12636 20244 12664 20411
rect 12820 20312 12848 20411
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 13076 20451 13134 20457
rect 13076 20448 13088 20451
rect 12952 20420 13088 20448
rect 12952 20408 12958 20420
rect 13076 20417 13088 20420
rect 13122 20417 13134 20451
rect 13076 20411 13134 20417
rect 13096 20380 13124 20411
rect 13170 20408 13176 20460
rect 13228 20408 13234 20460
rect 13262 20408 13268 20460
rect 13320 20408 13326 20460
rect 13354 20408 13360 20460
rect 13412 20457 13418 20460
rect 13412 20451 13451 20457
rect 13439 20417 13451 20451
rect 13412 20411 13451 20417
rect 13412 20408 13418 20411
rect 13538 20408 13544 20460
rect 13596 20408 13602 20460
rect 13648 20457 13676 20488
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20417 13691 20451
rect 13633 20411 13691 20417
rect 13722 20408 13728 20460
rect 13780 20448 13786 20460
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13780 20420 13829 20448
rect 13780 20408 13786 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 13924 20448 13952 20556
rect 14274 20544 14280 20596
rect 14332 20544 14338 20596
rect 15013 20587 15071 20593
rect 15013 20553 15025 20587
rect 15059 20584 15071 20587
rect 15194 20584 15200 20596
rect 15059 20556 15200 20584
rect 15059 20553 15071 20556
rect 15013 20547 15071 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15562 20544 15568 20596
rect 15620 20544 15626 20596
rect 17589 20587 17647 20593
rect 15672 20556 17080 20584
rect 14001 20451 14059 20457
rect 14001 20448 14013 20451
rect 13924 20420 14013 20448
rect 13817 20411 13875 20417
rect 14001 20417 14013 20420
rect 14047 20417 14059 20451
rect 14001 20411 14059 20417
rect 14090 20408 14096 20460
rect 14148 20408 14154 20460
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 14550 20448 14556 20460
rect 14332 20420 14556 20448
rect 14332 20408 14338 20420
rect 14550 20408 14556 20420
rect 14608 20448 14614 20460
rect 15197 20451 15255 20457
rect 15197 20448 15209 20451
rect 14608 20420 15209 20448
rect 14608 20408 14614 20420
rect 15197 20417 15209 20420
rect 15243 20448 15255 20451
rect 15672 20448 15700 20556
rect 17052 20528 17080 20556
rect 17589 20553 17601 20587
rect 17635 20584 17647 20587
rect 17678 20584 17684 20596
rect 17635 20556 17684 20584
rect 17635 20553 17647 20556
rect 17589 20547 17647 20553
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 20438 20544 20444 20596
rect 20496 20544 20502 20596
rect 20898 20544 20904 20596
rect 20956 20544 20962 20596
rect 22281 20587 22339 20593
rect 22281 20553 22293 20587
rect 22327 20584 22339 20587
rect 22646 20584 22652 20596
rect 22327 20556 22652 20584
rect 22327 20553 22339 20556
rect 22281 20547 22339 20553
rect 17034 20476 17040 20528
rect 17092 20516 17098 20528
rect 17092 20488 17448 20516
rect 17092 20476 17098 20488
rect 15243 20420 15700 20448
rect 15243 20417 15255 20420
rect 15197 20411 15255 20417
rect 15746 20408 15752 20460
rect 15804 20408 15810 20460
rect 15856 20420 17172 20448
rect 13096 20352 13676 20380
rect 13648 20324 13676 20352
rect 12897 20315 12955 20321
rect 12897 20312 12909 20315
rect 12820 20284 12909 20312
rect 12897 20281 12909 20284
rect 12943 20281 12955 20315
rect 12897 20275 12955 20281
rect 13630 20272 13636 20324
rect 13688 20272 13694 20324
rect 13740 20244 13768 20408
rect 15470 20340 15476 20392
rect 15528 20380 15534 20392
rect 15856 20380 15884 20420
rect 15528 20352 15884 20380
rect 16025 20383 16083 20389
rect 15528 20340 15534 20352
rect 16025 20349 16037 20383
rect 16071 20380 16083 20383
rect 16298 20380 16304 20392
rect 16071 20352 16304 20380
rect 16071 20349 16083 20352
rect 16025 20343 16083 20349
rect 13814 20272 13820 20324
rect 13872 20312 13878 20324
rect 13909 20315 13967 20321
rect 13909 20312 13921 20315
rect 13872 20284 13921 20312
rect 13872 20272 13878 20284
rect 13909 20281 13921 20284
rect 13955 20281 13967 20315
rect 13909 20275 13967 20281
rect 14921 20315 14979 20321
rect 14921 20281 14933 20315
rect 14967 20312 14979 20315
rect 16040 20312 16068 20343
rect 16298 20340 16304 20352
rect 16356 20340 16362 20392
rect 14967 20284 16068 20312
rect 14967 20281 14979 20284
rect 14921 20275 14979 20281
rect 12636 20216 13768 20244
rect 15381 20247 15439 20253
rect 15381 20213 15393 20247
rect 15427 20244 15439 20247
rect 15838 20244 15844 20256
rect 15427 20216 15844 20244
rect 15427 20213 15439 20216
rect 15381 20207 15439 20213
rect 15838 20204 15844 20216
rect 15896 20244 15902 20256
rect 15933 20247 15991 20253
rect 15933 20244 15945 20247
rect 15896 20216 15945 20244
rect 15896 20204 15902 20216
rect 15933 20213 15945 20216
rect 15979 20213 15991 20247
rect 15933 20207 15991 20213
rect 16393 20247 16451 20253
rect 16393 20213 16405 20247
rect 16439 20244 16451 20247
rect 17034 20244 17040 20256
rect 16439 20216 17040 20244
rect 16439 20213 16451 20216
rect 16393 20207 16451 20213
rect 17034 20204 17040 20216
rect 17092 20204 17098 20256
rect 17144 20244 17172 20420
rect 17218 20408 17224 20460
rect 17276 20408 17282 20460
rect 17420 20457 17448 20488
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17696 20448 17724 20544
rect 20456 20516 20484 20544
rect 21361 20519 21419 20525
rect 20456 20488 20668 20516
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17696 20420 18061 20448
rect 17405 20411 17463 20417
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18969 20451 19027 20457
rect 18969 20448 18981 20451
rect 18049 20411 18107 20417
rect 18248 20420 18981 20448
rect 17954 20340 17960 20392
rect 18012 20340 18018 20392
rect 17310 20272 17316 20324
rect 17368 20312 17374 20324
rect 18248 20312 18276 20420
rect 18969 20417 18981 20420
rect 19015 20417 19027 20451
rect 18969 20411 19027 20417
rect 20346 20408 20352 20460
rect 20404 20448 20410 20460
rect 20441 20451 20499 20457
rect 20441 20448 20453 20451
rect 20404 20420 20453 20448
rect 20404 20408 20410 20420
rect 20441 20417 20453 20420
rect 20487 20417 20499 20451
rect 20441 20411 20499 20417
rect 20530 20408 20536 20460
rect 20588 20408 20594 20460
rect 20640 20457 20668 20488
rect 21361 20485 21373 20519
rect 21407 20516 21419 20519
rect 21726 20516 21732 20528
rect 21407 20488 21732 20516
rect 21407 20485 21419 20488
rect 21361 20479 21419 20485
rect 21726 20476 21732 20488
rect 21784 20476 21790 20528
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20448 20683 20451
rect 20993 20451 21051 20457
rect 20993 20448 21005 20451
rect 20671 20420 21005 20448
rect 20671 20417 20683 20420
rect 20625 20411 20683 20417
rect 20993 20417 21005 20420
rect 21039 20417 21051 20451
rect 21177 20451 21235 20457
rect 21177 20448 21189 20451
rect 20993 20411 21051 20417
rect 21100 20420 21189 20448
rect 18877 20383 18935 20389
rect 18877 20380 18889 20383
rect 18432 20352 18889 20380
rect 18432 20321 18460 20352
rect 18877 20349 18889 20352
rect 18923 20349 18935 20383
rect 18877 20343 18935 20349
rect 19797 20383 19855 20389
rect 19797 20349 19809 20383
rect 19843 20349 19855 20383
rect 19797 20343 19855 20349
rect 17368 20284 18276 20312
rect 18417 20315 18475 20321
rect 17368 20272 17374 20284
rect 18417 20281 18429 20315
rect 18463 20281 18475 20315
rect 19812 20312 19840 20343
rect 20346 20312 20352 20324
rect 19812 20284 20352 20312
rect 18417 20275 18475 20281
rect 20346 20272 20352 20284
rect 20404 20272 20410 20324
rect 20548 20312 20576 20408
rect 20717 20383 20775 20389
rect 20717 20349 20729 20383
rect 20763 20380 20775 20383
rect 20806 20380 20812 20392
rect 20763 20352 20812 20380
rect 20763 20349 20775 20352
rect 20717 20343 20775 20349
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 20622 20312 20628 20324
rect 20548 20284 20628 20312
rect 20622 20272 20628 20284
rect 20680 20312 20686 20324
rect 21100 20312 21128 20420
rect 21177 20417 21189 20420
rect 21223 20417 21235 20451
rect 21177 20411 21235 20417
rect 21266 20408 21272 20460
rect 21324 20448 21330 20460
rect 22296 20448 22324 20547
rect 22646 20544 22652 20556
rect 22704 20544 22710 20596
rect 24578 20544 24584 20596
rect 24636 20544 24642 20596
rect 24946 20544 24952 20596
rect 25004 20544 25010 20596
rect 33318 20544 33324 20596
rect 33376 20584 33382 20596
rect 33965 20587 34023 20593
rect 33965 20584 33977 20587
rect 33376 20556 33977 20584
rect 33376 20544 33382 20556
rect 33965 20553 33977 20556
rect 34011 20553 34023 20587
rect 33965 20547 34023 20553
rect 24857 20519 24915 20525
rect 24857 20516 24869 20519
rect 21324 20420 22324 20448
rect 22480 20488 23152 20516
rect 21324 20408 21330 20420
rect 22480 20312 22508 20488
rect 23124 20457 23152 20488
rect 24688 20488 24869 20516
rect 24688 20460 24716 20488
rect 24857 20485 24869 20488
rect 24903 20485 24915 20519
rect 24964 20516 24992 20544
rect 24964 20488 25268 20516
rect 24857 20479 24915 20485
rect 22925 20451 22983 20457
rect 22925 20448 22937 20451
rect 20680 20284 21128 20312
rect 22066 20284 22508 20312
rect 20680 20272 20686 20284
rect 17770 20244 17776 20256
rect 17144 20216 17776 20244
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 22066 20244 22094 20284
rect 22480 20256 22508 20284
rect 22572 20420 22937 20448
rect 22572 20256 22600 20420
rect 22925 20417 22937 20420
rect 22971 20417 22983 20451
rect 22925 20411 22983 20417
rect 23109 20451 23167 20457
rect 23109 20417 23121 20451
rect 23155 20448 23167 20451
rect 23385 20451 23443 20457
rect 23385 20448 23397 20451
rect 23155 20420 23397 20448
rect 23155 20417 23167 20420
rect 23109 20411 23167 20417
rect 23385 20417 23397 20420
rect 23431 20417 23443 20451
rect 23385 20411 23443 20417
rect 24670 20408 24676 20460
rect 24728 20408 24734 20460
rect 24765 20451 24823 20457
rect 24765 20417 24777 20451
rect 24811 20417 24823 20451
rect 24765 20411 24823 20417
rect 24949 20451 25007 20457
rect 24949 20417 24961 20451
rect 24995 20417 25007 20451
rect 24949 20411 25007 20417
rect 24780 20380 24808 20411
rect 24964 20380 24992 20411
rect 25130 20408 25136 20460
rect 25188 20408 25194 20460
rect 25240 20457 25268 20488
rect 33226 20476 33232 20528
rect 33284 20476 33290 20528
rect 25225 20451 25283 20457
rect 25225 20417 25237 20451
rect 25271 20417 25283 20451
rect 25774 20448 25780 20460
rect 25225 20411 25283 20417
rect 25332 20420 25780 20448
rect 25332 20380 25360 20420
rect 25774 20408 25780 20420
rect 25832 20408 25838 20460
rect 26237 20451 26295 20457
rect 26237 20417 26249 20451
rect 26283 20448 26295 20451
rect 26326 20448 26332 20460
rect 26283 20420 26332 20448
rect 26283 20417 26295 20420
rect 26237 20411 26295 20417
rect 26326 20408 26332 20420
rect 26384 20408 26390 20460
rect 26145 20383 26203 20389
rect 26145 20380 26157 20383
rect 24780 20352 24900 20380
rect 24872 20324 24900 20352
rect 24964 20352 25360 20380
rect 25608 20352 26157 20380
rect 24854 20272 24860 20324
rect 24912 20272 24918 20324
rect 19576 20216 22094 20244
rect 19576 20204 19582 20216
rect 22462 20204 22468 20256
rect 22520 20204 22526 20256
rect 22554 20204 22560 20256
rect 22612 20204 22618 20256
rect 23014 20204 23020 20256
rect 23072 20204 23078 20256
rect 23750 20204 23756 20256
rect 23808 20244 23814 20256
rect 24964 20244 24992 20352
rect 25608 20324 25636 20352
rect 26145 20349 26157 20352
rect 26191 20349 26203 20383
rect 26145 20343 26203 20349
rect 32217 20383 32275 20389
rect 32217 20349 32229 20383
rect 32263 20349 32275 20383
rect 32217 20343 32275 20349
rect 25590 20272 25596 20324
rect 25648 20272 25654 20324
rect 23808 20216 24992 20244
rect 23808 20204 23814 20216
rect 26510 20204 26516 20256
rect 26568 20204 26574 20256
rect 31941 20247 31999 20253
rect 31941 20213 31953 20247
rect 31987 20244 31999 20247
rect 32232 20244 32260 20343
rect 32490 20340 32496 20392
rect 32548 20340 32554 20392
rect 32674 20244 32680 20256
rect 31987 20216 32680 20244
rect 31987 20213 31999 20216
rect 31941 20207 31999 20213
rect 32674 20204 32680 20216
rect 32732 20204 32738 20256
rect 1104 20154 35248 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 35248 20154
rect 1104 20080 35248 20102
rect 7374 20000 7380 20052
rect 7432 20000 7438 20052
rect 8294 20000 8300 20052
rect 8352 20000 8358 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 13173 20043 13231 20049
rect 13173 20009 13185 20043
rect 13219 20040 13231 20043
rect 13722 20040 13728 20052
rect 13219 20012 13728 20040
rect 13219 20009 13231 20012
rect 13173 20003 13231 20009
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14090 20000 14096 20052
rect 14148 20000 14154 20052
rect 14274 20000 14280 20052
rect 14332 20000 14338 20052
rect 14366 20000 14372 20052
rect 14424 20040 14430 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14424 20012 14933 20040
rect 14424 20000 14430 20012
rect 14921 20009 14933 20012
rect 14967 20040 14979 20043
rect 15470 20040 15476 20052
rect 14967 20012 15476 20040
rect 14967 20009 14979 20012
rect 14921 20003 14979 20009
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 16298 20000 16304 20052
rect 16356 20040 16362 20052
rect 16945 20043 17003 20049
rect 16945 20040 16957 20043
rect 16356 20012 16957 20040
rect 16356 20000 16362 20012
rect 16945 20009 16957 20012
rect 16991 20009 17003 20043
rect 16945 20003 17003 20009
rect 17129 20043 17187 20049
rect 17129 20009 17141 20043
rect 17175 20040 17187 20043
rect 17586 20040 17592 20052
rect 17175 20012 17592 20040
rect 17175 20009 17187 20012
rect 17129 20003 17187 20009
rect 10778 19932 10784 19984
rect 10836 19972 10842 19984
rect 12066 19972 12072 19984
rect 10836 19944 12072 19972
rect 10836 19932 10842 19944
rect 12066 19932 12072 19944
rect 12124 19972 12130 19984
rect 13262 19972 13268 19984
rect 12124 19944 13268 19972
rect 12124 19932 12130 19944
rect 13262 19932 13268 19944
rect 13320 19932 13326 19984
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 14108 19904 14136 20000
rect 16960 19972 16988 20003
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 20438 20000 20444 20052
rect 20496 20040 20502 20052
rect 20809 20043 20867 20049
rect 20809 20040 20821 20043
rect 20496 20012 20821 20040
rect 20496 20000 20502 20012
rect 20809 20009 20821 20012
rect 20855 20009 20867 20043
rect 20809 20003 20867 20009
rect 21542 20000 21548 20052
rect 21600 20040 21606 20052
rect 21637 20043 21695 20049
rect 21637 20040 21649 20043
rect 21600 20012 21649 20040
rect 21600 20000 21606 20012
rect 21637 20009 21649 20012
rect 21683 20040 21695 20043
rect 21683 20012 22094 20040
rect 21683 20009 21695 20012
rect 21637 20003 21695 20009
rect 18506 19972 18512 19984
rect 16960 19944 18512 19972
rect 18506 19932 18512 19944
rect 18564 19972 18570 19984
rect 18564 19944 20576 19972
rect 18564 19932 18570 19944
rect 11112 19876 11928 19904
rect 11112 19864 11118 19876
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 7285 19839 7343 19845
rect 7285 19805 7297 19839
rect 7331 19836 7343 19839
rect 7331 19808 7604 19836
rect 7331 19805 7343 19808
rect 7285 19799 7343 19805
rect 7576 19712 7604 19808
rect 11790 19796 11796 19848
rect 11848 19796 11854 19848
rect 11900 19845 11928 19876
rect 13372 19876 14136 19904
rect 17497 19907 17555 19913
rect 11885 19839 11943 19845
rect 11885 19805 11897 19839
rect 11931 19805 11943 19839
rect 11885 19799 11943 19805
rect 11974 19796 11980 19848
rect 12032 19836 12038 19848
rect 13372 19845 13400 19876
rect 17497 19873 17509 19907
rect 17543 19904 17555 19907
rect 17770 19904 17776 19916
rect 17543 19876 17776 19904
rect 17543 19873 17555 19876
rect 17497 19867 17555 19873
rect 17770 19864 17776 19876
rect 17828 19904 17834 19916
rect 19518 19904 19524 19916
rect 17828 19876 19524 19904
rect 17828 19864 17834 19876
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 20548 19904 20576 19944
rect 20622 19932 20628 19984
rect 20680 19972 20686 19984
rect 20901 19975 20959 19981
rect 20901 19972 20913 19975
rect 20680 19944 20913 19972
rect 20680 19932 20686 19944
rect 20901 19941 20913 19944
rect 20947 19941 20959 19975
rect 22066 19972 22094 20012
rect 23014 20000 23020 20052
rect 23072 20000 23078 20052
rect 24949 20043 25007 20049
rect 24949 20009 24961 20043
rect 24995 20040 25007 20043
rect 25130 20040 25136 20052
rect 24995 20012 25136 20040
rect 24995 20009 25007 20012
rect 24949 20003 25007 20009
rect 25130 20000 25136 20012
rect 25188 20000 25194 20052
rect 25866 20000 25872 20052
rect 25924 20000 25930 20052
rect 26053 20043 26111 20049
rect 26053 20009 26065 20043
rect 26099 20009 26111 20043
rect 26053 20003 26111 20009
rect 22554 19972 22560 19984
rect 22066 19944 22560 19972
rect 20901 19935 20959 19941
rect 22554 19932 22560 19944
rect 22612 19972 22618 19984
rect 23032 19972 23060 20000
rect 26068 19972 26096 20003
rect 26510 20000 26516 20052
rect 26568 20040 26574 20052
rect 26568 20012 27292 20040
rect 26568 20000 26574 20012
rect 27154 19972 27160 19984
rect 22612 19944 22876 19972
rect 23032 19944 23428 19972
rect 26068 19944 27160 19972
rect 22612 19932 22618 19944
rect 22186 19904 22192 19916
rect 20548 19876 22192 19904
rect 22186 19864 22192 19876
rect 22244 19864 22250 19916
rect 13357 19839 13415 19845
rect 13357 19836 13369 19839
rect 12032 19808 13369 19836
rect 12032 19796 12038 19808
rect 13357 19805 13369 19808
rect 13403 19805 13415 19839
rect 13357 19799 13415 19805
rect 13446 19796 13452 19848
rect 13504 19796 13510 19848
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 11425 19771 11483 19777
rect 11425 19737 11437 19771
rect 11471 19768 11483 19771
rect 11606 19768 11612 19780
rect 11471 19740 11612 19768
rect 11471 19737 11483 19740
rect 11425 19731 11483 19737
rect 11606 19728 11612 19740
rect 11664 19768 11670 19780
rect 12713 19771 12771 19777
rect 12713 19768 12725 19771
rect 11664 19740 12725 19768
rect 11664 19728 11670 19740
rect 12713 19737 12725 19740
rect 12759 19768 12771 19771
rect 13464 19768 13492 19796
rect 12759 19740 13492 19768
rect 13541 19771 13599 19777
rect 12759 19737 12771 19740
rect 12713 19731 12771 19737
rect 13541 19737 13553 19771
rect 13587 19737 13599 19771
rect 13541 19731 13599 19737
rect 1578 19660 1584 19712
rect 1636 19660 1642 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7616 19672 7757 19700
rect 7616 19660 7622 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 12069 19703 12127 19709
rect 12069 19669 12081 19703
rect 12115 19700 12127 19703
rect 12618 19700 12624 19712
rect 12115 19672 12624 19700
rect 12115 19669 12127 19672
rect 12069 19663 12127 19669
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 13081 19703 13139 19709
rect 13081 19669 13093 19703
rect 13127 19700 13139 19703
rect 13556 19700 13584 19731
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 13740 19768 13768 19799
rect 13814 19796 13820 19848
rect 13872 19796 13878 19848
rect 15838 19796 15844 19848
rect 15896 19796 15902 19848
rect 20349 19839 20407 19845
rect 20349 19805 20361 19839
rect 20395 19805 20407 19839
rect 20349 19799 20407 19805
rect 15856 19768 15884 19796
rect 16761 19771 16819 19777
rect 16761 19768 16773 19771
rect 13688 19740 15884 19768
rect 16684 19740 16773 19768
rect 13688 19728 13694 19740
rect 14366 19700 14372 19712
rect 13127 19672 14372 19700
rect 13127 19669 13139 19672
rect 13081 19663 13139 19669
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 15473 19703 15531 19709
rect 15473 19669 15485 19703
rect 15519 19700 15531 19703
rect 15562 19700 15568 19712
rect 15519 19672 15568 19700
rect 15519 19669 15531 19672
rect 15473 19663 15531 19669
rect 15562 19660 15568 19672
rect 15620 19660 15626 19712
rect 16574 19660 16580 19712
rect 16632 19700 16638 19712
rect 16684 19709 16712 19740
rect 16761 19737 16773 19740
rect 16807 19737 16819 19771
rect 16761 19731 16819 19737
rect 20364 19712 20392 19799
rect 20622 19796 20628 19848
rect 20680 19796 20686 19848
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19836 22155 19839
rect 22370 19836 22376 19848
rect 22143 19808 22376 19836
rect 22143 19805 22155 19808
rect 22097 19799 22155 19805
rect 22370 19796 22376 19808
rect 22428 19796 22434 19848
rect 22557 19839 22615 19845
rect 22557 19805 22569 19839
rect 22603 19836 22615 19839
rect 22646 19836 22652 19848
rect 22603 19808 22652 19836
rect 22603 19805 22615 19808
rect 22557 19799 22615 19805
rect 22646 19796 22652 19808
rect 22704 19796 22710 19848
rect 22848 19845 22876 19944
rect 23400 19913 23428 19944
rect 27154 19932 27160 19944
rect 27212 19932 27218 19984
rect 23385 19907 23443 19913
rect 23385 19873 23397 19907
rect 23431 19873 23443 19907
rect 23385 19867 23443 19873
rect 24213 19907 24271 19913
rect 24213 19873 24225 19907
rect 24259 19904 24271 19907
rect 24854 19904 24860 19916
rect 24259 19876 24860 19904
rect 24259 19873 24271 19876
rect 24213 19867 24271 19873
rect 24854 19864 24860 19876
rect 24912 19904 24918 19916
rect 24912 19876 25452 19904
rect 24912 19864 24918 19876
rect 25424 19845 25452 19876
rect 25774 19864 25780 19916
rect 25832 19864 25838 19916
rect 27264 19913 27292 20012
rect 30098 20000 30104 20052
rect 30156 20000 30162 20052
rect 31665 20043 31723 20049
rect 31665 20040 31677 20043
rect 31220 20012 31677 20040
rect 27249 19907 27307 19913
rect 27249 19873 27261 19907
rect 27295 19873 27307 19907
rect 27249 19867 27307 19873
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19805 22891 19839
rect 25225 19839 25283 19845
rect 22833 19799 22891 19805
rect 20438 19728 20444 19780
rect 20496 19768 20502 19780
rect 21085 19771 21143 19777
rect 21085 19768 21097 19771
rect 20496 19740 21097 19768
rect 20496 19728 20502 19740
rect 21085 19737 21097 19740
rect 21131 19737 21143 19771
rect 21085 19731 21143 19737
rect 21269 19771 21327 19777
rect 21269 19737 21281 19771
rect 21315 19737 21327 19771
rect 21269 19731 21327 19737
rect 22465 19771 22523 19777
rect 22465 19737 22477 19771
rect 22511 19768 22523 19771
rect 23308 19768 23336 19822
rect 25225 19805 25237 19839
rect 25271 19805 25283 19839
rect 25225 19799 25283 19805
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 22511 19740 23336 19768
rect 22511 19737 22523 19740
rect 22465 19731 22523 19737
rect 16669 19703 16727 19709
rect 16669 19700 16681 19703
rect 16632 19672 16681 19700
rect 16632 19660 16638 19672
rect 16669 19669 16681 19672
rect 16715 19669 16727 19703
rect 16669 19663 16727 19669
rect 16971 19703 17029 19709
rect 16971 19669 16983 19703
rect 17017 19700 17029 19703
rect 17494 19700 17500 19712
rect 17017 19672 17500 19700
rect 17017 19669 17029 19672
rect 16971 19663 17029 19669
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 20346 19660 20352 19712
rect 20404 19700 20410 19712
rect 21284 19700 21312 19731
rect 23750 19728 23756 19780
rect 23808 19728 23814 19780
rect 20404 19672 21312 19700
rect 23017 19703 23075 19709
rect 20404 19660 20410 19672
rect 23017 19669 23029 19703
rect 23063 19700 23075 19703
rect 23768 19700 23796 19728
rect 25240 19712 25268 19799
rect 25590 19796 25596 19848
rect 25648 19796 25654 19848
rect 25685 19839 25743 19845
rect 25685 19805 25697 19839
rect 25731 19836 25743 19839
rect 25792 19836 25820 19864
rect 26881 19839 26939 19845
rect 26881 19836 26893 19839
rect 25731 19808 25820 19836
rect 26804 19808 26893 19836
rect 25731 19805 25743 19808
rect 25685 19799 25743 19805
rect 25314 19728 25320 19780
rect 25372 19768 25378 19780
rect 26237 19771 26295 19777
rect 26237 19768 26249 19771
rect 25372 19740 26249 19768
rect 25372 19728 25378 19740
rect 26237 19737 26249 19740
rect 26283 19768 26295 19771
rect 26804 19768 26832 19808
rect 26881 19805 26893 19808
rect 26927 19805 26939 19839
rect 26881 19799 26939 19805
rect 27065 19839 27123 19845
rect 27065 19805 27077 19839
rect 27111 19836 27123 19839
rect 27154 19836 27160 19848
rect 27111 19808 27160 19836
rect 27111 19805 27123 19808
rect 27065 19799 27123 19805
rect 27154 19796 27160 19808
rect 27212 19796 27218 19848
rect 27341 19839 27399 19845
rect 27341 19805 27353 19839
rect 27387 19805 27399 19839
rect 27341 19799 27399 19805
rect 29733 19839 29791 19845
rect 29733 19805 29745 19839
rect 29779 19836 29791 19839
rect 30116 19836 30144 20000
rect 31110 19864 31116 19916
rect 31168 19864 31174 19916
rect 31220 19845 31248 20012
rect 31665 20009 31677 20012
rect 31711 20009 31723 20043
rect 31665 20003 31723 20009
rect 32030 20000 32036 20052
rect 32088 20000 32094 20052
rect 32490 20000 32496 20052
rect 32548 20000 32554 20052
rect 33226 20000 33232 20052
rect 33284 20040 33290 20052
rect 33321 20043 33379 20049
rect 33321 20040 33333 20043
rect 33284 20012 33333 20040
rect 33284 20000 33290 20012
rect 33321 20009 33333 20012
rect 33367 20009 33379 20043
rect 33321 20003 33379 20009
rect 31573 19975 31631 19981
rect 31573 19941 31585 19975
rect 31619 19972 31631 19975
rect 32508 19972 32536 20000
rect 31619 19944 32536 19972
rect 31619 19941 31631 19944
rect 31573 19935 31631 19941
rect 31386 19864 31392 19916
rect 31444 19904 31450 19916
rect 31757 19907 31815 19913
rect 31757 19904 31769 19907
rect 31444 19876 31769 19904
rect 31444 19864 31450 19876
rect 31757 19873 31769 19876
rect 31803 19873 31815 19907
rect 31757 19867 31815 19873
rect 31205 19839 31263 19845
rect 31205 19836 31217 19839
rect 29779 19808 30144 19836
rect 30208 19808 31217 19836
rect 29779 19805 29791 19808
rect 29733 19799 29791 19805
rect 26283 19740 26832 19768
rect 26283 19737 26295 19740
rect 26237 19731 26295 19737
rect 26804 19712 26832 19740
rect 26973 19771 27031 19777
rect 26973 19737 26985 19771
rect 27019 19768 27031 19771
rect 27356 19768 27384 19799
rect 27019 19740 27384 19768
rect 27019 19737 27031 19740
rect 26973 19731 27031 19737
rect 30208 19712 30236 19808
rect 31205 19805 31217 19808
rect 31251 19805 31263 19839
rect 31665 19839 31723 19845
rect 31665 19836 31677 19839
rect 31205 19799 31263 19805
rect 31496 19808 31677 19836
rect 31496 19712 31524 19808
rect 31665 19805 31677 19808
rect 31711 19805 31723 19839
rect 31665 19799 31723 19805
rect 33134 19796 33140 19848
rect 33192 19836 33198 19848
rect 33229 19839 33287 19845
rect 33229 19836 33241 19839
rect 33192 19808 33241 19836
rect 33192 19796 33198 19808
rect 33229 19805 33241 19808
rect 33275 19805 33287 19839
rect 33229 19799 33287 19805
rect 23063 19672 23796 19700
rect 23063 19669 23075 19672
rect 23017 19663 23075 19669
rect 25222 19660 25228 19712
rect 25280 19660 25286 19712
rect 25590 19660 25596 19712
rect 25648 19700 25654 19712
rect 26053 19703 26111 19709
rect 26053 19700 26065 19703
rect 25648 19672 26065 19700
rect 25648 19660 25654 19672
rect 26053 19669 26065 19672
rect 26099 19669 26111 19703
rect 26053 19663 26111 19669
rect 26786 19660 26792 19712
rect 26844 19660 26850 19712
rect 27706 19660 27712 19712
rect 27764 19660 27770 19712
rect 29641 19703 29699 19709
rect 29641 19669 29653 19703
rect 29687 19700 29699 19703
rect 29730 19700 29736 19712
rect 29687 19672 29736 19700
rect 29687 19669 29699 19672
rect 29641 19663 29699 19669
rect 29730 19660 29736 19672
rect 29788 19660 29794 19712
rect 30190 19660 30196 19712
rect 30248 19660 30254 19712
rect 31478 19660 31484 19712
rect 31536 19660 31542 19712
rect 33137 19703 33195 19709
rect 33137 19669 33149 19703
rect 33183 19700 33195 19703
rect 33244 19700 33272 19799
rect 33594 19700 33600 19712
rect 33183 19672 33600 19700
rect 33183 19669 33195 19672
rect 33137 19663 33195 19669
rect 33594 19660 33600 19672
rect 33652 19660 33658 19712
rect 1104 19610 35236 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 35236 19610
rect 1104 19536 35236 19558
rect 9766 19456 9772 19508
rect 9824 19496 9830 19508
rect 9861 19499 9919 19505
rect 9861 19496 9873 19499
rect 9824 19468 9873 19496
rect 9824 19456 9830 19468
rect 9861 19465 9873 19468
rect 9907 19465 9919 19499
rect 9861 19459 9919 19465
rect 10042 19456 10048 19508
rect 10100 19496 10106 19508
rect 10229 19499 10287 19505
rect 10229 19496 10241 19499
rect 10100 19468 10241 19496
rect 10100 19456 10106 19468
rect 10229 19465 10241 19468
rect 10275 19465 10287 19499
rect 10229 19459 10287 19465
rect 11974 19456 11980 19508
rect 12032 19456 12038 19508
rect 12066 19456 12072 19508
rect 12124 19456 12130 19508
rect 12158 19456 12164 19508
rect 12216 19496 12222 19508
rect 13354 19496 13360 19508
rect 12216 19468 13360 19496
rect 12216 19456 12222 19468
rect 13354 19456 13360 19468
rect 13412 19456 13418 19508
rect 13814 19456 13820 19508
rect 13872 19456 13878 19508
rect 15562 19456 15568 19508
rect 15620 19496 15626 19508
rect 16114 19496 16120 19508
rect 15620 19468 16120 19496
rect 15620 19456 15626 19468
rect 16114 19456 16120 19468
rect 16172 19496 16178 19508
rect 16485 19499 16543 19505
rect 16485 19496 16497 19499
rect 16172 19468 16497 19496
rect 16172 19456 16178 19468
rect 16485 19465 16497 19468
rect 16531 19496 16543 19499
rect 16574 19496 16580 19508
rect 16531 19468 16580 19496
rect 16531 19465 16543 19468
rect 16485 19459 16543 19465
rect 16574 19456 16580 19468
rect 16632 19456 16638 19508
rect 16666 19456 16672 19508
rect 16724 19496 16730 19508
rect 16853 19499 16911 19505
rect 16853 19496 16865 19499
rect 16724 19468 16865 19496
rect 16724 19456 16730 19468
rect 16853 19465 16865 19468
rect 16899 19465 16911 19499
rect 16853 19459 16911 19465
rect 17494 19456 17500 19508
rect 17552 19456 17558 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18012 19468 19472 19496
rect 18012 19456 18018 19468
rect 9953 19431 10011 19437
rect 9953 19428 9965 19431
rect 9784 19400 9965 19428
rect 9784 19292 9812 19400
rect 9953 19397 9965 19400
rect 9999 19397 10011 19431
rect 14921 19431 14979 19437
rect 14921 19428 14933 19431
rect 9953 19391 10011 19397
rect 11440 19400 14933 19428
rect 9858 19320 9864 19372
rect 9916 19320 9922 19372
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19329 10103 19363
rect 10045 19323 10103 19329
rect 9232 19264 9812 19292
rect 9876 19292 9904 19320
rect 10060 19292 10088 19323
rect 10505 19295 10563 19301
rect 10505 19292 10517 19295
rect 9876 19264 10517 19292
rect 9232 19168 9260 19264
rect 10505 19261 10517 19264
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 10962 19252 10968 19304
rect 11020 19292 11026 19304
rect 11440 19292 11468 19400
rect 11624 19332 11928 19360
rect 11624 19304 11652 19332
rect 11020 19264 11468 19292
rect 11020 19252 11026 19264
rect 11514 19252 11520 19304
rect 11572 19252 11578 19304
rect 11606 19252 11612 19304
rect 11664 19252 11670 19304
rect 11701 19295 11759 19301
rect 11701 19261 11713 19295
rect 11747 19261 11759 19295
rect 11701 19255 11759 19261
rect 9585 19227 9643 19233
rect 9585 19193 9597 19227
rect 9631 19224 9643 19227
rect 9674 19224 9680 19236
rect 9631 19196 9680 19224
rect 9631 19193 9643 19196
rect 9585 19187 9643 19193
rect 9674 19184 9680 19196
rect 9732 19224 9738 19236
rect 11716 19224 11744 19255
rect 11790 19252 11796 19304
rect 11848 19252 11854 19304
rect 11900 19292 11928 19332
rect 12434 19320 12440 19372
rect 12492 19320 12498 19372
rect 12618 19320 12624 19372
rect 12676 19320 12682 19372
rect 12710 19320 12716 19372
rect 12768 19320 12774 19372
rect 12912 19369 12940 19400
rect 14921 19397 14933 19400
rect 14967 19428 14979 19431
rect 15194 19428 15200 19440
rect 14967 19400 15200 19428
rect 14967 19397 14979 19400
rect 14921 19391 14979 19397
rect 15194 19388 15200 19400
rect 15252 19388 15258 19440
rect 16761 19431 16819 19437
rect 16761 19428 16773 19431
rect 15488 19400 16773 19428
rect 12897 19363 12955 19369
rect 12897 19329 12909 19363
rect 12943 19329 12955 19363
rect 13725 19363 13783 19369
rect 13725 19360 13737 19363
rect 12897 19323 12955 19329
rect 13556 19332 13737 19360
rect 12158 19292 12164 19304
rect 11900 19264 12164 19292
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12342 19252 12348 19304
rect 12400 19292 12406 19304
rect 12400 19252 12434 19292
rect 12253 19227 12311 19233
rect 12253 19224 12265 19227
rect 9732 19196 11560 19224
rect 11716 19196 12265 19224
rect 9732 19184 9738 19196
rect 9214 19116 9220 19168
rect 9272 19116 9278 19168
rect 10965 19159 11023 19165
rect 10965 19125 10977 19159
rect 11011 19156 11023 19159
rect 11146 19156 11152 19168
rect 11011 19128 11152 19156
rect 11011 19125 11023 19128
rect 10965 19119 11023 19125
rect 11146 19116 11152 19128
rect 11204 19156 11210 19168
rect 11241 19159 11299 19165
rect 11241 19156 11253 19159
rect 11204 19128 11253 19156
rect 11204 19116 11210 19128
rect 11241 19125 11253 19128
rect 11287 19125 11299 19159
rect 11532 19156 11560 19196
rect 12253 19193 12265 19196
rect 12299 19193 12311 19227
rect 12253 19187 12311 19193
rect 12406 19156 12434 19252
rect 12526 19184 12532 19236
rect 12584 19184 12590 19236
rect 13556 19233 13584 19332
rect 13725 19329 13737 19332
rect 13771 19329 13783 19363
rect 13725 19323 13783 19329
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 15105 19363 15163 19369
rect 13955 19332 14320 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 13541 19227 13599 19233
rect 13541 19224 13553 19227
rect 12636 19196 13553 19224
rect 12636 19168 12664 19196
rect 13541 19193 13553 19196
rect 13587 19193 13599 19227
rect 13541 19187 13599 19193
rect 12618 19156 12624 19168
rect 11532 19128 12624 19156
rect 11241 19119 11299 19125
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 13262 19116 13268 19168
rect 13320 19116 13326 19168
rect 14292 19165 14320 19332
rect 15105 19329 15117 19363
rect 15151 19360 15163 19363
rect 15286 19360 15292 19372
rect 15151 19332 15292 19360
rect 15151 19329 15163 19332
rect 15105 19323 15163 19329
rect 15286 19320 15292 19332
rect 15344 19320 15350 19372
rect 15378 19252 15384 19304
rect 15436 19292 15442 19304
rect 15488 19301 15516 19400
rect 16761 19397 16773 19400
rect 16807 19397 16819 19431
rect 19444 19428 19472 19468
rect 20346 19456 20352 19508
rect 20404 19496 20410 19508
rect 20404 19468 22140 19496
rect 20404 19456 20410 19468
rect 21266 19428 21272 19440
rect 16761 19391 16819 19397
rect 18800 19400 19380 19428
rect 19444 19400 21272 19428
rect 15746 19320 15752 19372
rect 15804 19320 15810 19372
rect 16666 19360 16672 19372
rect 16592 19332 16672 19360
rect 16592 19304 16620 19332
rect 16666 19320 16672 19332
rect 16724 19320 16730 19372
rect 17954 19360 17960 19372
rect 16960 19332 17960 19360
rect 15473 19295 15531 19301
rect 15473 19292 15485 19295
rect 15436 19264 15485 19292
rect 15436 19252 15442 19264
rect 15473 19261 15485 19264
rect 15519 19261 15531 19295
rect 15473 19255 15531 19261
rect 15654 19252 15660 19304
rect 15712 19252 15718 19304
rect 16574 19252 16580 19304
rect 16632 19252 16638 19304
rect 16853 19295 16911 19301
rect 16853 19261 16865 19295
rect 16899 19261 16911 19295
rect 16853 19255 16911 19261
rect 15289 19227 15347 19233
rect 15289 19193 15301 19227
rect 15335 19224 15347 19227
rect 16880 19224 16908 19255
rect 15335 19196 16908 19224
rect 15335 19193 15347 19196
rect 15289 19187 15347 19193
rect 14277 19159 14335 19165
rect 14277 19125 14289 19159
rect 14323 19156 14335 19159
rect 14734 19156 14740 19168
rect 14323 19128 14740 19156
rect 14323 19125 14335 19128
rect 14277 19119 14335 19125
rect 14734 19116 14740 19128
rect 14792 19116 14798 19168
rect 15194 19116 15200 19168
rect 15252 19156 15258 19168
rect 15930 19156 15936 19168
rect 15252 19128 15936 19156
rect 15252 19116 15258 19128
rect 15930 19116 15936 19128
rect 15988 19116 15994 19168
rect 16117 19159 16175 19165
rect 16117 19125 16129 19159
rect 16163 19156 16175 19159
rect 16960 19156 16988 19332
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18046 19320 18052 19372
rect 18104 19360 18110 19372
rect 18800 19369 18828 19400
rect 18785 19363 18843 19369
rect 18104 19332 18276 19360
rect 18104 19320 18110 19332
rect 17678 19252 17684 19304
rect 17736 19252 17742 19304
rect 17770 19252 17776 19304
rect 17828 19252 17834 19304
rect 18138 19252 18144 19304
rect 18196 19252 18202 19304
rect 18248 19292 18276 19332
rect 18785 19329 18797 19363
rect 18831 19329 18843 19363
rect 18785 19323 18843 19329
rect 18874 19320 18880 19372
rect 18932 19320 18938 19372
rect 19061 19363 19119 19369
rect 19061 19329 19073 19363
rect 19107 19329 19119 19363
rect 19352 19360 19380 19400
rect 21266 19388 21272 19400
rect 21324 19388 21330 19440
rect 20070 19360 20076 19372
rect 19352 19332 20076 19360
rect 19061 19323 19119 19329
rect 18966 19292 18972 19304
rect 18248 19264 18972 19292
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 16163 19128 16988 19156
rect 16163 19125 16175 19128
rect 16117 19119 16175 19125
rect 17310 19116 17316 19168
rect 17368 19156 17374 19168
rect 18322 19156 18328 19168
rect 17368 19128 18328 19156
rect 17368 19116 17374 19128
rect 18322 19116 18328 19128
rect 18380 19116 18386 19168
rect 18414 19116 18420 19168
rect 18472 19156 18478 19168
rect 19076 19156 19104 19323
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 22112 19369 22140 19468
rect 22186 19456 22192 19508
rect 22244 19496 22250 19508
rect 23566 19496 23572 19508
rect 22244 19468 23572 19496
rect 22244 19456 22250 19468
rect 23566 19456 23572 19468
rect 23624 19456 23630 19508
rect 25314 19456 25320 19508
rect 25372 19456 25378 19508
rect 25498 19505 25504 19508
rect 25494 19459 25504 19505
rect 25498 19456 25504 19459
rect 25556 19456 25562 19508
rect 28350 19456 28356 19508
rect 28408 19456 28414 19508
rect 30190 19456 30196 19508
rect 30248 19456 30254 19508
rect 31110 19456 31116 19508
rect 31168 19456 31174 19508
rect 25332 19428 25360 19456
rect 25409 19431 25467 19437
rect 25409 19428 25421 19431
rect 25332 19400 25421 19428
rect 25409 19397 25421 19400
rect 25455 19397 25467 19431
rect 25409 19391 25467 19397
rect 27706 19388 27712 19440
rect 27764 19428 27770 19440
rect 28721 19431 28779 19437
rect 28721 19428 28733 19431
rect 27764 19400 28733 19428
rect 27764 19388 27770 19400
rect 28721 19397 28733 19400
rect 28767 19397 28779 19431
rect 28721 19391 28779 19397
rect 29730 19388 29736 19440
rect 29788 19388 29794 19440
rect 31386 19388 31392 19440
rect 31444 19388 31450 19440
rect 31388 19385 31446 19388
rect 20625 19363 20683 19369
rect 20625 19360 20637 19363
rect 20496 19332 20637 19360
rect 20496 19320 20502 19332
rect 20625 19329 20637 19332
rect 20671 19329 20683 19363
rect 20625 19323 20683 19329
rect 22097 19363 22155 19369
rect 22097 19329 22109 19363
rect 22143 19329 22155 19363
rect 22097 19323 22155 19329
rect 25314 19320 25320 19372
rect 25372 19320 25378 19372
rect 25590 19360 25596 19372
rect 25424 19332 25596 19360
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 22005 19295 22063 19301
rect 22005 19292 22017 19295
rect 20579 19264 20668 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 20640 19168 20668 19264
rect 21008 19264 22017 19292
rect 21008 19233 21036 19264
rect 22005 19261 22017 19264
rect 22051 19261 22063 19295
rect 22005 19255 22063 19261
rect 22925 19295 22983 19301
rect 22925 19261 22937 19295
rect 22971 19292 22983 19295
rect 24670 19292 24676 19304
rect 22971 19264 24676 19292
rect 22971 19261 22983 19264
rect 22925 19255 22983 19261
rect 24670 19252 24676 19264
rect 24728 19292 24734 19304
rect 25424 19292 25452 19332
rect 25590 19320 25596 19332
rect 25648 19320 25654 19372
rect 28350 19320 28356 19372
rect 28408 19360 28414 19372
rect 28445 19363 28503 19369
rect 28445 19360 28457 19363
rect 28408 19332 28457 19360
rect 28408 19320 28414 19332
rect 28445 19329 28457 19332
rect 28491 19329 28503 19363
rect 31388 19351 31400 19385
rect 31434 19351 31446 19385
rect 31388 19345 31446 19351
rect 28445 19323 28503 19329
rect 24728 19264 25452 19292
rect 24728 19252 24734 19264
rect 31018 19252 31024 19304
rect 31076 19292 31082 19304
rect 31113 19295 31171 19301
rect 31113 19292 31125 19295
rect 31076 19264 31125 19292
rect 31076 19252 31082 19264
rect 31113 19261 31125 19264
rect 31159 19292 31171 19295
rect 31159 19264 31754 19292
rect 31159 19261 31171 19264
rect 31113 19255 31171 19261
rect 20993 19227 21051 19233
rect 20993 19193 21005 19227
rect 21039 19193 21051 19227
rect 31726 19224 31754 19264
rect 32214 19224 32220 19236
rect 31726 19196 32220 19224
rect 20993 19187 21051 19193
rect 32214 19184 32220 19196
rect 32272 19184 32278 19236
rect 18472 19128 19104 19156
rect 18472 19116 18478 19128
rect 19242 19116 19248 19168
rect 19300 19116 19306 19168
rect 20622 19116 20628 19168
rect 20680 19116 20686 19168
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 23198 19156 23204 19168
rect 22704 19128 23204 19156
rect 22704 19116 22710 19128
rect 23198 19116 23204 19128
rect 23256 19116 23262 19168
rect 31297 19159 31355 19165
rect 31297 19125 31309 19159
rect 31343 19156 31355 19159
rect 31478 19156 31484 19168
rect 31343 19128 31484 19156
rect 31343 19125 31355 19128
rect 31297 19119 31355 19125
rect 31478 19116 31484 19128
rect 31536 19116 31542 19168
rect 1104 19066 35248 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 35248 19066
rect 1104 18992 35248 19014
rect 12066 18912 12072 18964
rect 12124 18912 12130 18964
rect 12529 18955 12587 18961
rect 12529 18921 12541 18955
rect 12575 18952 12587 18955
rect 12710 18952 12716 18964
rect 12575 18924 12716 18952
rect 12575 18921 12587 18924
rect 12529 18915 12587 18921
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 13262 18912 13268 18964
rect 13320 18952 13326 18964
rect 13538 18952 13544 18964
rect 13320 18924 13544 18952
rect 13320 18912 13326 18924
rect 13538 18912 13544 18924
rect 13596 18952 13602 18964
rect 14369 18955 14427 18961
rect 14369 18952 14381 18955
rect 13596 18924 14381 18952
rect 13596 18912 13602 18924
rect 14369 18921 14381 18924
rect 14415 18952 14427 18955
rect 14458 18952 14464 18964
rect 14415 18924 14464 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 14458 18912 14464 18924
rect 14516 18952 14522 18964
rect 14921 18955 14979 18961
rect 14921 18952 14933 18955
rect 14516 18924 14933 18952
rect 14516 18912 14522 18924
rect 14921 18921 14933 18924
rect 14967 18952 14979 18955
rect 15562 18952 15568 18964
rect 14967 18924 15568 18952
rect 14967 18921 14979 18924
rect 14921 18915 14979 18921
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 15654 18912 15660 18964
rect 15712 18912 15718 18964
rect 15746 18912 15752 18964
rect 15804 18952 15810 18964
rect 16117 18955 16175 18961
rect 16117 18952 16129 18955
rect 15804 18924 16129 18952
rect 15804 18912 15810 18924
rect 16117 18921 16129 18924
rect 16163 18921 16175 18955
rect 16117 18915 16175 18921
rect 17129 18955 17187 18961
rect 17129 18921 17141 18955
rect 17175 18952 17187 18955
rect 17678 18952 17684 18964
rect 17175 18924 17684 18952
rect 17175 18921 17187 18924
rect 17129 18915 17187 18921
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 18046 18912 18052 18964
rect 18104 18912 18110 18964
rect 19058 18912 19064 18964
rect 19116 18912 19122 18964
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 19300 18924 22094 18952
rect 19300 18912 19306 18924
rect 9493 18887 9551 18893
rect 9493 18853 9505 18887
rect 9539 18884 9551 18887
rect 12084 18884 12112 18912
rect 9539 18856 9812 18884
rect 12084 18856 12296 18884
rect 9539 18853 9551 18856
rect 9493 18847 9551 18853
rect 9416 18788 9720 18816
rect 9416 18757 9444 18788
rect 9692 18760 9720 18788
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 9508 18612 9536 18711
rect 9674 18708 9680 18760
rect 9732 18708 9738 18760
rect 9784 18757 9812 18856
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 12268 18825 12296 18856
rect 12161 18819 12219 18825
rect 12161 18816 12173 18819
rect 11572 18788 12173 18816
rect 11572 18776 11578 18788
rect 12161 18785 12173 18788
rect 12207 18785 12219 18819
rect 12161 18779 12219 18785
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18785 12311 18819
rect 12253 18779 12311 18785
rect 9769 18751 9827 18757
rect 9769 18717 9781 18751
rect 9815 18717 9827 18751
rect 9769 18711 9827 18717
rect 10318 18708 10324 18760
rect 10376 18708 10382 18760
rect 12069 18751 12127 18757
rect 12069 18748 12081 18751
rect 11992 18720 12081 18748
rect 10962 18640 10968 18692
rect 11020 18640 11026 18692
rect 11992 18680 12020 18720
rect 12069 18717 12081 18720
rect 12115 18717 12127 18751
rect 12176 18748 12204 18779
rect 12342 18776 12348 18828
rect 12400 18776 12406 18828
rect 13280 18748 13308 18912
rect 15841 18887 15899 18893
rect 15841 18853 15853 18887
rect 15887 18884 15899 18887
rect 16574 18884 16580 18896
rect 15887 18856 16580 18884
rect 15887 18853 15899 18856
rect 15841 18847 15899 18853
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 18064 18884 18092 18912
rect 17604 18856 18092 18884
rect 15286 18776 15292 18828
rect 15344 18816 15350 18828
rect 16761 18819 16819 18825
rect 15344 18788 16068 18816
rect 15344 18776 15350 18788
rect 12176 18720 13308 18748
rect 12069 18711 12127 18717
rect 15194 18708 15200 18760
rect 15252 18748 15258 18760
rect 15764 18757 15884 18758
rect 15749 18751 15884 18757
rect 15252 18720 15332 18748
rect 15252 18708 15258 18720
rect 12250 18680 12256 18692
rect 11992 18652 12256 18680
rect 12250 18640 12256 18652
rect 12308 18680 12314 18692
rect 14366 18680 14372 18692
rect 12308 18652 14372 18680
rect 12308 18640 12314 18652
rect 14366 18640 14372 18652
rect 14424 18640 14430 18692
rect 15102 18640 15108 18692
rect 15160 18640 15166 18692
rect 15304 18689 15332 18720
rect 15749 18717 15761 18751
rect 15795 18730 15884 18751
rect 15795 18717 15807 18730
rect 15749 18711 15807 18717
rect 15289 18683 15347 18689
rect 15289 18649 15301 18683
rect 15335 18649 15347 18683
rect 15289 18643 15347 18649
rect 15473 18683 15531 18689
rect 15473 18649 15485 18683
rect 15519 18680 15531 18683
rect 15856 18680 15884 18730
rect 15930 18708 15936 18760
rect 15988 18708 15994 18760
rect 16040 18757 16068 18788
rect 16761 18785 16773 18819
rect 16807 18816 16819 18819
rect 17604 18816 17632 18856
rect 18966 18844 18972 18896
rect 19024 18884 19030 18896
rect 19024 18856 20300 18884
rect 19024 18844 19030 18856
rect 16807 18788 17632 18816
rect 16807 18785 16819 18788
rect 16761 18779 16819 18785
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18717 16083 18751
rect 16025 18711 16083 18717
rect 16209 18751 16267 18757
rect 16209 18717 16221 18751
rect 16255 18717 16267 18751
rect 16776 18748 16804 18779
rect 17954 18776 17960 18828
rect 18012 18816 18018 18828
rect 19245 18819 19303 18825
rect 19245 18816 19257 18819
rect 18012 18788 19257 18816
rect 18012 18776 18018 18788
rect 16209 18711 16267 18717
rect 16316 18720 16804 18748
rect 15519 18652 15884 18680
rect 15948 18680 15976 18708
rect 16224 18680 16252 18711
rect 15948 18652 16252 18680
rect 15519 18649 15531 18652
rect 15473 18643 15531 18649
rect 9858 18612 9864 18624
rect 9508 18584 9864 18612
rect 9858 18572 9864 18584
rect 9916 18572 9922 18624
rect 11698 18572 11704 18624
rect 11756 18612 11762 18624
rect 12342 18612 12348 18624
rect 11756 18584 12348 18612
rect 11756 18572 11762 18584
rect 12342 18572 12348 18584
rect 12400 18612 12406 18624
rect 13078 18612 13084 18624
rect 12400 18584 13084 18612
rect 12400 18572 12406 18584
rect 13078 18572 13084 18584
rect 13136 18572 13142 18624
rect 13173 18615 13231 18621
rect 13173 18581 13185 18615
rect 13219 18612 13231 18615
rect 13446 18612 13452 18624
rect 13219 18584 13452 18612
rect 13219 18581 13231 18584
rect 13173 18575 13231 18581
rect 13446 18572 13452 18584
rect 13504 18572 13510 18624
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 14734 18612 14740 18624
rect 13964 18584 14740 18612
rect 13964 18572 13970 18584
rect 14734 18572 14740 18584
rect 14792 18572 14798 18624
rect 15120 18612 15148 18640
rect 15488 18612 15516 18643
rect 15120 18584 15516 18612
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16316 18612 16344 18720
rect 17034 18708 17040 18760
rect 17092 18708 17098 18760
rect 17218 18708 17224 18760
rect 17276 18708 17282 18760
rect 18248 18757 18276 18788
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18524 18757 18552 18788
rect 19245 18785 19257 18788
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19628 18825 19656 18856
rect 19613 18819 19671 18825
rect 19392 18788 19564 18816
rect 19392 18776 19398 18788
rect 18417 18751 18475 18757
rect 18417 18748 18429 18751
rect 18380 18720 18429 18748
rect 18380 18708 18386 18720
rect 18417 18717 18429 18720
rect 18463 18717 18475 18751
rect 18417 18711 18475 18717
rect 18509 18751 18567 18757
rect 18509 18717 18521 18751
rect 18555 18717 18567 18751
rect 18509 18711 18567 18717
rect 18877 18751 18935 18757
rect 18877 18717 18889 18751
rect 18923 18748 18935 18751
rect 19426 18748 19432 18760
rect 18923 18720 19432 18748
rect 18923 18717 18935 18720
rect 18877 18711 18935 18717
rect 16574 18640 16580 18692
rect 16632 18680 16638 18692
rect 17236 18680 17264 18708
rect 16632 18652 17264 18680
rect 18432 18680 18460 18711
rect 19426 18708 19432 18720
rect 19484 18708 19490 18760
rect 19536 18748 19564 18788
rect 19613 18785 19625 18819
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18816 19947 18819
rect 20272 18816 20300 18856
rect 20346 18844 20352 18896
rect 20404 18844 20410 18896
rect 22066 18884 22094 18924
rect 25314 18912 25320 18964
rect 25372 18952 25378 18964
rect 25501 18955 25559 18961
rect 25501 18952 25513 18955
rect 25372 18924 25513 18952
rect 25372 18912 25378 18924
rect 25501 18921 25513 18924
rect 25547 18952 25559 18955
rect 25547 18924 26188 18952
rect 25547 18921 25559 18924
rect 25501 18915 25559 18921
rect 25961 18887 26019 18893
rect 22066 18856 24992 18884
rect 24964 18816 24992 18856
rect 25961 18853 25973 18887
rect 26007 18853 26019 18887
rect 26160 18884 26188 18924
rect 26786 18912 26792 18964
rect 26844 18912 26850 18964
rect 31297 18955 31355 18961
rect 31297 18921 31309 18955
rect 31343 18952 31355 18955
rect 31386 18952 31392 18964
rect 31343 18924 31392 18952
rect 31343 18921 31355 18924
rect 31297 18915 31355 18921
rect 31386 18912 31392 18924
rect 31444 18912 31450 18964
rect 27154 18884 27160 18896
rect 26160 18856 27160 18884
rect 25961 18847 26019 18853
rect 25976 18816 26004 18847
rect 27154 18844 27160 18856
rect 27212 18884 27218 18896
rect 27709 18887 27767 18893
rect 27709 18884 27721 18887
rect 27212 18856 27721 18884
rect 27212 18844 27218 18856
rect 27709 18853 27721 18856
rect 27755 18853 27767 18887
rect 27709 18847 27767 18853
rect 28629 18887 28687 18893
rect 28629 18853 28641 18887
rect 28675 18853 28687 18887
rect 28629 18847 28687 18853
rect 27893 18819 27951 18825
rect 19935 18788 20208 18816
rect 20272 18788 20760 18816
rect 19935 18785 19947 18788
rect 19889 18779 19947 18785
rect 20180 18757 20208 18788
rect 20732 18760 20760 18788
rect 24964 18788 25728 18816
rect 25976 18788 27384 18816
rect 22836 18760 22888 18766
rect 19705 18751 19763 18757
rect 19705 18748 19717 18751
rect 19536 18720 19717 18748
rect 19705 18717 19717 18720
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18717 20039 18751
rect 19981 18711 20039 18717
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 18693 18683 18751 18689
rect 18693 18680 18705 18683
rect 18432 18652 18705 18680
rect 16632 18640 16638 18652
rect 18693 18649 18705 18652
rect 18739 18649 18751 18683
rect 18693 18643 18751 18649
rect 18785 18683 18843 18689
rect 18785 18649 18797 18683
rect 18831 18680 18843 18683
rect 18966 18680 18972 18692
rect 18831 18652 18972 18680
rect 18831 18649 18843 18652
rect 18785 18643 18843 18649
rect 15804 18584 16344 18612
rect 17589 18615 17647 18621
rect 15804 18572 15810 18584
rect 17589 18581 17601 18615
rect 17635 18612 17647 18615
rect 17954 18612 17960 18624
rect 17635 18584 17960 18612
rect 17635 18581 17647 18584
rect 17589 18575 17647 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18414 18572 18420 18624
rect 18472 18572 18478 18624
rect 18708 18612 18736 18643
rect 18966 18640 18972 18652
rect 19024 18640 19030 18692
rect 19058 18640 19064 18692
rect 19116 18680 19122 18692
rect 19996 18680 20024 18711
rect 20714 18708 20720 18760
rect 20772 18708 20778 18760
rect 22373 18751 22431 18757
rect 22373 18748 22385 18751
rect 22020 18720 22385 18748
rect 19116 18652 20024 18680
rect 19116 18640 19122 18652
rect 19337 18615 19395 18621
rect 19337 18612 19349 18615
rect 18708 18584 19349 18612
rect 19337 18581 19349 18584
rect 19383 18581 19395 18615
rect 19337 18575 19395 18581
rect 19426 18572 19432 18624
rect 19484 18572 19490 18624
rect 20438 18572 20444 18624
rect 20496 18612 20502 18624
rect 22020 18621 22048 18720
rect 22373 18717 22385 18720
rect 22419 18717 22431 18751
rect 22373 18711 22431 18717
rect 22554 18708 22560 18760
rect 22612 18708 22618 18760
rect 22741 18751 22799 18757
rect 22741 18717 22753 18751
rect 22787 18717 22799 18751
rect 22741 18711 22799 18717
rect 22465 18683 22523 18689
rect 22465 18649 22477 18683
rect 22511 18680 22523 18683
rect 22756 18680 22784 18711
rect 24964 18757 24992 18788
rect 25700 18757 25728 18788
rect 27356 18757 27384 18788
rect 27893 18785 27905 18819
rect 27939 18816 27951 18819
rect 28077 18819 28135 18825
rect 28077 18816 28089 18819
rect 27939 18788 28089 18816
rect 27939 18785 27951 18788
rect 27893 18779 27951 18785
rect 28077 18785 28089 18788
rect 28123 18785 28135 18819
rect 28077 18779 28135 18785
rect 24949 18751 25007 18757
rect 24949 18717 24961 18751
rect 24995 18717 25007 18751
rect 25225 18751 25283 18757
rect 25225 18748 25237 18751
rect 24949 18711 25007 18717
rect 25056 18720 25237 18748
rect 22836 18702 22888 18708
rect 22511 18652 22784 18680
rect 22511 18649 22523 18652
rect 22465 18643 22523 18649
rect 23658 18640 23664 18692
rect 23716 18680 23722 18692
rect 23753 18683 23811 18689
rect 23753 18680 23765 18683
rect 23716 18652 23765 18680
rect 23716 18640 23722 18652
rect 23753 18649 23765 18652
rect 23799 18649 23811 18683
rect 23753 18643 23811 18649
rect 22005 18615 22063 18621
rect 22005 18612 22017 18615
rect 20496 18584 22017 18612
rect 20496 18572 20502 18584
rect 22005 18581 22017 18584
rect 22051 18581 22063 18615
rect 22005 18575 22063 18581
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 25056 18612 25084 18720
rect 25225 18717 25237 18720
rect 25271 18717 25283 18751
rect 25225 18711 25283 18717
rect 25593 18751 25651 18757
rect 25593 18717 25605 18751
rect 25639 18717 25651 18751
rect 25593 18711 25651 18717
rect 25685 18751 25743 18757
rect 25685 18717 25697 18751
rect 25731 18717 25743 18751
rect 25685 18711 25743 18717
rect 26973 18751 27031 18757
rect 26973 18717 26985 18751
rect 27019 18717 27031 18751
rect 26973 18711 27031 18717
rect 27065 18751 27123 18757
rect 27065 18717 27077 18751
rect 27111 18748 27123 18751
rect 27249 18751 27307 18757
rect 27111 18720 27200 18748
rect 27111 18717 27123 18720
rect 27065 18711 27123 18717
rect 25608 18680 25636 18711
rect 25961 18683 26019 18689
rect 25961 18680 25973 18683
rect 25608 18652 25973 18680
rect 25961 18649 25973 18652
rect 26007 18649 26019 18683
rect 25961 18643 26019 18649
rect 25777 18615 25835 18621
rect 25777 18612 25789 18615
rect 22796 18584 25789 18612
rect 22796 18572 22802 18584
rect 25777 18581 25789 18584
rect 25823 18581 25835 18615
rect 25777 18575 25835 18581
rect 25866 18572 25872 18624
rect 25924 18612 25930 18624
rect 25976 18612 26004 18643
rect 25924 18584 26004 18612
rect 26988 18612 27016 18711
rect 27172 18692 27200 18720
rect 27249 18717 27261 18751
rect 27295 18717 27307 18751
rect 27249 18711 27307 18717
rect 27341 18751 27399 18757
rect 27341 18717 27353 18751
rect 27387 18748 27399 18751
rect 27433 18751 27491 18757
rect 27433 18748 27445 18751
rect 27387 18720 27445 18748
rect 27387 18717 27399 18720
rect 27341 18711 27399 18717
rect 27433 18717 27445 18720
rect 27479 18717 27491 18751
rect 27433 18711 27491 18717
rect 28169 18751 28227 18757
rect 28169 18717 28181 18751
rect 28215 18748 28227 18751
rect 28644 18748 28672 18847
rect 28215 18720 28672 18748
rect 28215 18717 28227 18720
rect 28169 18711 28227 18717
rect 27154 18640 27160 18692
rect 27212 18640 27218 18692
rect 27264 18680 27292 18711
rect 28718 18708 28724 18760
rect 28776 18748 28782 18760
rect 28905 18751 28963 18757
rect 28905 18748 28917 18751
rect 28776 18720 28917 18748
rect 28776 18708 28782 18720
rect 28905 18717 28917 18720
rect 28951 18717 28963 18751
rect 28905 18711 28963 18717
rect 29362 18708 29368 18760
rect 29420 18748 29426 18760
rect 29549 18751 29607 18757
rect 29549 18748 29561 18751
rect 29420 18720 29561 18748
rect 29420 18708 29426 18720
rect 29549 18717 29561 18720
rect 29595 18717 29607 18751
rect 31404 18748 31432 18912
rect 31665 18819 31723 18825
rect 31665 18785 31677 18819
rect 31711 18816 31723 18819
rect 32125 18819 32183 18825
rect 32125 18816 32137 18819
rect 31711 18788 32137 18816
rect 31711 18785 31723 18788
rect 31665 18779 31723 18785
rect 32125 18785 32137 18788
rect 32171 18785 32183 18819
rect 32125 18779 32183 18785
rect 34057 18819 34115 18825
rect 34057 18785 34069 18819
rect 34103 18785 34115 18819
rect 34057 18779 34115 18785
rect 31573 18751 31631 18757
rect 31573 18748 31585 18751
rect 31404 18720 31585 18748
rect 29549 18711 29607 18717
rect 31573 18717 31585 18720
rect 31619 18717 31631 18751
rect 32033 18751 32091 18757
rect 32033 18748 32045 18751
rect 31573 18711 31631 18717
rect 31726 18720 32045 18748
rect 27522 18680 27528 18692
rect 27264 18652 27528 18680
rect 27522 18640 27528 18652
rect 27580 18680 27586 18692
rect 28629 18683 28687 18689
rect 28629 18680 28641 18683
rect 27580 18652 28641 18680
rect 27580 18640 27586 18652
rect 28629 18649 28641 18652
rect 28675 18649 28687 18683
rect 29825 18683 29883 18689
rect 29825 18680 29837 18683
rect 28629 18643 28687 18649
rect 28736 18652 29837 18680
rect 27706 18612 27712 18624
rect 26988 18584 27712 18612
rect 25924 18572 25930 18584
rect 27706 18572 27712 18584
rect 27764 18572 27770 18624
rect 28537 18615 28595 18621
rect 28537 18581 28549 18615
rect 28583 18612 28595 18615
rect 28736 18612 28764 18652
rect 29825 18649 29837 18652
rect 29871 18649 29883 18683
rect 29825 18643 29883 18649
rect 30282 18640 30288 18692
rect 30340 18640 30346 18692
rect 31478 18640 31484 18692
rect 31536 18680 31542 18692
rect 31726 18680 31754 18720
rect 32033 18717 32045 18720
rect 32079 18717 32091 18751
rect 32033 18711 32091 18717
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32493 18751 32551 18757
rect 32493 18748 32505 18751
rect 32272 18720 32505 18748
rect 32272 18708 32278 18720
rect 32493 18717 32505 18720
rect 32539 18717 32551 18751
rect 32493 18711 32551 18717
rect 31536 18652 31754 18680
rect 34072 18680 34100 18779
rect 34514 18708 34520 18760
rect 34572 18708 34578 18760
rect 34606 18680 34612 18692
rect 34072 18652 34612 18680
rect 31536 18640 31542 18652
rect 34606 18640 34612 18652
rect 34664 18640 34670 18692
rect 28583 18584 28764 18612
rect 28813 18615 28871 18621
rect 28583 18581 28595 18584
rect 28537 18575 28595 18581
rect 28813 18581 28825 18615
rect 28859 18612 28871 18615
rect 28902 18612 28908 18624
rect 28859 18584 28908 18612
rect 28859 18581 28871 18584
rect 28813 18575 28871 18581
rect 28902 18572 28908 18584
rect 28960 18572 28966 18624
rect 31938 18572 31944 18624
rect 31996 18572 32002 18624
rect 1104 18522 35236 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 35236 18522
rect 1104 18448 35236 18470
rect 4157 18411 4215 18417
rect 4157 18377 4169 18411
rect 4203 18408 4215 18411
rect 6362 18408 6368 18420
rect 4203 18380 6368 18408
rect 4203 18377 4215 18380
rect 4157 18371 4215 18377
rect 6362 18368 6368 18380
rect 6420 18368 6426 18420
rect 9401 18411 9459 18417
rect 9401 18377 9413 18411
rect 9447 18408 9459 18411
rect 9674 18408 9680 18420
rect 9447 18380 9680 18408
rect 9447 18377 9459 18380
rect 9401 18371 9459 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 10318 18368 10324 18420
rect 10376 18368 10382 18420
rect 10778 18368 10784 18420
rect 10836 18368 10842 18420
rect 11606 18368 11612 18420
rect 11664 18368 11670 18420
rect 12069 18411 12127 18417
rect 12069 18377 12081 18411
rect 12115 18408 12127 18411
rect 12434 18408 12440 18420
rect 12115 18380 12440 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 13078 18368 13084 18420
rect 13136 18408 13142 18420
rect 13906 18408 13912 18420
rect 13136 18380 13912 18408
rect 13136 18368 13142 18380
rect 13906 18368 13912 18380
rect 13964 18368 13970 18420
rect 13998 18368 14004 18420
rect 14056 18368 14062 18420
rect 14366 18368 14372 18420
rect 14424 18408 14430 18420
rect 14737 18411 14795 18417
rect 14737 18408 14749 18411
rect 14424 18380 14749 18408
rect 14424 18368 14430 18380
rect 14737 18377 14749 18380
rect 14783 18377 14795 18411
rect 14737 18371 14795 18377
rect 15102 18368 15108 18420
rect 15160 18368 15166 18420
rect 16574 18408 16580 18420
rect 15212 18380 16580 18408
rect 1578 18300 1584 18352
rect 1636 18340 1642 18352
rect 1673 18343 1731 18349
rect 1673 18340 1685 18343
rect 1636 18312 1685 18340
rect 1636 18300 1642 18312
rect 1673 18309 1685 18312
rect 1719 18309 1731 18343
rect 1673 18303 1731 18309
rect 10229 18343 10287 18349
rect 10229 18309 10241 18343
rect 10275 18340 10287 18343
rect 10336 18340 10364 18368
rect 10275 18312 10364 18340
rect 10796 18340 10824 18368
rect 10873 18343 10931 18349
rect 10873 18340 10885 18343
rect 10796 18312 10885 18340
rect 10275 18309 10287 18312
rect 10229 18303 10287 18309
rect 10873 18309 10885 18312
rect 10919 18309 10931 18343
rect 10873 18303 10931 18309
rect 11517 18343 11575 18349
rect 11517 18309 11529 18343
rect 11563 18340 11575 18343
rect 11624 18340 11652 18368
rect 12802 18340 12808 18352
rect 11563 18312 11652 18340
rect 12268 18312 12808 18340
rect 11563 18309 11575 18312
rect 11517 18303 11575 18309
rect 3329 18275 3387 18281
rect 3329 18272 3341 18275
rect 2806 18244 3341 18272
rect 3329 18241 3341 18244
rect 3375 18241 3387 18275
rect 3329 18235 3387 18241
rect 3418 18232 3424 18284
rect 3476 18232 3482 18284
rect 9033 18275 9091 18281
rect 9033 18241 9045 18275
rect 9079 18272 9091 18275
rect 9214 18272 9220 18284
rect 9079 18244 9220 18272
rect 9079 18241 9091 18244
rect 9033 18235 9091 18241
rect 9214 18232 9220 18244
rect 9272 18272 9278 18284
rect 9582 18272 9588 18284
rect 9272 18244 9588 18272
rect 9272 18232 9278 18244
rect 9582 18232 9588 18244
rect 9640 18272 9646 18284
rect 9861 18275 9919 18281
rect 9861 18272 9873 18275
rect 9640 18244 9873 18272
rect 9640 18232 9646 18244
rect 9861 18241 9873 18244
rect 9907 18241 9919 18275
rect 9861 18235 9919 18241
rect 10137 18275 10195 18281
rect 10137 18241 10149 18275
rect 10183 18272 10195 18275
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10183 18244 10977 18272
rect 10183 18241 10195 18244
rect 10137 18235 10195 18241
rect 10965 18241 10977 18244
rect 11011 18272 11023 18275
rect 11054 18272 11060 18284
rect 11011 18244 11060 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 11054 18232 11060 18244
rect 11112 18232 11118 18284
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18241 11207 18275
rect 11149 18235 11207 18241
rect 1394 18164 1400 18216
rect 1452 18164 1458 18216
rect 3436 18204 3464 18232
rect 11164 18204 11192 18235
rect 11698 18232 11704 18284
rect 11756 18232 11762 18284
rect 11790 18232 11796 18284
rect 11848 18272 11854 18284
rect 11977 18275 12035 18281
rect 11977 18272 11989 18275
rect 11848 18244 11989 18272
rect 11848 18232 11854 18244
rect 11977 18241 11989 18244
rect 12023 18241 12035 18275
rect 11977 18235 12035 18241
rect 3436 18176 3740 18204
rect 3712 18080 3740 18176
rect 9876 18176 11192 18204
rect 9876 18080 9904 18176
rect 11808 18136 11836 18232
rect 11885 18207 11943 18213
rect 11885 18173 11897 18207
rect 11931 18173 11943 18207
rect 11992 18204 12020 18235
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12268 18272 12296 18312
rect 12802 18300 12808 18312
rect 12860 18340 12866 18352
rect 13357 18343 13415 18349
rect 13357 18340 13369 18343
rect 12860 18312 13369 18340
rect 12860 18300 12866 18312
rect 13357 18309 13369 18312
rect 13403 18340 13415 18343
rect 13446 18340 13452 18352
rect 13403 18312 13452 18340
rect 13403 18309 13415 18312
rect 13357 18303 13415 18309
rect 13446 18300 13452 18312
rect 13504 18340 13510 18352
rect 14016 18340 14044 18368
rect 15212 18340 15240 18380
rect 16574 18368 16580 18380
rect 16632 18368 16638 18420
rect 18874 18408 18880 18420
rect 18708 18380 18880 18408
rect 13504 18312 13676 18340
rect 14016 18312 15240 18340
rect 13504 18300 13510 18312
rect 12124 18244 12296 18272
rect 12124 18232 12130 18244
rect 12342 18232 12348 18284
rect 12400 18232 12406 18284
rect 12529 18275 12587 18281
rect 12529 18241 12541 18275
rect 12575 18241 12587 18275
rect 12529 18235 12587 18241
rect 12621 18275 12679 18281
rect 12621 18241 12633 18275
rect 12667 18241 12679 18275
rect 12621 18235 12679 18241
rect 12250 18204 12256 18216
rect 11992 18176 12256 18204
rect 11885 18167 11943 18173
rect 11164 18108 11836 18136
rect 11900 18136 11928 18167
rect 12250 18164 12256 18176
rect 12308 18204 12314 18216
rect 12544 18204 12572 18235
rect 12308 18176 12572 18204
rect 12636 18204 12664 18235
rect 12894 18232 12900 18284
rect 12952 18232 12958 18284
rect 12986 18232 12992 18284
rect 13044 18232 13050 18284
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18241 13599 18275
rect 13648 18272 13676 18312
rect 15286 18300 15292 18352
rect 15344 18300 15350 18352
rect 15580 18312 18000 18340
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13648 18244 14013 18272
rect 13541 18235 13599 18241
rect 14001 18241 14013 18244
rect 14047 18272 14059 18275
rect 14645 18275 14703 18281
rect 14047 18244 14596 18272
rect 14047 18241 14059 18244
rect 14001 18235 14059 18241
rect 13262 18204 13268 18216
rect 12636 18176 13268 18204
rect 12308 18164 12314 18176
rect 13262 18164 13268 18176
rect 13320 18164 13326 18216
rect 13556 18204 13584 18235
rect 13722 18204 13728 18216
rect 13556 18176 13728 18204
rect 13722 18164 13728 18176
rect 13780 18164 13786 18216
rect 13817 18207 13875 18213
rect 13817 18173 13829 18207
rect 13863 18204 13875 18207
rect 13906 18204 13912 18216
rect 13863 18176 13912 18204
rect 13863 18173 13875 18176
rect 13817 18167 13875 18173
rect 13906 18164 13912 18176
rect 13964 18164 13970 18216
rect 14369 18207 14427 18213
rect 14369 18173 14381 18207
rect 14415 18204 14427 18207
rect 14458 18204 14464 18216
rect 14415 18176 14464 18204
rect 14415 18173 14427 18176
rect 14369 18167 14427 18173
rect 14458 18164 14464 18176
rect 14516 18164 14522 18216
rect 14568 18204 14596 18244
rect 14645 18241 14657 18275
rect 14691 18272 14703 18275
rect 14734 18272 14740 18284
rect 14691 18244 14740 18272
rect 14691 18241 14703 18244
rect 14645 18235 14703 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 15197 18275 15255 18281
rect 15197 18272 15209 18275
rect 14884 18244 15209 18272
rect 14884 18232 14890 18244
rect 15197 18241 15209 18244
rect 15243 18241 15255 18275
rect 15197 18235 15255 18241
rect 15470 18232 15476 18284
rect 15528 18232 15534 18284
rect 15580 18204 15608 18312
rect 17972 18284 18000 18312
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 16114 18232 16120 18284
rect 16172 18232 16178 18284
rect 17954 18232 17960 18284
rect 18012 18232 18018 18284
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 18196 18244 18613 18272
rect 18196 18232 18202 18244
rect 14568 18176 15608 18204
rect 12618 18136 12624 18148
rect 11900 18108 12624 18136
rect 11164 18080 11192 18108
rect 12618 18096 12624 18108
rect 12676 18096 12682 18148
rect 14826 18136 14832 18148
rect 13832 18108 14832 18136
rect 13832 18080 13860 18108
rect 14826 18096 14832 18108
rect 14884 18096 14890 18148
rect 15102 18096 15108 18148
rect 15160 18136 15166 18148
rect 15764 18136 15792 18232
rect 15160 18108 15792 18136
rect 15160 18096 15166 18108
rect 3142 18028 3148 18080
rect 3200 18028 3206 18080
rect 3694 18028 3700 18080
rect 3752 18028 3758 18080
rect 9769 18071 9827 18077
rect 9769 18037 9781 18071
rect 9815 18068 9827 18071
rect 9858 18068 9864 18080
rect 9815 18040 9864 18068
rect 9815 18037 9827 18040
rect 9769 18031 9827 18037
rect 9858 18028 9864 18040
rect 9916 18028 9922 18080
rect 10689 18071 10747 18077
rect 10689 18037 10701 18071
rect 10735 18068 10747 18071
rect 11146 18068 11152 18080
rect 10735 18040 11152 18068
rect 10735 18037 10747 18040
rect 10689 18031 10747 18037
rect 11146 18028 11152 18040
rect 11204 18028 11210 18080
rect 12434 18028 12440 18080
rect 12492 18028 12498 18080
rect 12710 18028 12716 18080
rect 12768 18028 12774 18080
rect 13170 18028 13176 18080
rect 13228 18028 13234 18080
rect 13725 18071 13783 18077
rect 13725 18037 13737 18071
rect 13771 18068 13783 18071
rect 13814 18068 13820 18080
rect 13771 18040 13820 18068
rect 13771 18037 13783 18040
rect 13725 18031 13783 18037
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14185 18071 14243 18077
rect 14185 18037 14197 18071
rect 14231 18068 14243 18071
rect 14461 18071 14519 18077
rect 14461 18068 14473 18071
rect 14231 18040 14473 18068
rect 14231 18037 14243 18040
rect 14185 18031 14243 18037
rect 14461 18037 14473 18040
rect 14507 18068 14519 18071
rect 15856 18068 15884 18232
rect 14507 18040 15884 18068
rect 16945 18071 17003 18077
rect 14507 18037 14519 18040
rect 14461 18031 14519 18037
rect 16945 18037 16957 18071
rect 16991 18068 17003 18071
rect 17034 18068 17040 18080
rect 16991 18040 17040 18068
rect 16991 18037 17003 18040
rect 16945 18031 17003 18037
rect 17034 18028 17040 18040
rect 17092 18068 17098 18080
rect 17862 18068 17868 18080
rect 17092 18040 17868 18068
rect 17092 18028 17098 18040
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 18340 18068 18368 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18708 18204 18736 18380
rect 18874 18368 18880 18380
rect 18932 18368 18938 18420
rect 18966 18368 18972 18420
rect 19024 18408 19030 18420
rect 19061 18411 19119 18417
rect 19061 18408 19073 18411
rect 19024 18380 19073 18408
rect 19024 18368 19030 18380
rect 19061 18377 19073 18380
rect 19107 18377 19119 18411
rect 19061 18371 19119 18377
rect 19429 18411 19487 18417
rect 19429 18377 19441 18411
rect 19475 18408 19487 18411
rect 19797 18411 19855 18417
rect 19475 18380 19564 18408
rect 19475 18377 19487 18380
rect 19429 18371 19487 18377
rect 19536 18349 19564 18380
rect 19797 18377 19809 18411
rect 19843 18408 19855 18411
rect 22738 18408 22744 18420
rect 19843 18380 22744 18408
rect 19843 18377 19855 18380
rect 19797 18371 19855 18377
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 22830 18368 22836 18420
rect 22888 18368 22894 18420
rect 30098 18368 30104 18420
rect 30156 18368 30162 18420
rect 30282 18368 30288 18420
rect 30340 18368 30346 18420
rect 31938 18368 31944 18420
rect 31996 18368 32002 18420
rect 34514 18368 34520 18420
rect 34572 18368 34578 18420
rect 18785 18343 18843 18349
rect 18785 18309 18797 18343
rect 18831 18340 18843 18343
rect 19521 18343 19579 18349
rect 18831 18312 19472 18340
rect 18831 18309 18843 18312
rect 18785 18303 18843 18309
rect 18874 18232 18880 18284
rect 18932 18232 18938 18284
rect 18984 18281 19012 18312
rect 19444 18284 19472 18312
rect 19521 18309 19533 18343
rect 19567 18340 19579 18343
rect 20070 18340 20076 18352
rect 19567 18312 20076 18340
rect 19567 18309 19579 18312
rect 19521 18303 19579 18309
rect 20070 18300 20076 18312
rect 20128 18300 20134 18352
rect 18969 18275 19027 18281
rect 18969 18241 18981 18275
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19242 18272 19248 18284
rect 19116 18244 19248 18272
rect 19116 18232 19122 18244
rect 19242 18232 19248 18244
rect 19300 18232 19306 18284
rect 19426 18232 19432 18284
rect 19484 18232 19490 18284
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18241 19763 18275
rect 19705 18235 19763 18241
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18241 19855 18275
rect 22741 18275 22799 18281
rect 22741 18272 22753 18275
rect 19797 18235 19855 18241
rect 22204 18244 22753 18272
rect 19720 18204 19748 18235
rect 18708 18176 19748 18204
rect 18414 18096 18420 18148
rect 18472 18136 18478 18148
rect 19812 18136 19840 18235
rect 18472 18108 19840 18136
rect 18472 18096 18478 18108
rect 19058 18068 19064 18080
rect 18340 18040 19064 18068
rect 19058 18028 19064 18040
rect 19116 18028 19122 18080
rect 19150 18028 19156 18080
rect 19208 18068 19214 18080
rect 21358 18068 21364 18080
rect 19208 18040 21364 18068
rect 19208 18028 19214 18040
rect 21358 18028 21364 18040
rect 21416 18068 21422 18080
rect 22204 18068 22232 18244
rect 22741 18241 22753 18244
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18272 22983 18275
rect 23198 18272 23204 18284
rect 22971 18244 23204 18272
rect 22971 18241 22983 18244
rect 22925 18235 22983 18241
rect 22281 18207 22339 18213
rect 22281 18173 22293 18207
rect 22327 18204 22339 18207
rect 22554 18204 22560 18216
rect 22327 18176 22560 18204
rect 22327 18173 22339 18176
rect 22281 18167 22339 18173
rect 22554 18164 22560 18176
rect 22612 18164 22618 18216
rect 22646 18164 22652 18216
rect 22704 18204 22710 18216
rect 22940 18204 22968 18235
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 27154 18232 27160 18284
rect 27212 18272 27218 18284
rect 27890 18272 27896 18284
rect 27212 18244 27896 18272
rect 27212 18232 27218 18244
rect 27890 18232 27896 18244
rect 27948 18232 27954 18284
rect 30116 18272 30144 18368
rect 31956 18340 31984 18368
rect 33045 18343 33103 18349
rect 33045 18340 33057 18343
rect 31956 18312 33057 18340
rect 33045 18309 33057 18312
rect 33091 18309 33103 18343
rect 33045 18303 33103 18309
rect 33778 18300 33784 18352
rect 33836 18300 33842 18352
rect 30193 18275 30251 18281
rect 30193 18272 30205 18275
rect 30116 18244 30205 18272
rect 30193 18241 30205 18244
rect 30239 18241 30251 18275
rect 30193 18235 30251 18241
rect 22704 18176 22968 18204
rect 32769 18207 32827 18213
rect 22704 18164 22710 18176
rect 32769 18173 32781 18207
rect 32815 18173 32827 18207
rect 32769 18167 32827 18173
rect 32784 18080 32812 18167
rect 22557 18071 22615 18077
rect 22557 18068 22569 18071
rect 21416 18040 22569 18068
rect 21416 18028 21422 18040
rect 22557 18037 22569 18040
rect 22603 18037 22615 18071
rect 22557 18031 22615 18037
rect 32677 18071 32735 18077
rect 32677 18037 32689 18071
rect 32723 18068 32735 18071
rect 32766 18068 32772 18080
rect 32723 18040 32772 18068
rect 32723 18037 32735 18040
rect 32677 18031 32735 18037
rect 32766 18028 32772 18040
rect 32824 18028 32830 18080
rect 1104 17978 35248 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 35248 17978
rect 1104 17904 35248 17926
rect 4062 17824 4068 17876
rect 4120 17824 4126 17876
rect 4341 17867 4399 17873
rect 4341 17833 4353 17867
rect 4387 17864 4399 17867
rect 4706 17864 4712 17876
rect 4387 17836 4712 17864
rect 4387 17833 4399 17836
rect 4341 17827 4399 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 9732 17836 10609 17864
rect 9732 17824 9738 17836
rect 10597 17833 10609 17836
rect 10643 17833 10655 17867
rect 10597 17827 10655 17833
rect 11057 17867 11115 17873
rect 11057 17833 11069 17867
rect 11103 17864 11115 17867
rect 11146 17864 11152 17876
rect 11103 17836 11152 17864
rect 11103 17833 11115 17836
rect 11057 17827 11115 17833
rect 11146 17824 11152 17836
rect 11204 17824 11210 17876
rect 11977 17867 12035 17873
rect 11977 17833 11989 17867
rect 12023 17864 12035 17867
rect 12710 17864 12716 17876
rect 12023 17836 12716 17864
rect 12023 17833 12035 17836
rect 11977 17827 12035 17833
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 12894 17824 12900 17876
rect 12952 17824 12958 17876
rect 12986 17824 12992 17876
rect 13044 17864 13050 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 13044 17836 13277 17864
rect 13044 17824 13050 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 14366 17824 14372 17876
rect 14424 17864 14430 17876
rect 15013 17867 15071 17873
rect 15013 17864 15025 17867
rect 14424 17836 15025 17864
rect 14424 17824 14430 17836
rect 15013 17833 15025 17836
rect 15059 17833 15071 17867
rect 15013 17827 15071 17833
rect 15102 17824 15108 17876
rect 15160 17824 15166 17876
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19613 17867 19671 17873
rect 19613 17864 19625 17867
rect 19484 17836 19625 17864
rect 19484 17824 19490 17836
rect 19613 17833 19625 17836
rect 19659 17833 19671 17867
rect 19613 17827 19671 17833
rect 20714 17824 20720 17876
rect 20772 17824 20778 17876
rect 27341 17867 27399 17873
rect 22204 17836 24808 17864
rect 11514 17756 11520 17808
rect 11572 17756 11578 17808
rect 11609 17799 11667 17805
rect 11609 17765 11621 17799
rect 11655 17796 11667 17799
rect 11885 17799 11943 17805
rect 11885 17796 11897 17799
rect 11655 17768 11897 17796
rect 11655 17765 11667 17768
rect 11609 17759 11667 17765
rect 11885 17765 11897 17768
rect 11931 17796 11943 17799
rect 12526 17796 12532 17808
rect 11931 17768 12532 17796
rect 11931 17765 11943 17768
rect 11885 17759 11943 17765
rect 12526 17756 12532 17768
rect 12584 17756 12590 17808
rect 12912 17796 12940 17824
rect 13173 17799 13231 17805
rect 13173 17796 13185 17799
rect 12912 17768 13185 17796
rect 13173 17765 13185 17768
rect 13219 17765 13231 17799
rect 13173 17759 13231 17765
rect 14734 17756 14740 17808
rect 14792 17796 14798 17808
rect 15120 17796 15148 17824
rect 20898 17796 20904 17808
rect 14792 17768 15148 17796
rect 20180 17768 20904 17796
rect 14792 17756 14798 17768
rect 3602 17688 3608 17740
rect 3660 17728 3666 17740
rect 3973 17731 4031 17737
rect 3973 17728 3985 17731
rect 3660 17700 3985 17728
rect 3660 17688 3666 17700
rect 3973 17697 3985 17700
rect 4019 17697 4031 17731
rect 3973 17691 4031 17697
rect 5166 17688 5172 17740
rect 5224 17728 5230 17740
rect 5445 17731 5503 17737
rect 5445 17728 5457 17731
rect 5224 17700 5457 17728
rect 5224 17688 5230 17700
rect 5445 17697 5457 17700
rect 5491 17697 5503 17731
rect 5445 17691 5503 17697
rect 5721 17731 5779 17737
rect 5721 17697 5733 17731
rect 5767 17728 5779 17731
rect 5767 17700 6316 17728
rect 5767 17697 5779 17700
rect 5721 17691 5779 17697
rect 934 17620 940 17672
rect 992 17660 998 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 992 17632 1409 17660
rect 992 17620 998 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 3142 17620 3148 17672
rect 3200 17660 3206 17672
rect 3878 17660 3884 17672
rect 3200 17632 3884 17660
rect 3200 17620 3206 17632
rect 3878 17620 3884 17632
rect 3936 17620 3942 17672
rect 4157 17663 4215 17669
rect 4157 17629 4169 17663
rect 4203 17629 4215 17663
rect 4157 17623 4215 17629
rect 4172 17592 4200 17623
rect 4614 17620 4620 17672
rect 4672 17660 4678 17672
rect 5258 17660 5264 17672
rect 4672 17632 5264 17660
rect 4672 17620 4678 17632
rect 5258 17620 5264 17632
rect 5316 17660 5322 17672
rect 5353 17663 5411 17669
rect 5353 17660 5365 17663
rect 5316 17632 5365 17660
rect 5316 17620 5322 17632
rect 5353 17629 5365 17632
rect 5399 17629 5411 17663
rect 5353 17623 5411 17629
rect 6086 17620 6092 17672
rect 6144 17660 6150 17672
rect 6288 17669 6316 17700
rect 12066 17688 12072 17740
rect 12124 17688 12130 17740
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 12894 17728 12900 17740
rect 12492 17700 12900 17728
rect 12492 17688 12498 17700
rect 12894 17688 12900 17700
rect 12952 17728 12958 17740
rect 20180 17737 20208 17768
rect 20898 17756 20904 17768
rect 20956 17756 20962 17808
rect 20165 17731 20223 17737
rect 20165 17728 20177 17731
rect 12952 17700 13768 17728
rect 12952 17688 12958 17700
rect 6181 17663 6239 17669
rect 6181 17660 6193 17663
rect 6144 17632 6193 17660
rect 6144 17620 6150 17632
rect 6181 17629 6193 17632
rect 6227 17629 6239 17663
rect 6181 17623 6239 17629
rect 6273 17663 6331 17669
rect 6273 17629 6285 17663
rect 6319 17629 6331 17663
rect 6273 17623 6331 17629
rect 3988 17564 4200 17592
rect 6196 17592 6224 17623
rect 11054 17620 11060 17672
rect 11112 17660 11118 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11112 17632 11805 17660
rect 11112 17620 11118 17632
rect 11793 17629 11805 17632
rect 11839 17660 11851 17663
rect 12342 17660 12348 17672
rect 11839 17632 12348 17660
rect 11839 17629 11851 17632
rect 11793 17623 11851 17629
rect 12342 17620 12348 17632
rect 12400 17620 12406 17672
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12618 17660 12624 17672
rect 12575 17632 12624 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 13004 17669 13032 17700
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 12713 17623 12771 17629
rect 12989 17663 13047 17669
rect 12989 17629 13001 17663
rect 13035 17629 13047 17663
rect 12989 17623 13047 17629
rect 9953 17595 10011 17601
rect 6196 17564 6776 17592
rect 3988 17536 4016 17564
rect 6748 17536 6776 17564
rect 9953 17561 9965 17595
rect 9999 17592 10011 17595
rect 11149 17595 11207 17601
rect 9999 17564 10916 17592
rect 9999 17561 10011 17564
rect 9953 17555 10011 17561
rect 10888 17536 10916 17564
rect 11149 17561 11161 17595
rect 11195 17561 11207 17595
rect 11149 17555 11207 17561
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17524 1639 17527
rect 1670 17524 1676 17536
rect 1627 17496 1676 17524
rect 1627 17493 1639 17496
rect 1581 17487 1639 17493
rect 1670 17484 1676 17496
rect 1728 17484 1734 17536
rect 3970 17484 3976 17536
rect 4028 17484 4034 17536
rect 6454 17484 6460 17536
rect 6512 17484 6518 17536
rect 6730 17484 6736 17536
rect 6788 17484 6794 17536
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 9309 17527 9367 17533
rect 9309 17524 9321 17527
rect 9272 17496 9321 17524
rect 9272 17484 9278 17496
rect 9309 17493 9321 17496
rect 9355 17493 9367 17527
rect 9309 17487 9367 17493
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 10229 17527 10287 17533
rect 10229 17524 10241 17527
rect 9916 17496 10241 17524
rect 9916 17484 9922 17496
rect 10229 17493 10241 17496
rect 10275 17493 10287 17527
rect 10229 17487 10287 17493
rect 10870 17484 10876 17536
rect 10928 17524 10934 17536
rect 11164 17524 11192 17555
rect 11974 17552 11980 17604
rect 12032 17592 12038 17604
rect 12728 17592 12756 17623
rect 13538 17620 13544 17672
rect 13596 17620 13602 17672
rect 13630 17620 13636 17672
rect 13688 17620 13694 17672
rect 13740 17669 13768 17700
rect 19996 17700 20177 17728
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 13909 17663 13967 17669
rect 13909 17660 13921 17663
rect 13872 17632 13921 17660
rect 13872 17620 13878 17632
rect 13909 17629 13921 17632
rect 13955 17629 13967 17663
rect 13909 17623 13967 17629
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 16853 17663 16911 17669
rect 16853 17629 16865 17663
rect 16899 17629 16911 17663
rect 16853 17623 16911 17629
rect 12032 17564 12756 17592
rect 12032 17552 12038 17564
rect 12434 17524 12440 17536
rect 10928 17496 12440 17524
rect 10928 17484 10934 17496
rect 12434 17484 12440 17496
rect 12492 17524 12498 17536
rect 13722 17524 13728 17536
rect 12492 17496 13728 17524
rect 12492 17484 12498 17496
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16868 17524 16896 17623
rect 19334 17620 19340 17672
rect 19392 17660 19398 17672
rect 19996 17669 20024 17700
rect 20165 17697 20177 17700
rect 20211 17697 20223 17731
rect 21082 17728 21088 17740
rect 20165 17691 20223 17697
rect 20456 17700 21088 17728
rect 20456 17669 20484 17700
rect 21082 17688 21088 17700
rect 21140 17688 21146 17740
rect 19797 17663 19855 17669
rect 19797 17660 19809 17663
rect 19392 17632 19809 17660
rect 19392 17620 19398 17632
rect 19797 17629 19809 17632
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17629 20499 17663
rect 20441 17623 20499 17629
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 19812 17592 19840 17623
rect 20070 17592 20076 17604
rect 19812 17564 20076 17592
rect 20070 17552 20076 17564
rect 20128 17552 20134 17604
rect 20548 17592 20576 17623
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 20993 17663 21051 17669
rect 20993 17660 21005 17663
rect 20956 17632 21005 17660
rect 20956 17620 20962 17632
rect 20993 17629 21005 17632
rect 21039 17629 21051 17663
rect 20993 17623 21051 17629
rect 21174 17620 21180 17672
rect 21232 17620 21238 17672
rect 21450 17620 21456 17672
rect 21508 17620 21514 17672
rect 22204 17669 22232 17836
rect 23014 17756 23020 17808
rect 23072 17756 23078 17808
rect 22557 17731 22615 17737
rect 22557 17728 22569 17731
rect 22388 17700 22569 17728
rect 22189 17663 22247 17669
rect 22189 17629 22201 17663
rect 22235 17629 22247 17663
rect 22189 17623 22247 17629
rect 21266 17592 21272 17604
rect 20548 17564 21272 17592
rect 21266 17552 21272 17564
rect 21324 17592 21330 17604
rect 22388 17592 22416 17700
rect 22557 17697 22569 17700
rect 22603 17728 22615 17731
rect 23201 17731 23259 17737
rect 22603 17700 23152 17728
rect 22603 17697 22615 17700
rect 22557 17691 22615 17697
rect 22465 17663 22523 17669
rect 22465 17629 22477 17663
rect 22511 17660 22523 17663
rect 22649 17663 22707 17669
rect 22511 17632 22600 17660
rect 22511 17629 22523 17632
rect 22465 17623 22523 17629
rect 21324 17564 22416 17592
rect 21324 17552 21330 17564
rect 22572 17536 22600 17632
rect 22649 17629 22661 17663
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 22664 17592 22692 17623
rect 22738 17620 22744 17672
rect 22796 17620 22802 17672
rect 23124 17669 23152 17700
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 24581 17731 24639 17737
rect 24581 17728 24593 17731
rect 23247 17700 24593 17728
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 24581 17697 24593 17700
rect 24627 17697 24639 17731
rect 24780 17728 24808 17836
rect 27341 17833 27353 17867
rect 27387 17864 27399 17867
rect 27522 17864 27528 17876
rect 27387 17836 27528 17864
rect 27387 17833 27399 17836
rect 27341 17827 27399 17833
rect 27522 17824 27528 17836
rect 27580 17824 27586 17876
rect 27706 17824 27712 17876
rect 27764 17864 27770 17876
rect 28261 17867 28319 17873
rect 28261 17864 28273 17867
rect 27764 17836 28273 17864
rect 27764 17824 27770 17836
rect 28261 17833 28273 17836
rect 28307 17833 28319 17867
rect 28261 17827 28319 17833
rect 27356 17768 28028 17796
rect 27356 17728 27384 17768
rect 24780 17700 27384 17728
rect 24581 17691 24639 17697
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17629 23167 17663
rect 23109 17623 23167 17629
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23474 17620 23480 17672
rect 23532 17660 23538 17672
rect 23569 17663 23627 17669
rect 23569 17660 23581 17663
rect 23532 17632 23581 17660
rect 23532 17620 23538 17632
rect 23569 17629 23581 17632
rect 23615 17629 23627 17663
rect 23569 17623 23627 17629
rect 23750 17620 23756 17672
rect 23808 17620 23814 17672
rect 24673 17663 24731 17669
rect 24673 17629 24685 17663
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 23017 17595 23075 17601
rect 22664 17564 22876 17592
rect 16172 17496 16896 17524
rect 17589 17527 17647 17533
rect 16172 17484 16178 17496
rect 17589 17493 17601 17527
rect 17635 17524 17647 17527
rect 20714 17524 20720 17536
rect 17635 17496 20720 17524
rect 17635 17493 17647 17496
rect 17589 17487 17647 17493
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 20806 17484 20812 17536
rect 20864 17484 20870 17536
rect 22554 17484 22560 17536
rect 22612 17524 22618 17536
rect 22738 17524 22744 17536
rect 22612 17496 22744 17524
rect 22612 17484 22618 17496
rect 22738 17484 22744 17496
rect 22796 17484 22802 17536
rect 22848 17533 22876 17564
rect 23017 17561 23029 17595
rect 23063 17592 23075 17595
rect 23658 17592 23664 17604
rect 23063 17564 23664 17592
rect 23063 17561 23075 17564
rect 23017 17555 23075 17561
rect 23658 17552 23664 17564
rect 23716 17592 23722 17604
rect 24688 17592 24716 17623
rect 27356 17601 27384 17700
rect 27632 17700 27844 17728
rect 27522 17620 27528 17672
rect 27580 17660 27586 17672
rect 27632 17669 27660 17700
rect 27816 17669 27844 17700
rect 28000 17669 28028 17768
rect 28276 17728 28304 17827
rect 33778 17824 33784 17876
rect 33836 17824 33842 17876
rect 28810 17756 28816 17808
rect 28868 17756 28874 17808
rect 28718 17728 28724 17740
rect 28276 17700 28724 17728
rect 28644 17669 28672 17700
rect 28718 17688 28724 17700
rect 28776 17688 28782 17740
rect 27617 17663 27675 17669
rect 27617 17660 27629 17663
rect 27580 17632 27629 17660
rect 27580 17620 27586 17632
rect 27617 17629 27629 17632
rect 27663 17629 27675 17663
rect 27617 17623 27675 17629
rect 27709 17663 27767 17669
rect 27709 17629 27721 17663
rect 27755 17629 27767 17663
rect 27709 17623 27767 17629
rect 27801 17663 27859 17669
rect 27801 17629 27813 17663
rect 27847 17629 27859 17663
rect 27801 17623 27859 17629
rect 27985 17663 28043 17669
rect 27985 17629 27997 17663
rect 28031 17629 28043 17663
rect 28537 17663 28595 17669
rect 28537 17660 28549 17663
rect 27985 17623 28043 17629
rect 28276 17632 28549 17660
rect 23716 17564 24716 17592
rect 27341 17595 27399 17601
rect 23716 17552 23722 17564
rect 27341 17561 27353 17595
rect 27387 17592 27399 17595
rect 27430 17592 27436 17604
rect 27387 17564 27436 17592
rect 27387 17561 27399 17564
rect 27341 17555 27399 17561
rect 27430 17552 27436 17564
rect 27488 17552 27494 17604
rect 27724 17592 27752 17623
rect 27632 17564 27752 17592
rect 27632 17536 27660 17564
rect 27890 17552 27896 17604
rect 27948 17592 27954 17604
rect 28077 17595 28135 17601
rect 28077 17592 28089 17595
rect 27948 17564 28089 17592
rect 27948 17552 27954 17564
rect 28077 17561 28089 17564
rect 28123 17592 28135 17595
rect 28166 17592 28172 17604
rect 28123 17564 28172 17592
rect 28123 17561 28135 17564
rect 28077 17555 28135 17561
rect 28166 17552 28172 17564
rect 28224 17552 28230 17604
rect 22833 17527 22891 17533
rect 22833 17493 22845 17527
rect 22879 17524 22891 17527
rect 23106 17524 23112 17536
rect 22879 17496 23112 17524
rect 22879 17493 22891 17496
rect 22833 17487 22891 17493
rect 23106 17484 23112 17496
rect 23164 17524 23170 17536
rect 23385 17527 23443 17533
rect 23385 17524 23397 17527
rect 23164 17496 23397 17524
rect 23164 17484 23170 17496
rect 23385 17493 23397 17496
rect 23431 17493 23443 17527
rect 23385 17487 23443 17493
rect 25501 17527 25559 17533
rect 25501 17493 25513 17527
rect 25547 17524 25559 17527
rect 26970 17524 26976 17536
rect 25547 17496 26976 17524
rect 25547 17493 25559 17496
rect 25501 17487 25559 17493
rect 26970 17484 26976 17496
rect 27028 17484 27034 17536
rect 27525 17527 27583 17533
rect 27525 17493 27537 17527
rect 27571 17524 27583 17527
rect 27614 17524 27620 17536
rect 27571 17496 27620 17524
rect 27571 17493 27583 17496
rect 27525 17487 27583 17493
rect 27614 17484 27620 17496
rect 27672 17484 27678 17536
rect 27798 17484 27804 17536
rect 27856 17524 27862 17536
rect 28276 17533 28304 17632
rect 28537 17629 28549 17632
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 28629 17663 28687 17669
rect 28629 17629 28641 17663
rect 28675 17629 28687 17663
rect 33689 17663 33747 17669
rect 33689 17660 33701 17663
rect 28629 17623 28687 17629
rect 33612 17632 33701 17660
rect 28813 17595 28871 17601
rect 28813 17561 28825 17595
rect 28859 17592 28871 17595
rect 28902 17592 28908 17604
rect 28859 17564 28908 17592
rect 28859 17561 28871 17564
rect 28813 17555 28871 17561
rect 28276 17527 28335 17533
rect 28276 17524 28289 17527
rect 27856 17496 28289 17524
rect 27856 17484 27862 17496
rect 28277 17493 28289 17496
rect 28323 17493 28335 17527
rect 28277 17487 28335 17493
rect 28442 17484 28448 17536
rect 28500 17484 28506 17536
rect 28534 17484 28540 17536
rect 28592 17524 28598 17536
rect 28828 17524 28856 17555
rect 28902 17552 28908 17564
rect 28960 17552 28966 17604
rect 33612 17536 33640 17632
rect 33689 17629 33701 17632
rect 33735 17629 33747 17663
rect 33689 17623 33747 17629
rect 28592 17496 28856 17524
rect 28592 17484 28598 17496
rect 33594 17484 33600 17536
rect 33652 17484 33658 17536
rect 1104 17434 35236 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 35236 17434
rect 1104 17360 35236 17382
rect 3234 17280 3240 17332
rect 3292 17320 3298 17332
rect 3513 17323 3571 17329
rect 3513 17320 3525 17323
rect 3292 17292 3525 17320
rect 3292 17280 3298 17292
rect 3513 17289 3525 17292
rect 3559 17289 3571 17323
rect 3513 17283 3571 17289
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 22922 17320 22928 17332
rect 6512 17292 22928 17320
rect 6512 17280 6518 17292
rect 22922 17280 22928 17292
rect 22980 17280 22986 17332
rect 23014 17280 23020 17332
rect 23072 17280 23078 17332
rect 23106 17280 23112 17332
rect 23164 17280 23170 17332
rect 23290 17280 23296 17332
rect 23348 17320 23354 17332
rect 23477 17323 23535 17329
rect 23477 17320 23489 17323
rect 23348 17292 23489 17320
rect 23348 17280 23354 17292
rect 23477 17289 23489 17292
rect 23523 17289 23535 17323
rect 23477 17283 23535 17289
rect 25685 17323 25743 17329
rect 25685 17289 25697 17323
rect 25731 17320 25743 17323
rect 25866 17320 25872 17332
rect 25731 17292 25872 17320
rect 25731 17289 25743 17292
rect 25685 17283 25743 17289
rect 25866 17280 25872 17292
rect 25924 17280 25930 17332
rect 27614 17280 27620 17332
rect 27672 17280 27678 17332
rect 27798 17280 27804 17332
rect 27856 17280 27862 17332
rect 28442 17280 28448 17332
rect 28500 17280 28506 17332
rect 28810 17280 28816 17332
rect 28868 17280 28874 17332
rect 29273 17323 29331 17329
rect 29273 17289 29285 17323
rect 29319 17320 29331 17323
rect 29362 17320 29368 17332
rect 29319 17292 29368 17320
rect 29319 17289 29331 17292
rect 29273 17283 29331 17289
rect 29362 17280 29368 17292
rect 29420 17280 29426 17332
rect 31478 17280 31484 17332
rect 31536 17280 31542 17332
rect 6825 17255 6883 17261
rect 3620 17224 5028 17252
rect 3620 17196 3648 17224
rect 3602 17144 3608 17196
rect 3660 17144 3666 17196
rect 3878 17144 3884 17196
rect 3936 17144 3942 17196
rect 5000 17193 5028 17224
rect 6825 17221 6837 17255
rect 6871 17252 6883 17255
rect 7558 17252 7564 17264
rect 6871 17224 7564 17252
rect 6871 17221 6883 17224
rect 6825 17215 6883 17221
rect 4985 17187 5043 17193
rect 4985 17153 4997 17187
rect 5031 17153 5043 17187
rect 4985 17147 5043 17153
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 6932 17193 6960 17224
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 8694 17224 9137 17252
rect 9125 17221 9137 17224
rect 9171 17221 9183 17255
rect 9125 17215 9183 17221
rect 10137 17255 10195 17261
rect 10137 17221 10149 17255
rect 10183 17252 10195 17255
rect 10870 17252 10876 17264
rect 10183 17224 10876 17252
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 10870 17212 10876 17224
rect 10928 17212 10934 17264
rect 12176 17224 12756 17252
rect 6917 17187 6975 17193
rect 6917 17153 6929 17187
rect 6963 17153 6975 17187
rect 9214 17184 9220 17196
rect 6917 17147 6975 17153
rect 8772 17156 9220 17184
rect 3786 17076 3792 17128
rect 3844 17076 3850 17128
rect 5074 17076 5080 17128
rect 5132 17076 5138 17128
rect 6380 17116 6408 17144
rect 8772 17128 8800 17156
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9309 17187 9367 17193
rect 9309 17153 9321 17187
rect 9355 17153 9367 17187
rect 9309 17147 9367 17153
rect 6822 17116 6828 17128
rect 6380 17088 6828 17116
rect 6822 17076 6828 17088
rect 6880 17116 6886 17128
rect 7193 17119 7251 17125
rect 7193 17116 7205 17119
rect 6880 17088 7205 17116
rect 6880 17076 6886 17088
rect 7193 17085 7205 17088
rect 7239 17085 7251 17119
rect 7469 17119 7527 17125
rect 7469 17116 7481 17119
rect 7193 17079 7251 17085
rect 7300 17088 7481 17116
rect 5353 17051 5411 17057
rect 5353 17017 5365 17051
rect 5399 17048 5411 17051
rect 7300 17048 7328 17088
rect 7469 17085 7481 17088
rect 7515 17085 7527 17119
rect 7469 17079 7527 17085
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 8754 17116 8760 17128
rect 7616 17088 8760 17116
rect 7616 17076 7622 17088
rect 8754 17076 8760 17088
rect 8812 17076 8818 17128
rect 8941 17119 8999 17125
rect 8941 17085 8953 17119
rect 8987 17116 8999 17119
rect 9324 17116 9352 17147
rect 11514 17144 11520 17196
rect 11572 17184 11578 17196
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11572 17156 11989 17184
rect 11572 17144 11578 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 8987 17088 9352 17116
rect 8987 17085 8999 17088
rect 8941 17079 8999 17085
rect 5399 17020 7328 17048
rect 5399 17017 5411 17020
rect 5353 17011 5411 17017
rect 11974 17008 11980 17060
rect 12032 17048 12038 17060
rect 12176 17057 12204 17224
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 12268 17116 12296 17147
rect 12342 17144 12348 17196
rect 12400 17184 12406 17196
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12400 17156 12633 17184
rect 12400 17144 12406 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12728 17184 12756 17224
rect 13262 17212 13268 17264
rect 13320 17212 13326 17264
rect 13538 17212 13544 17264
rect 13596 17212 13602 17264
rect 16574 17212 16580 17264
rect 16632 17212 16638 17264
rect 18322 17212 18328 17264
rect 18380 17212 18386 17264
rect 20806 17212 20812 17264
rect 20864 17212 20870 17264
rect 21082 17212 21088 17264
rect 21140 17212 21146 17264
rect 21266 17212 21272 17264
rect 21324 17212 21330 17264
rect 21450 17212 21456 17264
rect 21508 17212 21514 17264
rect 12784 17187 12842 17193
rect 12784 17184 12796 17187
rect 12728 17156 12796 17184
rect 12621 17147 12679 17153
rect 12784 17153 12796 17156
rect 12830 17153 12842 17187
rect 12784 17147 12842 17153
rect 12434 17116 12440 17128
rect 12268 17088 12440 17116
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 12636 17116 12664 17147
rect 12894 17144 12900 17196
rect 12952 17144 12958 17196
rect 12986 17144 12992 17196
rect 13044 17184 13050 17196
rect 13556 17184 13584 17212
rect 13044 17156 13584 17184
rect 15841 17187 15899 17193
rect 13044 17144 13050 17156
rect 15841 17153 15853 17187
rect 15887 17184 15899 17187
rect 15930 17184 15936 17196
rect 15887 17156 15936 17184
rect 15887 17153 15899 17156
rect 15841 17147 15899 17153
rect 15930 17144 15936 17156
rect 15988 17184 15994 17196
rect 16301 17187 16359 17193
rect 16301 17184 16313 17187
rect 15988 17156 16313 17184
rect 15988 17144 15994 17156
rect 16301 17153 16313 17156
rect 16347 17153 16359 17187
rect 16301 17147 16359 17153
rect 16485 17187 16543 17193
rect 16485 17153 16497 17187
rect 16531 17153 16543 17187
rect 16485 17147 16543 17153
rect 13906 17116 13912 17128
rect 12636 17088 13912 17116
rect 13906 17076 13912 17088
rect 13964 17076 13970 17128
rect 15746 17076 15752 17128
rect 15804 17116 15810 17128
rect 16500 17116 16528 17147
rect 15804 17088 16528 17116
rect 15804 17076 15810 17088
rect 12161 17051 12219 17057
rect 12161 17048 12173 17051
rect 12032 17020 12173 17048
rect 12032 17008 12038 17020
rect 12161 17017 12173 17020
rect 12207 17017 12219 17051
rect 12161 17011 12219 17017
rect 16209 17051 16267 17057
rect 16209 17017 16221 17051
rect 16255 17048 16267 17051
rect 16592 17048 16620 17212
rect 17954 17144 17960 17196
rect 18012 17184 18018 17196
rect 18012 17156 18920 17184
rect 18012 17144 18018 17156
rect 18230 17076 18236 17128
rect 18288 17076 18294 17128
rect 18325 17119 18383 17125
rect 18325 17085 18337 17119
rect 18371 17085 18383 17119
rect 18325 17079 18383 17085
rect 16255 17020 16620 17048
rect 16255 17017 16267 17020
rect 16209 17011 16267 17017
rect 17402 17008 17408 17060
rect 17460 17048 17466 17060
rect 18340 17048 18368 17079
rect 17460 17020 18368 17048
rect 18785 17051 18843 17057
rect 17460 17008 17466 17020
rect 18785 17017 18797 17051
rect 18831 17017 18843 17051
rect 18892 17048 18920 17156
rect 20070 17144 20076 17196
rect 20128 17184 20134 17196
rect 20441 17187 20499 17193
rect 20441 17184 20453 17187
rect 20128 17156 20453 17184
rect 20128 17144 20134 17156
rect 20441 17153 20453 17156
rect 20487 17153 20499 17187
rect 20441 17147 20499 17153
rect 20533 17119 20591 17125
rect 20533 17085 20545 17119
rect 20579 17116 20591 17119
rect 20824 17116 20852 17212
rect 21100 17184 21128 17212
rect 23032 17184 23060 17280
rect 23124 17193 23152 17280
rect 27433 17255 27491 17261
rect 27433 17221 27445 17255
rect 27479 17252 27491 17255
rect 27632 17252 27660 17280
rect 27479 17224 27844 17252
rect 27479 17221 27491 17224
rect 27433 17215 27491 17221
rect 27816 17196 27844 17224
rect 21100 17156 23060 17184
rect 23109 17187 23167 17193
rect 23109 17153 23121 17187
rect 23155 17153 23167 17187
rect 23109 17147 23167 17153
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17153 23351 17187
rect 23293 17147 23351 17153
rect 20579 17088 20852 17116
rect 20579 17085 20591 17088
rect 20533 17079 20591 17085
rect 21174 17076 21180 17128
rect 21232 17076 21238 17128
rect 22554 17076 22560 17128
rect 22612 17116 22618 17128
rect 23308 17116 23336 17147
rect 25222 17144 25228 17196
rect 25280 17144 25286 17196
rect 25406 17144 25412 17196
rect 25464 17184 25470 17196
rect 26145 17187 26203 17193
rect 26145 17184 26157 17187
rect 25464 17156 26157 17184
rect 25464 17144 25470 17156
rect 26145 17153 26157 17156
rect 26191 17153 26203 17187
rect 27341 17187 27399 17193
rect 27341 17184 27353 17187
rect 26145 17147 26203 17153
rect 26252 17156 27353 17184
rect 22612 17088 23336 17116
rect 24765 17119 24823 17125
rect 22612 17076 22618 17088
rect 24765 17085 24777 17119
rect 24811 17116 24823 17119
rect 25038 17116 25044 17128
rect 24811 17088 25044 17116
rect 24811 17085 24823 17088
rect 24765 17079 24823 17085
rect 25038 17076 25044 17088
rect 25096 17076 25102 17128
rect 25130 17076 25136 17128
rect 25188 17076 25194 17128
rect 25866 17076 25872 17128
rect 25924 17076 25930 17128
rect 25961 17119 26019 17125
rect 25961 17085 25973 17119
rect 26007 17085 26019 17119
rect 25961 17079 26019 17085
rect 26053 17119 26111 17125
rect 26053 17085 26065 17119
rect 26099 17085 26111 17119
rect 26053 17079 26111 17085
rect 20438 17048 20444 17060
rect 18892 17020 20444 17048
rect 18785 17011 18843 17017
rect 4249 16983 4307 16989
rect 4249 16949 4261 16983
rect 4295 16980 4307 16983
rect 6454 16980 6460 16992
rect 4295 16952 6460 16980
rect 4295 16949 4307 16952
rect 4249 16943 4307 16949
rect 6454 16940 6460 16952
rect 6512 16940 6518 16992
rect 7006 16940 7012 16992
rect 7064 16940 7070 16992
rect 9582 16940 9588 16992
rect 9640 16980 9646 16992
rect 11149 16983 11207 16989
rect 11149 16980 11161 16983
rect 9640 16952 11161 16980
rect 9640 16940 9646 16952
rect 11149 16949 11161 16952
rect 11195 16980 11207 16983
rect 11698 16980 11704 16992
rect 11195 16952 11704 16980
rect 11195 16949 11207 16952
rect 11149 16943 11207 16949
rect 11698 16940 11704 16952
rect 11756 16940 11762 16992
rect 16390 16940 16396 16992
rect 16448 16940 16454 16992
rect 18800 16980 18828 17011
rect 20438 17008 20444 17020
rect 20496 17008 20502 17060
rect 20809 17051 20867 17057
rect 20809 17017 20821 17051
rect 20855 17048 20867 17051
rect 21192 17048 21220 17076
rect 20855 17020 21220 17048
rect 24581 17051 24639 17057
rect 20855 17017 20867 17020
rect 20809 17011 20867 17017
rect 24581 17017 24593 17051
rect 24627 17048 24639 17051
rect 25976 17048 26004 17079
rect 24627 17020 26004 17048
rect 24627 17017 24639 17020
rect 24581 17011 24639 17017
rect 20990 16980 20996 16992
rect 18800 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 25590 16940 25596 16992
rect 25648 16940 25654 16992
rect 25958 16940 25964 16992
rect 26016 16980 26022 16992
rect 26068 16980 26096 17079
rect 26252 16992 26280 17156
rect 27341 17153 27353 17156
rect 27387 17184 27399 17187
rect 27522 17184 27528 17196
rect 27387 17156 27528 17184
rect 27387 17153 27399 17156
rect 27341 17147 27399 17153
rect 27522 17144 27528 17156
rect 27580 17144 27586 17196
rect 27617 17187 27675 17193
rect 27617 17153 27629 17187
rect 27663 17153 27675 17187
rect 27617 17147 27675 17153
rect 27430 17076 27436 17128
rect 27488 17116 27494 17128
rect 27632 17116 27660 17147
rect 27798 17144 27804 17196
rect 27856 17144 27862 17196
rect 28460 17184 28488 17280
rect 28828 17193 28856 17280
rect 29380 17193 29408 17280
rect 30374 17212 30380 17264
rect 30432 17212 30438 17264
rect 28629 17187 28687 17193
rect 28629 17184 28641 17187
rect 28460 17156 28641 17184
rect 28629 17153 28641 17156
rect 28675 17153 28687 17187
rect 28629 17147 28687 17153
rect 28813 17187 28871 17193
rect 28813 17153 28825 17187
rect 28859 17153 28871 17187
rect 28813 17147 28871 17153
rect 29365 17187 29423 17193
rect 29365 17153 29377 17187
rect 29411 17153 29423 17187
rect 31665 17187 31723 17193
rect 31665 17184 31677 17187
rect 29365 17147 29423 17153
rect 31128 17156 31677 17184
rect 31128 17125 31156 17156
rect 31665 17153 31677 17156
rect 31711 17184 31723 17187
rect 31754 17184 31760 17196
rect 31711 17156 31760 17184
rect 31711 17153 31723 17156
rect 31665 17147 31723 17153
rect 31754 17144 31760 17156
rect 31812 17144 31818 17196
rect 31849 17187 31907 17193
rect 31849 17153 31861 17187
rect 31895 17184 31907 17187
rect 31938 17184 31944 17196
rect 31895 17156 31944 17184
rect 31895 17153 31907 17156
rect 31849 17147 31907 17153
rect 31938 17144 31944 17156
rect 31996 17144 32002 17196
rect 29641 17119 29699 17125
rect 29641 17116 29653 17119
rect 27488 17088 27660 17116
rect 29472 17088 29653 17116
rect 27488 17076 27494 17088
rect 28629 17051 28687 17057
rect 28629 17017 28641 17051
rect 28675 17048 28687 17051
rect 29472 17048 29500 17088
rect 29641 17085 29653 17088
rect 29687 17085 29699 17119
rect 29641 17079 29699 17085
rect 31113 17119 31171 17125
rect 31113 17085 31125 17119
rect 31159 17085 31171 17119
rect 31113 17079 31171 17085
rect 28675 17020 29500 17048
rect 28675 17017 28687 17020
rect 28629 17011 28687 17017
rect 26016 16952 26096 16980
rect 26016 16940 26022 16952
rect 26234 16940 26240 16992
rect 26292 16940 26298 16992
rect 1104 16890 35248 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 35248 16890
rect 1104 16816 35248 16838
rect 3234 16736 3240 16788
rect 3292 16736 3298 16788
rect 3786 16736 3792 16788
rect 3844 16736 3850 16788
rect 4172 16748 4844 16776
rect 1670 16600 1676 16652
rect 1728 16600 1734 16652
rect 3252 16640 3280 16736
rect 3970 16708 3976 16720
rect 3896 16680 3976 16708
rect 3252 16612 3464 16640
rect 1394 16532 1400 16584
rect 1452 16532 1458 16584
rect 3436 16581 3464 16612
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16541 3479 16575
rect 3896 16574 3924 16680
rect 3970 16668 3976 16680
rect 4028 16668 4034 16720
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 4172 16640 4200 16748
rect 4614 16708 4620 16720
rect 4120 16612 4200 16640
rect 4264 16680 4620 16708
rect 4264 16640 4292 16680
rect 4614 16668 4620 16680
rect 4672 16668 4678 16720
rect 4264 16612 4568 16640
rect 4120 16600 4126 16612
rect 3965 16575 4023 16581
rect 3965 16574 3977 16575
rect 3896 16546 3977 16574
rect 3421 16535 3479 16541
rect 3965 16541 3977 16546
rect 4011 16541 4023 16575
rect 3965 16535 4023 16541
rect 4154 16532 4160 16584
rect 4212 16532 4218 16584
rect 4264 16581 4292 16612
rect 4540 16581 4568 16612
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 4525 16575 4583 16581
rect 4525 16541 4537 16575
rect 4571 16541 4583 16575
rect 4688 16575 4746 16581
rect 4816 16578 4844 16748
rect 5074 16736 5080 16788
rect 5132 16776 5138 16788
rect 5169 16779 5227 16785
rect 5169 16776 5181 16779
rect 5132 16748 5181 16776
rect 5132 16736 5138 16748
rect 5169 16745 5181 16748
rect 5215 16745 5227 16779
rect 6822 16776 6828 16788
rect 5169 16739 5227 16745
rect 6196 16748 6828 16776
rect 5534 16668 5540 16720
rect 5592 16708 5598 16720
rect 6196 16708 6224 16748
rect 6822 16736 6828 16748
rect 6880 16776 6886 16788
rect 8205 16779 8263 16785
rect 8205 16776 8217 16779
rect 6880 16748 8217 16776
rect 6880 16736 6886 16748
rect 8205 16745 8217 16748
rect 8251 16776 8263 16779
rect 8662 16776 8668 16788
rect 8251 16748 8668 16776
rect 8251 16745 8263 16748
rect 8205 16739 8263 16745
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 9858 16736 9864 16788
rect 9916 16776 9922 16788
rect 11609 16779 11667 16785
rect 11609 16776 11621 16779
rect 9916 16748 11621 16776
rect 9916 16736 9922 16748
rect 11609 16745 11621 16748
rect 11655 16776 11667 16779
rect 12066 16776 12072 16788
rect 11655 16748 12072 16776
rect 11655 16745 11667 16748
rect 11609 16739 11667 16745
rect 12066 16736 12072 16748
rect 12124 16776 12130 16788
rect 12345 16779 12403 16785
rect 12345 16776 12357 16779
rect 12124 16748 12357 16776
rect 12124 16736 12130 16748
rect 12345 16745 12357 16748
rect 12391 16745 12403 16779
rect 12345 16739 12403 16745
rect 12805 16779 12863 16785
rect 12805 16745 12817 16779
rect 12851 16776 12863 16779
rect 12986 16776 12992 16788
rect 12851 16748 12992 16776
rect 12851 16745 12863 16748
rect 12805 16739 12863 16745
rect 12820 16708 12848 16739
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 15746 16736 15752 16788
rect 15804 16736 15810 16788
rect 16485 16779 16543 16785
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 17402 16776 17408 16788
rect 16531 16748 17408 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 17402 16736 17408 16748
rect 17460 16736 17466 16788
rect 18230 16736 18236 16788
rect 18288 16776 18294 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 18288 16748 19257 16776
rect 18288 16736 18294 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 19245 16739 19303 16745
rect 19978 16736 19984 16788
rect 20036 16736 20042 16788
rect 20438 16736 20444 16788
rect 20496 16736 20502 16788
rect 22370 16736 22376 16788
rect 22428 16776 22434 16788
rect 22465 16779 22523 16785
rect 22465 16776 22477 16779
rect 22428 16748 22477 16776
rect 22428 16736 22434 16748
rect 22465 16745 22477 16748
rect 22511 16745 22523 16779
rect 22465 16739 22523 16745
rect 22922 16736 22928 16788
rect 22980 16736 22986 16788
rect 23566 16736 23572 16788
rect 23624 16736 23630 16788
rect 25222 16736 25228 16788
rect 25280 16776 25286 16788
rect 25501 16779 25559 16785
rect 25501 16776 25513 16779
rect 25280 16748 25513 16776
rect 25280 16736 25286 16748
rect 25501 16745 25513 16748
rect 25547 16745 25559 16779
rect 25501 16739 25559 16745
rect 26234 16736 26240 16788
rect 26292 16736 26298 16788
rect 30098 16736 30104 16788
rect 30156 16736 30162 16788
rect 30374 16736 30380 16788
rect 30432 16736 30438 16788
rect 32214 16776 32220 16788
rect 31726 16748 32220 16776
rect 5592 16680 6224 16708
rect 5592 16668 5598 16680
rect 4688 16572 4700 16575
rect 4525 16535 4583 16541
rect 4632 16544 4700 16572
rect 3329 16507 3387 16513
rect 3329 16504 3341 16507
rect 2898 16476 3341 16504
rect 3329 16473 3341 16476
rect 3375 16473 3387 16507
rect 4448 16504 4476 16535
rect 4632 16504 4660 16544
rect 4688 16541 4700 16544
rect 4734 16541 4746 16575
rect 4688 16535 4746 16541
rect 4801 16572 4859 16578
rect 4801 16538 4813 16572
rect 4847 16538 4859 16572
rect 4801 16532 4859 16538
rect 4893 16575 4951 16581
rect 4893 16541 4905 16575
rect 4939 16574 4951 16575
rect 4982 16574 4988 16584
rect 4939 16546 4988 16574
rect 4939 16541 4951 16546
rect 4893 16535 4951 16541
rect 4982 16532 4988 16546
rect 5040 16532 5046 16584
rect 6196 16581 6224 16680
rect 12406 16680 12848 16708
rect 6454 16600 6460 16652
rect 6512 16600 6518 16652
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 9456 16612 9689 16640
rect 9456 16600 9462 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16640 11115 16643
rect 11977 16643 12035 16649
rect 11977 16640 11989 16643
rect 11103 16612 11989 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 11977 16609 11989 16612
rect 12023 16640 12035 16643
rect 12406 16640 12434 16680
rect 12023 16612 12434 16640
rect 15197 16643 15255 16649
rect 12023 16609 12035 16612
rect 11977 16603 12035 16609
rect 15197 16609 15209 16643
rect 15243 16640 15255 16643
rect 15764 16640 15792 16736
rect 15243 16612 15792 16640
rect 15243 16609 15255 16612
rect 15197 16603 15255 16609
rect 6181 16575 6239 16581
rect 6181 16541 6193 16575
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 14182 16532 14188 16584
rect 14240 16532 14246 16584
rect 14366 16532 14372 16584
rect 14424 16532 14430 16584
rect 15764 16581 15792 16612
rect 15841 16643 15899 16649
rect 15841 16609 15853 16643
rect 15887 16640 15899 16643
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 15887 16612 16037 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 16025 16609 16037 16612
rect 16071 16640 16083 16643
rect 16071 16612 17172 16640
rect 16071 16609 16083 16612
rect 16025 16603 16083 16609
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15749 16535 15807 16541
rect 15930 16532 15936 16584
rect 15988 16532 15994 16584
rect 16114 16532 16120 16584
rect 16172 16532 16178 16584
rect 16301 16575 16359 16581
rect 16301 16541 16313 16575
rect 16347 16572 16359 16575
rect 16390 16572 16396 16584
rect 16347 16544 16396 16572
rect 16347 16541 16359 16544
rect 16301 16535 16359 16541
rect 16390 16532 16396 16544
rect 16448 16532 16454 16584
rect 16666 16532 16672 16584
rect 16724 16532 16730 16584
rect 16850 16532 16856 16584
rect 16908 16532 16914 16584
rect 17144 16581 17172 16612
rect 19058 16600 19064 16652
rect 19116 16640 19122 16652
rect 19116 16612 19564 16640
rect 19116 16600 19122 16612
rect 17129 16575 17187 16581
rect 17129 16541 17141 16575
rect 17175 16541 17187 16575
rect 17129 16535 17187 16541
rect 17313 16575 17371 16581
rect 17313 16541 17325 16575
rect 17359 16572 17371 16575
rect 18322 16572 18328 16584
rect 17359 16544 18328 16572
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 18322 16532 18328 16544
rect 18380 16572 18386 16584
rect 18601 16575 18659 16581
rect 18601 16572 18613 16575
rect 18380 16544 18613 16572
rect 18380 16532 18386 16544
rect 18601 16541 18613 16544
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 18877 16575 18935 16581
rect 18877 16572 18889 16575
rect 18840 16544 18889 16572
rect 18840 16532 18846 16544
rect 18877 16541 18889 16544
rect 18923 16572 18935 16575
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 18923 16544 19441 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19536 16572 19564 16612
rect 19705 16575 19763 16581
rect 19705 16572 19717 16575
rect 19536 16544 19717 16572
rect 19429 16535 19487 16541
rect 19705 16541 19717 16544
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 3329 16467 3387 16473
rect 4080 16476 4660 16504
rect 4816 16504 4844 16532
rect 5258 16504 5264 16516
rect 4816 16476 5264 16504
rect 4080 16448 4108 16476
rect 3142 16396 3148 16448
rect 3200 16396 3206 16448
rect 4062 16396 4068 16448
rect 4120 16396 4126 16448
rect 4632 16436 4660 16476
rect 5258 16464 5264 16476
rect 5316 16464 5322 16516
rect 7006 16464 7012 16516
rect 7064 16464 7070 16516
rect 8941 16507 8999 16513
rect 8941 16504 8953 16507
rect 7944 16476 8953 16504
rect 6730 16436 6736 16448
rect 4632 16408 6736 16436
rect 6730 16396 6736 16408
rect 6788 16396 6794 16448
rect 7944 16445 7972 16476
rect 8941 16473 8953 16476
rect 8987 16473 8999 16507
rect 19904 16504 19932 16535
rect 8941 16467 8999 16473
rect 18708 16476 19932 16504
rect 18708 16448 18736 16476
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16405 7987 16439
rect 7929 16399 7987 16405
rect 10962 16396 10968 16448
rect 11020 16436 11026 16448
rect 13354 16436 13360 16448
rect 11020 16408 13360 16436
rect 11020 16396 11026 16408
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 18506 16396 18512 16448
rect 18564 16396 18570 16448
rect 18690 16396 18696 16448
rect 18748 16396 18754 16448
rect 19061 16439 19119 16445
rect 19061 16405 19073 16439
rect 19107 16436 19119 16439
rect 19996 16436 20024 16736
rect 20456 16572 20484 16736
rect 21361 16711 21419 16717
rect 21361 16677 21373 16711
rect 21407 16708 21419 16711
rect 22646 16708 22652 16720
rect 21407 16680 22652 16708
rect 21407 16677 21419 16680
rect 21361 16671 21419 16677
rect 21376 16640 21404 16671
rect 22646 16668 22652 16680
rect 22704 16668 22710 16720
rect 22940 16708 22968 16736
rect 29273 16711 29331 16717
rect 29273 16708 29285 16711
rect 22940 16680 29285 16708
rect 29273 16677 29285 16680
rect 29319 16677 29331 16711
rect 30116 16708 30144 16736
rect 30650 16708 30656 16720
rect 30116 16680 30656 16708
rect 29273 16671 29331 16677
rect 21008 16612 21404 16640
rect 20806 16572 20812 16584
rect 20456 16544 20812 16572
rect 20806 16532 20812 16544
rect 20864 16532 20870 16584
rect 21008 16581 21036 16612
rect 23566 16600 23572 16652
rect 23624 16600 23630 16652
rect 23658 16600 23664 16652
rect 23716 16640 23722 16652
rect 23716 16612 24164 16640
rect 23716 16600 23722 16612
rect 20993 16575 21051 16581
rect 20993 16541 21005 16575
rect 21039 16541 21051 16575
rect 23584 16572 23612 16600
rect 23750 16572 23756 16584
rect 23584 16544 23756 16572
rect 20993 16535 21051 16541
rect 23750 16532 23756 16544
rect 23808 16572 23814 16584
rect 24136 16581 24164 16612
rect 25406 16600 25412 16652
rect 25464 16600 25470 16652
rect 25590 16600 25596 16652
rect 25648 16640 25654 16652
rect 25777 16643 25835 16649
rect 25777 16640 25789 16643
rect 25648 16612 25789 16640
rect 25648 16600 25654 16612
rect 25777 16609 25789 16612
rect 25823 16609 25835 16643
rect 25777 16603 25835 16609
rect 23937 16575 23995 16581
rect 23937 16572 23949 16575
rect 23808 16544 23949 16572
rect 23808 16532 23814 16544
rect 23937 16541 23949 16544
rect 23983 16541 23995 16575
rect 23937 16535 23995 16541
rect 24121 16575 24179 16581
rect 24121 16541 24133 16575
rect 24167 16572 24179 16575
rect 24581 16575 24639 16581
rect 24581 16572 24593 16575
rect 24167 16544 24593 16572
rect 24167 16541 24179 16544
rect 24121 16535 24179 16541
rect 24581 16541 24593 16544
rect 24627 16541 24639 16575
rect 24581 16535 24639 16541
rect 24762 16532 24768 16584
rect 24820 16572 24826 16584
rect 24857 16575 24915 16581
rect 24857 16572 24869 16575
rect 24820 16544 24869 16572
rect 24820 16532 24826 16544
rect 24857 16541 24869 16544
rect 24903 16541 24915 16575
rect 24857 16535 24915 16541
rect 24946 16532 24952 16584
rect 25004 16572 25010 16584
rect 25041 16575 25099 16581
rect 25041 16572 25053 16575
rect 25004 16544 25053 16572
rect 25004 16532 25010 16544
rect 25041 16541 25053 16544
rect 25087 16541 25099 16575
rect 25041 16535 25099 16541
rect 25317 16575 25375 16581
rect 25317 16541 25329 16575
rect 25363 16572 25375 16575
rect 25424 16572 25452 16600
rect 25363 16544 25452 16572
rect 25363 16541 25375 16544
rect 25317 16535 25375 16541
rect 24029 16507 24087 16513
rect 24029 16473 24041 16507
rect 24075 16504 24087 16507
rect 25332 16504 25360 16535
rect 25866 16532 25872 16584
rect 25924 16572 25930 16584
rect 26142 16572 26148 16584
rect 25924 16544 26148 16572
rect 25924 16532 25930 16544
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 29288 16572 29316 16671
rect 30300 16581 30328 16680
rect 30650 16668 30656 16680
rect 30708 16708 30714 16720
rect 30745 16711 30803 16717
rect 30745 16708 30757 16711
rect 30708 16680 30757 16708
rect 30708 16668 30714 16680
rect 30745 16677 30757 16680
rect 30791 16677 30803 16711
rect 30745 16671 30803 16677
rect 31726 16640 31754 16748
rect 32214 16736 32220 16748
rect 32272 16776 32278 16788
rect 32674 16776 32680 16788
rect 32272 16748 32680 16776
rect 32272 16736 32278 16748
rect 32674 16736 32680 16748
rect 32732 16776 32738 16788
rect 32861 16779 32919 16785
rect 32861 16776 32873 16779
rect 32732 16748 32873 16776
rect 32732 16736 32738 16748
rect 32861 16745 32873 16748
rect 32907 16745 32919 16779
rect 32861 16739 32919 16745
rect 32309 16711 32367 16717
rect 32309 16677 32321 16711
rect 32355 16708 32367 16711
rect 33134 16708 33140 16720
rect 32355 16680 33140 16708
rect 32355 16677 32367 16680
rect 32309 16671 32367 16677
rect 33134 16668 33140 16680
rect 33192 16668 33198 16720
rect 31680 16612 31754 16640
rect 32033 16643 32091 16649
rect 29733 16575 29791 16581
rect 29733 16572 29745 16575
rect 29288 16544 29745 16572
rect 29733 16541 29745 16544
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16541 30067 16575
rect 30009 16535 30067 16541
rect 30285 16575 30343 16581
rect 30285 16541 30297 16575
rect 30331 16541 30343 16575
rect 30285 16535 30343 16541
rect 24075 16476 25360 16504
rect 30024 16504 30052 16535
rect 31386 16504 31392 16516
rect 30024 16476 31392 16504
rect 24075 16473 24087 16476
rect 24029 16467 24087 16473
rect 31386 16464 31392 16476
rect 31444 16504 31450 16516
rect 31680 16504 31708 16612
rect 32033 16609 32045 16643
rect 32079 16640 32091 16643
rect 32493 16643 32551 16649
rect 32493 16640 32505 16643
rect 32079 16612 32505 16640
rect 32079 16609 32091 16612
rect 32033 16603 32091 16609
rect 32493 16609 32505 16612
rect 32539 16609 32551 16643
rect 32493 16603 32551 16609
rect 32674 16600 32680 16652
rect 32732 16600 32738 16652
rect 31754 16532 31760 16584
rect 31812 16572 31818 16584
rect 31941 16575 31999 16581
rect 31941 16572 31953 16575
rect 31812 16544 31953 16572
rect 31812 16532 31818 16544
rect 31941 16541 31953 16544
rect 31987 16541 31999 16575
rect 31941 16535 31999 16541
rect 32401 16575 32459 16581
rect 32401 16541 32413 16575
rect 32447 16541 32459 16575
rect 32401 16535 32459 16541
rect 32585 16575 32643 16581
rect 32585 16541 32597 16575
rect 32631 16572 32643 16575
rect 32692 16572 32720 16600
rect 32631 16544 32720 16572
rect 32631 16541 32643 16544
rect 32585 16535 32643 16541
rect 32416 16504 32444 16535
rect 34514 16532 34520 16584
rect 34572 16532 34578 16584
rect 31444 16476 31708 16504
rect 31956 16476 32444 16504
rect 33597 16507 33655 16513
rect 31444 16464 31450 16476
rect 31956 16448 31984 16476
rect 33597 16473 33609 16507
rect 33643 16504 33655 16507
rect 34606 16504 34612 16516
rect 33643 16476 34612 16504
rect 33643 16473 33655 16476
rect 33597 16467 33655 16473
rect 34606 16464 34612 16476
rect 34664 16464 34670 16516
rect 19107 16408 20024 16436
rect 19107 16405 19119 16408
rect 19061 16399 19119 16405
rect 20990 16396 20996 16448
rect 21048 16396 21054 16448
rect 31938 16396 31944 16448
rect 31996 16396 32002 16448
rect 1104 16346 35236 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 35236 16346
rect 1104 16272 35236 16294
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 4154 16232 4160 16244
rect 3660 16204 4160 16232
rect 3660 16192 3666 16204
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 10321 16235 10379 16241
rect 10321 16201 10333 16235
rect 10367 16232 10379 16235
rect 10962 16232 10968 16244
rect 10367 16204 10968 16232
rect 10367 16201 10379 16204
rect 10321 16195 10379 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 12345 16235 12403 16241
rect 12345 16232 12357 16235
rect 11440 16204 12357 16232
rect 11440 16176 11468 16204
rect 12345 16201 12357 16204
rect 12391 16232 12403 16235
rect 13633 16235 13691 16241
rect 13633 16232 13645 16235
rect 12391 16204 13645 16232
rect 12391 16201 12403 16204
rect 12345 16195 12403 16201
rect 13633 16201 13645 16204
rect 13679 16232 13691 16235
rect 13906 16232 13912 16244
rect 13679 16204 13912 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 13906 16192 13912 16204
rect 13964 16192 13970 16244
rect 14001 16235 14059 16241
rect 14001 16201 14013 16235
rect 14047 16232 14059 16235
rect 14182 16232 14188 16244
rect 14047 16204 14188 16232
rect 14047 16201 14059 16204
rect 14001 16195 14059 16201
rect 14182 16192 14188 16204
rect 14240 16192 14246 16244
rect 14277 16235 14335 16241
rect 14277 16201 14289 16235
rect 14323 16232 14335 16235
rect 14366 16232 14372 16244
rect 14323 16204 14372 16232
rect 14323 16201 14335 16204
rect 14277 16195 14335 16201
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 18233 16235 18291 16241
rect 18233 16232 18245 16235
rect 16080 16204 18245 16232
rect 16080 16192 16086 16204
rect 18233 16201 18245 16204
rect 18279 16201 18291 16235
rect 18233 16195 18291 16201
rect 3329 16167 3387 16173
rect 3329 16164 3341 16167
rect 2746 16136 3341 16164
rect 1394 15852 1400 15904
rect 1452 15892 1458 15904
rect 2746 15892 2774 16136
rect 3329 16133 3341 16136
rect 3375 16164 3387 16167
rect 3786 16164 3792 16176
rect 3375 16136 3792 16164
rect 3375 16133 3387 16136
rect 3329 16127 3387 16133
rect 3786 16124 3792 16136
rect 3844 16164 3850 16176
rect 5534 16164 5540 16176
rect 3844 16136 5540 16164
rect 3844 16124 3850 16136
rect 5534 16124 5540 16136
rect 5592 16124 5598 16176
rect 11422 16124 11428 16176
rect 11480 16124 11486 16176
rect 11514 16124 11520 16176
rect 11572 16164 11578 16176
rect 11572 16136 11836 16164
rect 11572 16124 11578 16136
rect 6362 16056 6368 16108
rect 6420 16056 6426 16108
rect 9953 16099 10011 16105
rect 9953 16065 9965 16099
rect 9999 16096 10011 16099
rect 11054 16096 11060 16108
rect 9999 16068 11060 16096
rect 9999 16065 10011 16068
rect 9953 16059 10011 16065
rect 11054 16056 11060 16068
rect 11112 16056 11118 16108
rect 11149 16099 11207 16105
rect 11149 16065 11161 16099
rect 11195 16096 11207 16099
rect 11238 16096 11244 16108
rect 11195 16068 11244 16096
rect 11195 16065 11207 16068
rect 11149 16059 11207 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16096 11391 16099
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 11379 16068 11713 16096
rect 11379 16065 11391 16068
rect 11333 16059 11391 16065
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11808 16096 11836 16136
rect 11882 16124 11888 16176
rect 11940 16164 11946 16176
rect 12526 16164 12532 16176
rect 11940 16136 12532 16164
rect 11940 16124 11946 16136
rect 12526 16124 12532 16136
rect 12584 16124 12590 16176
rect 13354 16124 13360 16176
rect 13412 16164 13418 16176
rect 18248 16164 18276 16195
rect 18690 16192 18696 16244
rect 18748 16232 18754 16244
rect 19245 16235 19303 16241
rect 19245 16232 19257 16235
rect 18748 16204 19257 16232
rect 18748 16192 18754 16204
rect 19245 16201 19257 16204
rect 19291 16201 19303 16235
rect 22925 16235 22983 16241
rect 22925 16232 22937 16235
rect 19245 16195 19303 16201
rect 22112 16204 22937 16232
rect 13412 16136 14228 16164
rect 18248 16136 18644 16164
rect 13412 16124 13418 16136
rect 12434 16096 12440 16108
rect 11808 16068 12440 16096
rect 11701 16059 11759 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 14016 16105 14044 16136
rect 14200 16108 14228 16136
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 14001 16099 14059 16105
rect 14001 16065 14013 16099
rect 14047 16065 14059 16099
rect 14001 16059 14059 16065
rect 11793 16031 11851 16037
rect 11793 15997 11805 16031
rect 11839 16028 11851 16031
rect 12161 16031 12219 16037
rect 12161 16028 12173 16031
rect 11839 16000 12173 16028
rect 11839 15997 11851 16000
rect 11793 15991 11851 15997
rect 12161 15997 12173 16000
rect 12207 15997 12219 16031
rect 12452 16028 12480 16056
rect 13832 16028 13860 16059
rect 14090 16056 14096 16108
rect 14148 16056 14154 16108
rect 14182 16056 14188 16108
rect 14240 16056 14246 16108
rect 14274 16056 14280 16108
rect 14332 16096 14338 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14332 16068 14657 16096
rect 14332 16056 14338 16068
rect 14645 16065 14657 16068
rect 14691 16096 14703 16099
rect 16022 16096 16028 16108
rect 14691 16068 16028 16096
rect 14691 16065 14703 16068
rect 14645 16059 14703 16065
rect 16022 16056 16028 16068
rect 16080 16056 16086 16108
rect 18616 16105 18644 16136
rect 18874 16124 18880 16176
rect 18932 16164 18938 16176
rect 19061 16167 19119 16173
rect 19061 16164 19073 16167
rect 18932 16136 19073 16164
rect 18932 16124 18938 16136
rect 19061 16133 19073 16136
rect 19107 16164 19119 16167
rect 19107 16136 19288 16164
rect 19107 16133 19119 16136
rect 19061 16127 19119 16133
rect 19260 16108 19288 16136
rect 18417 16099 18475 16105
rect 18417 16096 18429 16099
rect 17880 16068 18429 16096
rect 15378 16028 15384 16040
rect 12452 16000 15384 16028
rect 12161 15991 12219 15997
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 10689 15963 10747 15969
rect 10689 15929 10701 15963
rect 10735 15960 10747 15963
rect 10781 15963 10839 15969
rect 10781 15960 10793 15963
rect 10735 15932 10793 15960
rect 10735 15929 10747 15932
rect 10689 15923 10747 15929
rect 10781 15929 10793 15932
rect 10827 15960 10839 15963
rect 16301 15963 16359 15969
rect 16301 15960 16313 15963
rect 10827 15932 11836 15960
rect 10827 15929 10839 15932
rect 10781 15923 10839 15929
rect 11808 15904 11836 15932
rect 15580 15932 16313 15960
rect 1452 15864 2774 15892
rect 3697 15895 3755 15901
rect 1452 15852 1458 15864
rect 3697 15861 3709 15895
rect 3743 15892 3755 15895
rect 4062 15892 4068 15904
rect 3743 15864 4068 15892
rect 3743 15861 3755 15864
rect 3697 15855 3755 15861
rect 4062 15852 4068 15864
rect 4120 15892 4126 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 4120 15864 4353 15892
rect 4120 15852 4126 15864
rect 4341 15861 4353 15864
rect 4387 15861 4399 15895
rect 4341 15855 4399 15861
rect 6549 15895 6607 15901
rect 6549 15861 6561 15895
rect 6595 15892 6607 15895
rect 6914 15892 6920 15904
rect 6595 15864 6920 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 11790 15852 11796 15904
rect 11848 15852 11854 15904
rect 11974 15852 11980 15904
rect 12032 15852 12038 15904
rect 12158 15852 12164 15904
rect 12216 15892 12222 15904
rect 12710 15892 12716 15904
rect 12216 15864 12716 15892
rect 12216 15852 12222 15864
rect 12710 15852 12716 15864
rect 12768 15892 12774 15904
rect 15580 15892 15608 15932
rect 16301 15929 16313 15932
rect 16347 15960 16359 15963
rect 16758 15960 16764 15972
rect 16347 15932 16764 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 16758 15920 16764 15932
rect 16816 15960 16822 15972
rect 17218 15960 17224 15972
rect 16816 15932 17224 15960
rect 16816 15920 16822 15932
rect 17218 15920 17224 15932
rect 17276 15920 17282 15972
rect 12768 15864 15608 15892
rect 12768 15852 12774 15864
rect 15654 15852 15660 15904
rect 15712 15852 15718 15904
rect 17770 15852 17776 15904
rect 17828 15892 17834 15904
rect 17880 15901 17908 16068
rect 18417 16065 18429 16068
rect 18463 16065 18475 16099
rect 18417 16059 18475 16065
rect 18601 16099 18659 16105
rect 18601 16065 18613 16099
rect 18647 16065 18659 16099
rect 18601 16059 18659 16065
rect 19242 16056 19248 16108
rect 19300 16056 19306 16108
rect 19429 16099 19487 16105
rect 19429 16065 19441 16099
rect 19475 16096 19487 16099
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19475 16068 19717 16096
rect 19475 16065 19487 16068
rect 19429 16059 19487 16065
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 19334 15988 19340 16040
rect 19392 16028 19398 16040
rect 19444 16028 19472 16059
rect 22112 16037 22140 16204
rect 22925 16201 22937 16204
rect 22971 16201 22983 16235
rect 22925 16195 22983 16201
rect 25130 16192 25136 16244
rect 25188 16232 25194 16244
rect 25225 16235 25283 16241
rect 25225 16232 25237 16235
rect 25188 16204 25237 16232
rect 25188 16192 25194 16204
rect 25225 16201 25237 16204
rect 25271 16201 25283 16235
rect 27433 16235 27491 16241
rect 27433 16232 27445 16235
rect 25225 16195 25283 16201
rect 27080 16204 27445 16232
rect 22741 16167 22799 16173
rect 22741 16164 22753 16167
rect 22204 16136 22753 16164
rect 22204 16105 22232 16136
rect 22741 16133 22753 16136
rect 22787 16133 22799 16167
rect 22741 16127 22799 16133
rect 27080 16108 27108 16204
rect 27433 16201 27445 16204
rect 27479 16201 27491 16235
rect 27433 16195 27491 16201
rect 27798 16192 27804 16244
rect 27856 16192 27862 16244
rect 34514 16192 34520 16244
rect 34572 16232 34578 16244
rect 34701 16235 34759 16241
rect 34701 16232 34713 16235
rect 34572 16204 34713 16232
rect 34572 16192 34578 16204
rect 34701 16201 34713 16204
rect 34747 16201 34759 16235
rect 34701 16195 34759 16201
rect 27356 16136 28212 16164
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 22370 16056 22376 16108
rect 22428 16096 22434 16108
rect 22649 16099 22707 16105
rect 22649 16096 22661 16099
rect 22428 16068 22661 16096
rect 22428 16056 22434 16068
rect 22649 16065 22661 16068
rect 22695 16065 22707 16099
rect 22649 16059 22707 16065
rect 22833 16099 22891 16105
rect 22833 16065 22845 16099
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 19392 16000 19472 16028
rect 22097 16031 22155 16037
rect 19392 15988 19398 16000
rect 22097 15997 22109 16031
rect 22143 15997 22155 16031
rect 22097 15991 22155 15997
rect 22554 15988 22560 16040
rect 22612 15988 22618 16040
rect 22848 16028 22876 16059
rect 22922 16056 22928 16108
rect 22980 16056 22986 16108
rect 23106 16056 23112 16108
rect 23164 16096 23170 16108
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 23164 16068 23397 16096
rect 23164 16056 23170 16068
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 24118 16056 24124 16108
rect 24176 16096 24182 16108
rect 24762 16096 24768 16108
rect 24176 16068 24768 16096
rect 24176 16056 24182 16068
rect 24762 16056 24768 16068
rect 24820 16096 24826 16108
rect 25958 16096 25964 16108
rect 24820 16068 25964 16096
rect 24820 16056 24826 16068
rect 25958 16056 25964 16068
rect 26016 16056 26022 16108
rect 27062 16056 27068 16108
rect 27120 16056 27126 16108
rect 27154 16056 27160 16108
rect 27212 16096 27218 16108
rect 27356 16105 27384 16136
rect 27341 16099 27399 16105
rect 27341 16096 27353 16099
rect 27212 16068 27353 16096
rect 27212 16056 27218 16068
rect 27341 16065 27353 16068
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 27522 16056 27528 16108
rect 27580 16096 27586 16108
rect 28184 16105 28212 16136
rect 33134 16124 33140 16176
rect 33192 16164 33198 16176
rect 33229 16167 33287 16173
rect 33229 16164 33241 16167
rect 33192 16136 33241 16164
rect 33192 16124 33198 16136
rect 33229 16133 33241 16136
rect 33275 16133 33287 16167
rect 33229 16127 33287 16133
rect 33962 16124 33968 16176
rect 34020 16124 34026 16176
rect 27617 16099 27675 16105
rect 27617 16096 27629 16099
rect 27580 16068 27629 16096
rect 27580 16056 27586 16068
rect 27617 16065 27629 16068
rect 27663 16065 27675 16099
rect 27617 16059 27675 16065
rect 28169 16099 28227 16105
rect 28169 16065 28181 16099
rect 28215 16065 28227 16099
rect 28169 16059 28227 16065
rect 22664 16000 22876 16028
rect 22664 15972 22692 16000
rect 17954 15920 17960 15972
rect 18012 15960 18018 15972
rect 21450 15960 21456 15972
rect 18012 15932 21456 15960
rect 18012 15920 18018 15932
rect 21450 15920 21456 15932
rect 21508 15920 21514 15972
rect 22646 15920 22652 15972
rect 22704 15920 22710 15972
rect 17865 15895 17923 15901
rect 17865 15892 17877 15895
rect 17828 15864 17877 15892
rect 17828 15852 17834 15864
rect 17865 15861 17877 15864
rect 17911 15861 17923 15895
rect 17865 15855 17923 15861
rect 18414 15852 18420 15904
rect 18472 15892 18478 15904
rect 18509 15895 18567 15901
rect 18509 15892 18521 15895
rect 18472 15864 18521 15892
rect 18472 15852 18478 15864
rect 18509 15861 18521 15864
rect 18555 15892 18567 15895
rect 18782 15892 18788 15904
rect 18555 15864 18788 15892
rect 18555 15861 18567 15864
rect 18509 15855 18567 15861
rect 18782 15852 18788 15864
rect 18840 15852 18846 15904
rect 20165 15895 20223 15901
rect 20165 15861 20177 15895
rect 20211 15892 20223 15895
rect 20346 15892 20352 15904
rect 20211 15864 20352 15892
rect 20211 15861 20223 15864
rect 20165 15855 20223 15861
rect 20346 15852 20352 15864
rect 20404 15892 20410 15904
rect 22940 15892 22968 16056
rect 27080 16028 27108 16056
rect 27985 16031 28043 16037
rect 27985 16028 27997 16031
rect 27080 16000 27997 16028
rect 27985 15997 27997 16000
rect 28031 15997 28043 16031
rect 32953 16031 33011 16037
rect 32953 16028 32965 16031
rect 27985 15991 28043 15997
rect 32784 16000 32965 16028
rect 32784 15904 32812 16000
rect 32953 15997 32965 16000
rect 32999 15997 33011 16031
rect 32953 15991 33011 15997
rect 20404 15864 22968 15892
rect 23845 15895 23903 15901
rect 20404 15852 20410 15864
rect 23845 15861 23857 15895
rect 23891 15892 23903 15895
rect 23934 15892 23940 15904
rect 23891 15864 23940 15892
rect 23891 15861 23903 15864
rect 23845 15855 23903 15861
rect 23934 15852 23940 15864
rect 23992 15852 23998 15904
rect 25041 15895 25099 15901
rect 25041 15861 25053 15895
rect 25087 15892 25099 15895
rect 25406 15892 25412 15904
rect 25087 15864 25412 15892
rect 25087 15861 25099 15864
rect 25041 15855 25099 15861
rect 25406 15852 25412 15864
rect 25464 15852 25470 15904
rect 28350 15852 28356 15904
rect 28408 15852 28414 15904
rect 32766 15852 32772 15904
rect 32824 15852 32830 15904
rect 1104 15802 35248 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 35248 15802
rect 1104 15728 35248 15750
rect 3602 15648 3608 15700
rect 3660 15648 3666 15700
rect 4614 15648 4620 15700
rect 4672 15688 4678 15700
rect 4801 15691 4859 15697
rect 4801 15688 4813 15691
rect 4672 15660 4813 15688
rect 4672 15648 4678 15660
rect 4801 15657 4813 15660
rect 4847 15657 4859 15691
rect 4801 15651 4859 15657
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 9125 15691 9183 15697
rect 9125 15688 9137 15691
rect 8720 15660 9137 15688
rect 8720 15648 8726 15660
rect 9125 15657 9137 15660
rect 9171 15657 9183 15691
rect 9125 15651 9183 15657
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 13449 15691 13507 15697
rect 13449 15688 13461 15691
rect 12492 15660 13461 15688
rect 12492 15648 12498 15660
rect 13449 15657 13461 15660
rect 13495 15657 13507 15691
rect 15654 15688 15660 15700
rect 13449 15651 13507 15657
rect 15120 15660 15660 15688
rect 1394 15580 1400 15632
rect 1452 15620 1458 15632
rect 1452 15592 1900 15620
rect 1452 15580 1458 15592
rect 1872 15561 1900 15592
rect 11054 15580 11060 15632
rect 11112 15620 11118 15632
rect 15120 15620 15148 15660
rect 15654 15648 15660 15660
rect 15712 15648 15718 15700
rect 15930 15648 15936 15700
rect 15988 15648 15994 15700
rect 18138 15688 18144 15700
rect 16500 15660 18144 15688
rect 16500 15620 16528 15660
rect 18138 15648 18144 15660
rect 18196 15648 18202 15700
rect 21450 15648 21456 15700
rect 21508 15688 21514 15700
rect 22833 15691 22891 15697
rect 21508 15660 22094 15688
rect 21508 15648 21514 15660
rect 11112 15592 15148 15620
rect 15580 15592 16528 15620
rect 16577 15623 16635 15629
rect 11112 15580 11118 15592
rect 1857 15555 1915 15561
rect 1857 15521 1869 15555
rect 1903 15521 1915 15555
rect 1857 15515 1915 15521
rect 3694 15512 3700 15564
rect 3752 15552 3758 15564
rect 3878 15552 3884 15564
rect 3752 15524 3884 15552
rect 3752 15512 3758 15524
rect 3878 15512 3884 15524
rect 3936 15552 3942 15564
rect 3936 15524 4016 15552
rect 3936 15512 3942 15524
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 3988 15493 4016 15524
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 15105 15555 15163 15561
rect 12032 15524 13952 15552
rect 12032 15512 12038 15524
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 4982 15484 4988 15496
rect 4862 15459 4988 15484
rect 3973 15447 4031 15453
rect 4847 15456 4988 15459
rect 4847 15453 4905 15456
rect 2133 15419 2191 15425
rect 2133 15416 2145 15419
rect 1596 15388 2145 15416
rect 1596 15357 1624 15388
rect 2133 15385 2145 15388
rect 2179 15385 2191 15419
rect 3881 15419 3939 15425
rect 3881 15416 3893 15419
rect 3358 15388 3893 15416
rect 2133 15379 2191 15385
rect 3881 15385 3893 15388
rect 3927 15385 3939 15419
rect 3881 15379 3939 15385
rect 4062 15376 4068 15428
rect 4120 15416 4126 15428
rect 4433 15419 4491 15425
rect 4433 15416 4445 15419
rect 4120 15388 4445 15416
rect 4120 15376 4126 15388
rect 4433 15385 4445 15388
rect 4479 15416 4491 15419
rect 4617 15419 4675 15425
rect 4617 15416 4629 15419
rect 4479 15388 4629 15416
rect 4479 15385 4491 15388
rect 4433 15379 4491 15385
rect 4617 15385 4629 15388
rect 4663 15385 4675 15419
rect 4847 15419 4859 15453
rect 4893 15419 4905 15453
rect 4982 15444 4988 15456
rect 5040 15444 5046 15496
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 7837 15487 7895 15493
rect 7837 15484 7849 15487
rect 7515 15456 7849 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 7837 15453 7849 15456
rect 7883 15484 7895 15487
rect 8297 15487 8355 15493
rect 8297 15484 8309 15487
rect 7883 15456 8309 15484
rect 7883 15453 7895 15456
rect 7837 15447 7895 15453
rect 8297 15453 8309 15456
rect 8343 15484 8355 15487
rect 8343 15456 8708 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 4847 15416 4905 15419
rect 4617 15379 4675 15385
rect 4832 15413 4905 15416
rect 4832 15388 4890 15413
rect 4832 15360 4860 15388
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15317 1639 15351
rect 1581 15311 1639 15317
rect 3602 15308 3608 15360
rect 3660 15348 3666 15360
rect 3970 15348 3976 15360
rect 3660 15320 3976 15348
rect 3660 15308 3666 15320
rect 3970 15308 3976 15320
rect 4028 15348 4034 15360
rect 4798 15348 4804 15360
rect 4028 15320 4804 15348
rect 4028 15308 4034 15320
rect 4798 15308 4804 15320
rect 4856 15308 4862 15360
rect 4982 15308 4988 15360
rect 5040 15308 5046 15360
rect 7377 15351 7435 15357
rect 7377 15317 7389 15351
rect 7423 15348 7435 15351
rect 7466 15348 7472 15360
rect 7423 15320 7472 15348
rect 7423 15317 7435 15320
rect 7377 15311 7435 15317
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 8205 15351 8263 15357
rect 8205 15317 8217 15351
rect 8251 15348 8263 15351
rect 8294 15348 8300 15360
rect 8251 15320 8300 15348
rect 8251 15317 8263 15320
rect 8205 15311 8263 15317
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 8680 15357 8708 15456
rect 12526 15444 12532 15496
rect 12584 15444 12590 15496
rect 8665 15351 8723 15357
rect 8665 15317 8677 15351
rect 8711 15348 8723 15351
rect 8754 15348 8760 15360
rect 8711 15320 8760 15348
rect 8711 15317 8723 15320
rect 8665 15311 8723 15317
rect 8754 15308 8760 15320
rect 8812 15308 8818 15360
rect 10505 15351 10563 15357
rect 10505 15317 10517 15351
rect 10551 15348 10563 15351
rect 11238 15348 11244 15360
rect 10551 15320 11244 15348
rect 10551 15317 10563 15320
rect 10505 15311 10563 15317
rect 11238 15308 11244 15320
rect 11296 15308 11302 15360
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11422 15348 11428 15360
rect 11379 15320 11428 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11422 15308 11428 15320
rect 11480 15308 11486 15360
rect 11514 15308 11520 15360
rect 11572 15348 11578 15360
rect 11609 15351 11667 15357
rect 11609 15348 11621 15351
rect 11572 15320 11621 15348
rect 11572 15308 11578 15320
rect 11609 15317 11621 15320
rect 11655 15317 11667 15351
rect 11609 15311 11667 15317
rect 12069 15351 12127 15357
rect 12069 15317 12081 15351
rect 12115 15348 12127 15351
rect 12158 15348 12164 15360
rect 12115 15320 12164 15348
rect 12115 15317 12127 15320
rect 12069 15311 12127 15317
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 12437 15351 12495 15357
rect 12437 15317 12449 15351
rect 12483 15348 12495 15351
rect 12544 15348 12572 15444
rect 13924 15416 13952 15524
rect 15105 15521 15117 15555
rect 15151 15552 15163 15555
rect 15580 15552 15608 15592
rect 16577 15589 16589 15623
rect 16623 15589 16635 15623
rect 20254 15620 20260 15632
rect 16577 15583 16635 15589
rect 17788 15592 20260 15620
rect 16592 15552 16620 15583
rect 16942 15552 16948 15564
rect 15151 15524 15608 15552
rect 15672 15524 16948 15552
rect 15151 15521 15163 15524
rect 15105 15515 15163 15521
rect 15672 15496 15700 15524
rect 16942 15512 16948 15524
rect 17000 15512 17006 15564
rect 17052 15524 17448 15552
rect 17052 15496 17080 15524
rect 14182 15444 14188 15496
rect 14240 15444 14246 15496
rect 14366 15444 14372 15496
rect 14424 15444 14430 15496
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 15473 15487 15531 15493
rect 15473 15453 15485 15487
rect 15519 15453 15531 15487
rect 15473 15447 15531 15453
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15453 15623 15487
rect 15565 15447 15623 15453
rect 15488 15416 15516 15447
rect 13924 15388 15516 15416
rect 15580 15416 15608 15447
rect 15654 15444 15660 15496
rect 15712 15444 15718 15496
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 15804 15456 15976 15484
rect 15804 15444 15810 15456
rect 15948 15416 15976 15456
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15453 16267 15487
rect 16209 15447 16267 15453
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 16485 15487 16543 15493
rect 16485 15484 16497 15487
rect 16439 15456 16497 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 16485 15453 16497 15456
rect 16531 15453 16543 15487
rect 16485 15447 16543 15453
rect 16224 15416 16252 15447
rect 17034 15444 17040 15496
rect 17092 15444 17098 15496
rect 17126 15444 17132 15496
rect 17184 15444 17190 15496
rect 17218 15444 17224 15496
rect 17276 15484 17282 15496
rect 17420 15484 17448 15524
rect 17788 15496 17816 15592
rect 20254 15580 20260 15592
rect 20312 15580 20318 15632
rect 20438 15580 20444 15632
rect 20496 15620 20502 15632
rect 22066 15620 22094 15660
rect 22833 15657 22845 15691
rect 22879 15688 22891 15691
rect 22922 15688 22928 15700
rect 22879 15660 22928 15688
rect 22879 15657 22891 15660
rect 22833 15651 22891 15657
rect 22922 15648 22928 15660
rect 22980 15648 22986 15700
rect 26970 15648 26976 15700
rect 27028 15688 27034 15700
rect 27028 15660 28212 15688
rect 27028 15648 27034 15660
rect 22278 15620 22284 15632
rect 20496 15592 20944 15620
rect 22066 15592 22284 15620
rect 20496 15580 20502 15592
rect 20070 15512 20076 15564
rect 20128 15552 20134 15564
rect 20128 15524 20484 15552
rect 20128 15512 20134 15524
rect 17770 15484 17776 15496
rect 17276 15456 17356 15484
rect 17420 15481 17632 15484
rect 17696 15481 17776 15484
rect 17420 15456 17776 15481
rect 17276 15444 17282 15456
rect 15580 15388 15792 15416
rect 15948 15388 16252 15416
rect 17328 15416 17356 15456
rect 17604 15453 17724 15456
rect 17770 15444 17776 15456
rect 17828 15444 17834 15496
rect 18138 15444 18144 15496
rect 18196 15444 18202 15496
rect 18506 15444 18512 15496
rect 18564 15484 18570 15496
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 18564 15456 19533 15484
rect 18564 15444 18570 15456
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 20346 15484 20352 15496
rect 19659 15456 20352 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 20346 15444 20352 15456
rect 20404 15444 20410 15496
rect 20456 15493 20484 15524
rect 20916 15493 20944 15592
rect 22278 15580 22284 15592
rect 22336 15620 22342 15632
rect 23109 15623 23167 15629
rect 23109 15620 23121 15623
rect 22336 15592 23121 15620
rect 22336 15580 22342 15592
rect 23109 15589 23121 15592
rect 23155 15589 23167 15623
rect 23109 15583 23167 15589
rect 27249 15623 27307 15629
rect 27249 15589 27261 15623
rect 27295 15589 27307 15623
rect 27249 15583 27307 15589
rect 28184 15620 28212 15660
rect 33962 15648 33968 15700
rect 34020 15648 34026 15700
rect 28184 15592 29868 15620
rect 20990 15512 20996 15564
rect 21048 15512 21054 15564
rect 21729 15555 21787 15561
rect 21729 15521 21741 15555
rect 21775 15552 21787 15555
rect 21775 15524 22094 15552
rect 21775 15521 21787 15524
rect 21729 15515 21787 15521
rect 20441 15487 20499 15493
rect 20441 15453 20453 15487
rect 20487 15453 20499 15487
rect 20441 15447 20499 15453
rect 20901 15487 20959 15493
rect 20901 15453 20913 15487
rect 20947 15453 20959 15487
rect 22066 15484 22094 15524
rect 23124 15484 23152 15583
rect 23569 15555 23627 15561
rect 23569 15521 23581 15555
rect 23615 15552 23627 15555
rect 24673 15555 24731 15561
rect 24673 15552 24685 15555
rect 23615 15524 24685 15552
rect 23615 15521 23627 15524
rect 23569 15515 23627 15521
rect 24673 15521 24685 15524
rect 24719 15521 24731 15555
rect 24673 15515 24731 15521
rect 23477 15487 23535 15493
rect 23477 15484 23489 15487
rect 22066 15456 23060 15484
rect 23124 15456 23489 15484
rect 20901 15447 20959 15453
rect 18969 15419 19027 15425
rect 18969 15416 18981 15419
rect 17328 15388 18981 15416
rect 15764 15360 15792 15388
rect 12483 15320 12572 15348
rect 12483 15317 12495 15320
rect 12437 15311 12495 15317
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 14274 15348 14280 15360
rect 13044 15320 14280 15348
rect 13044 15308 13050 15320
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 15746 15308 15752 15360
rect 15804 15308 15810 15360
rect 16224 15348 16252 15388
rect 18969 15385 18981 15388
rect 19015 15416 19027 15419
rect 19797 15419 19855 15425
rect 19797 15416 19809 15419
rect 19015 15388 19809 15416
rect 19015 15385 19027 15388
rect 18969 15379 19027 15385
rect 19797 15385 19809 15388
rect 19843 15416 19855 15419
rect 22370 15416 22376 15428
rect 19843 15388 22376 15416
rect 19843 15385 19855 15388
rect 19797 15379 19855 15385
rect 22370 15376 22376 15388
rect 22428 15376 22434 15428
rect 16482 15348 16488 15360
rect 16224 15320 16488 15348
rect 16482 15308 16488 15320
rect 16540 15308 16546 15360
rect 19058 15308 19064 15360
rect 19116 15348 19122 15360
rect 19245 15351 19303 15357
rect 19245 15348 19257 15351
rect 19116 15320 19257 15348
rect 19116 15308 19122 15320
rect 19245 15317 19257 15320
rect 19291 15317 19303 15351
rect 19245 15311 19303 15317
rect 19426 15308 19432 15360
rect 19484 15308 19490 15360
rect 22281 15351 22339 15357
rect 22281 15317 22293 15351
rect 22327 15348 22339 15351
rect 22554 15348 22560 15360
rect 22327 15320 22560 15348
rect 22327 15317 22339 15320
rect 22281 15311 22339 15317
rect 22554 15308 22560 15320
rect 22612 15308 22618 15360
rect 23032 15348 23060 15456
rect 23477 15453 23489 15456
rect 23523 15453 23535 15487
rect 23477 15447 23535 15453
rect 23658 15444 23664 15496
rect 23716 15444 23722 15496
rect 23750 15444 23756 15496
rect 23808 15493 23814 15496
rect 23808 15484 23817 15493
rect 23808 15456 23853 15484
rect 23808 15447 23817 15456
rect 23808 15444 23814 15447
rect 23934 15444 23940 15496
rect 23992 15444 23998 15496
rect 25961 15487 26019 15493
rect 25961 15484 25973 15487
rect 23290 15376 23296 15428
rect 23348 15416 23354 15428
rect 23676 15416 23704 15444
rect 23348 15388 23704 15416
rect 23845 15419 23903 15425
rect 23348 15376 23354 15388
rect 23845 15385 23857 15419
rect 23891 15416 23903 15419
rect 24596 15416 24624 15470
rect 25608 15456 25973 15484
rect 25608 15428 25636 15456
rect 25961 15453 25973 15456
rect 26007 15453 26019 15487
rect 25961 15447 26019 15453
rect 26973 15487 27031 15493
rect 26973 15453 26985 15487
rect 27019 15484 27031 15487
rect 27154 15484 27160 15496
rect 27019 15456 27160 15484
rect 27019 15453 27031 15456
rect 26973 15447 27031 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27264 15484 27292 15583
rect 28074 15512 28080 15564
rect 28132 15512 28138 15564
rect 27341 15487 27399 15493
rect 27341 15484 27353 15487
rect 27264 15456 27353 15484
rect 27341 15453 27353 15456
rect 27387 15453 27399 15487
rect 27341 15447 27399 15453
rect 27890 15444 27896 15496
rect 27948 15444 27954 15496
rect 28184 15493 28212 15592
rect 28350 15512 28356 15564
rect 28408 15512 28414 15564
rect 29840 15561 29868 15592
rect 29825 15555 29883 15561
rect 28644 15524 29776 15552
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15453 28227 15487
rect 28368 15484 28396 15512
rect 28644 15493 28672 15524
rect 29748 15493 29776 15524
rect 29825 15521 29837 15555
rect 29871 15521 29883 15555
rect 29825 15515 29883 15521
rect 30101 15555 30159 15561
rect 30101 15521 30113 15555
rect 30147 15552 30159 15555
rect 30469 15555 30527 15561
rect 30469 15552 30481 15555
rect 30147 15524 30481 15552
rect 30147 15521 30159 15524
rect 30101 15515 30159 15521
rect 30469 15521 30481 15524
rect 30515 15521 30527 15555
rect 30469 15515 30527 15521
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 28368 15456 28641 15484
rect 28169 15447 28227 15453
rect 28629 15453 28641 15456
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 29181 15487 29239 15493
rect 29181 15453 29193 15487
rect 29227 15453 29239 15487
rect 29181 15447 29239 15453
rect 29733 15487 29791 15493
rect 29733 15453 29745 15487
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 30561 15487 30619 15493
rect 30561 15453 30573 15487
rect 30607 15453 30619 15487
rect 30561 15447 30619 15453
rect 23891 15388 24624 15416
rect 25501 15419 25559 15425
rect 23891 15385 23903 15388
rect 23845 15379 23903 15385
rect 25501 15385 25513 15419
rect 25547 15416 25559 15419
rect 25590 15416 25596 15428
rect 25547 15388 25596 15416
rect 25547 15385 25559 15388
rect 25501 15379 25559 15385
rect 25590 15376 25596 15388
rect 25648 15376 25654 15428
rect 25976 15388 27200 15416
rect 25976 15348 26004 15388
rect 23032 15320 26004 15348
rect 26050 15308 26056 15360
rect 26108 15308 26114 15360
rect 26234 15308 26240 15360
rect 26292 15348 26298 15360
rect 27062 15348 27068 15360
rect 26292 15320 27068 15348
rect 26292 15308 26298 15320
rect 27062 15308 27068 15320
rect 27120 15308 27126 15360
rect 27172 15348 27200 15388
rect 27246 15376 27252 15428
rect 27304 15416 27310 15428
rect 27522 15416 27528 15428
rect 27304 15388 27528 15416
rect 27304 15376 27310 15388
rect 27522 15376 27528 15388
rect 27580 15416 27586 15428
rect 28350 15416 28356 15428
rect 27580 15388 28356 15416
rect 27580 15376 27586 15388
rect 28350 15376 28356 15388
rect 28408 15376 28414 15428
rect 28718 15376 28724 15428
rect 28776 15416 28782 15428
rect 29196 15416 29224 15447
rect 30576 15416 30604 15447
rect 33594 15444 33600 15496
rect 33652 15484 33658 15496
rect 33781 15487 33839 15493
rect 33781 15484 33793 15487
rect 33652 15456 33793 15484
rect 33652 15444 33658 15456
rect 33781 15453 33793 15456
rect 33827 15484 33839 15487
rect 33873 15487 33931 15493
rect 33873 15484 33885 15487
rect 33827 15456 33885 15484
rect 33827 15453 33839 15456
rect 33781 15447 33839 15453
rect 33873 15453 33885 15456
rect 33919 15453 33931 15487
rect 33873 15447 33931 15453
rect 28776 15388 30604 15416
rect 28776 15376 28782 15388
rect 27982 15348 27988 15360
rect 27172 15320 27988 15348
rect 27982 15308 27988 15320
rect 28040 15308 28046 15360
rect 30190 15308 30196 15360
rect 30248 15308 30254 15360
rect 1104 15258 35236 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 35236 15258
rect 1104 15184 35236 15206
rect 1486 15104 1492 15156
rect 1544 15104 1550 15156
rect 3786 15104 3792 15156
rect 3844 15104 3850 15156
rect 4798 15104 4804 15156
rect 4856 15104 4862 15156
rect 5721 15147 5779 15153
rect 5721 15113 5733 15147
rect 5767 15144 5779 15147
rect 6362 15144 6368 15156
rect 5767 15116 6368 15144
rect 5767 15113 5779 15116
rect 5721 15107 5779 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 13449 15147 13507 15153
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 14366 15144 14372 15156
rect 13495 15116 14372 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 14366 15104 14372 15116
rect 14424 15104 14430 15156
rect 15013 15147 15071 15153
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15286 15144 15292 15156
rect 15059 15116 15292 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15286 15104 15292 15116
rect 15344 15104 15350 15156
rect 15378 15104 15384 15156
rect 15436 15144 15442 15156
rect 15933 15147 15991 15153
rect 15436 15116 15516 15144
rect 15436 15104 15442 15116
rect 1504 15076 1532 15104
rect 1412 15048 1532 15076
rect 1412 15017 1440 15048
rect 1578 15036 1584 15088
rect 1636 15076 1642 15088
rect 1673 15079 1731 15085
rect 1673 15076 1685 15079
rect 1636 15048 1685 15076
rect 1636 15036 1642 15048
rect 1673 15045 1685 15048
rect 1719 15045 1731 15079
rect 1673 15039 1731 15045
rect 2314 15036 2320 15088
rect 2372 15036 2378 15088
rect 3804 15076 3832 15104
rect 4433 15079 4491 15085
rect 4433 15076 4445 15079
rect 3804 15048 4445 15076
rect 4433 15045 4445 15048
rect 4479 15045 4491 15079
rect 4816 15076 4844 15104
rect 4816 15048 5580 15076
rect 4433 15039 4491 15045
rect 1397 15011 1455 15017
rect 1397 14977 1409 15011
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 4801 15011 4859 15017
rect 4801 14977 4813 15011
rect 4847 15008 4859 15011
rect 5258 15008 5264 15020
rect 4847 14980 5264 15008
rect 4847 14977 4859 14980
rect 4801 14971 4859 14977
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14940 3203 14943
rect 4816 14940 4844 14971
rect 5258 14968 5264 14980
rect 5316 14968 5322 15020
rect 5552 15017 5580 15048
rect 6914 15036 6920 15088
rect 6972 15076 6978 15088
rect 7285 15079 7343 15085
rect 7285 15076 7297 15079
rect 6972 15048 7297 15076
rect 6972 15036 6978 15048
rect 7285 15045 7297 15048
rect 7331 15045 7343 15079
rect 7285 15039 7343 15045
rect 8294 15036 8300 15088
rect 8352 15036 8358 15088
rect 9858 15036 9864 15088
rect 9916 15036 9922 15088
rect 12253 15079 12311 15085
rect 12253 15045 12265 15079
rect 12299 15076 12311 15079
rect 12986 15076 12992 15088
rect 12299 15048 12992 15076
rect 12299 15045 12311 15048
rect 12253 15039 12311 15045
rect 5537 15011 5595 15017
rect 5537 14977 5549 15011
rect 5583 14977 5595 15011
rect 5537 14971 5595 14977
rect 8662 14968 8668 15020
rect 8720 14968 8726 15020
rect 9033 15011 9091 15017
rect 9033 15008 9045 15011
rect 8772 14980 9045 15008
rect 3191 14912 4844 14940
rect 4893 14943 4951 14949
rect 3191 14909 3203 14912
rect 3145 14903 3203 14909
rect 4893 14909 4905 14943
rect 4939 14940 4951 14943
rect 4982 14940 4988 14952
rect 4939 14912 4988 14940
rect 4939 14909 4951 14912
rect 4893 14903 4951 14909
rect 4982 14900 4988 14912
rect 5040 14900 5046 14952
rect 7009 14943 7067 14949
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 8294 14940 8300 14952
rect 7055 14912 8300 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 8294 14900 8300 14912
rect 8352 14940 8358 14952
rect 8680 14940 8708 14968
rect 8772 14949 8800 14980
rect 9033 14977 9045 14980
rect 9079 14977 9091 15011
rect 9033 14971 9091 14977
rect 11609 15011 11667 15017
rect 11609 14977 11621 15011
rect 11655 14977 11667 15011
rect 11609 14971 11667 14977
rect 8352 14912 8708 14940
rect 8757 14943 8815 14949
rect 8352 14900 8358 14912
rect 8757 14909 8769 14943
rect 8803 14909 8815 14943
rect 8757 14903 8815 14909
rect 11238 14900 11244 14952
rect 11296 14940 11302 14952
rect 11624 14940 11652 14971
rect 11790 14968 11796 15020
rect 11848 15008 11854 15020
rect 12268 15008 12296 15039
rect 12986 15036 12992 15048
rect 13044 15036 13050 15088
rect 15102 15076 15108 15088
rect 13096 15048 15108 15076
rect 11848 14980 12296 15008
rect 11848 14968 11854 14980
rect 12342 14968 12348 15020
rect 12400 14968 12406 15020
rect 13096 15017 13124 15048
rect 15102 15036 15108 15048
rect 15160 15076 15166 15088
rect 15488 15076 15516 15116
rect 15933 15113 15945 15147
rect 15979 15144 15991 15147
rect 16022 15144 16028 15156
rect 15979 15116 16028 15144
rect 15979 15113 15991 15116
rect 15933 15107 15991 15113
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 16666 15104 16672 15156
rect 16724 15144 16730 15156
rect 18969 15147 19027 15153
rect 18969 15144 18981 15147
rect 16724 15116 18981 15144
rect 16724 15104 16730 15116
rect 18969 15113 18981 15116
rect 19015 15113 19027 15147
rect 18969 15107 19027 15113
rect 19797 15147 19855 15153
rect 19797 15113 19809 15147
rect 19843 15144 19855 15147
rect 20346 15144 20352 15156
rect 19843 15116 20352 15144
rect 19843 15113 19855 15116
rect 19797 15107 19855 15113
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 20806 15104 20812 15156
rect 20864 15144 20870 15156
rect 21177 15147 21235 15153
rect 21177 15144 21189 15147
rect 20864 15116 21189 15144
rect 20864 15104 20870 15116
rect 21177 15113 21189 15116
rect 21223 15144 21235 15147
rect 21818 15144 21824 15156
rect 21223 15116 21824 15144
rect 21223 15113 21235 15116
rect 21177 15107 21235 15113
rect 21818 15104 21824 15116
rect 21876 15144 21882 15156
rect 22925 15147 22983 15153
rect 22925 15144 22937 15147
rect 21876 15116 22937 15144
rect 21876 15104 21882 15116
rect 22925 15113 22937 15116
rect 22971 15113 22983 15147
rect 22925 15107 22983 15113
rect 23750 15104 23756 15156
rect 23808 15104 23814 15156
rect 26142 15104 26148 15156
rect 26200 15144 26206 15156
rect 26605 15147 26663 15153
rect 26605 15144 26617 15147
rect 26200 15116 26617 15144
rect 26200 15104 26206 15116
rect 26605 15113 26617 15116
rect 26651 15113 26663 15147
rect 26605 15107 26663 15113
rect 27617 15147 27675 15153
rect 27617 15113 27629 15147
rect 27663 15144 27675 15147
rect 28074 15144 28080 15156
rect 27663 15116 28080 15144
rect 27663 15113 27675 15116
rect 27617 15107 27675 15113
rect 28074 15104 28080 15116
rect 28132 15104 28138 15156
rect 28350 15104 28356 15156
rect 28408 15104 28414 15156
rect 28718 15104 28724 15156
rect 28776 15104 28782 15156
rect 29362 15104 29368 15156
rect 29420 15144 29426 15156
rect 29825 15147 29883 15153
rect 29825 15144 29837 15147
rect 29420 15116 29837 15144
rect 29420 15104 29426 15116
rect 29825 15113 29837 15116
rect 29871 15113 29883 15147
rect 29825 15107 29883 15113
rect 16853 15079 16911 15085
rect 16853 15076 16865 15079
rect 15160 15048 15424 15076
rect 15488 15048 16865 15076
rect 15160 15036 15166 15048
rect 13081 15011 13139 15017
rect 13081 14977 13093 15011
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 14918 14968 14924 15020
rect 14976 14968 14982 15020
rect 15194 14968 15200 15020
rect 15252 14968 15258 15020
rect 15396 15017 15424 15048
rect 16853 15045 16865 15048
rect 16899 15076 16911 15079
rect 17034 15076 17040 15088
rect 16899 15048 17040 15076
rect 16899 15045 16911 15048
rect 16853 15039 16911 15045
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 18138 15076 18144 15088
rect 17328 15048 18144 15076
rect 15381 15011 15439 15017
rect 15381 14977 15393 15011
rect 15427 14977 15439 15011
rect 15381 14971 15439 14977
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 12360 14940 12388 14968
rect 11296 14912 12388 14940
rect 13173 14943 13231 14949
rect 11296 14900 11302 14912
rect 13173 14909 13185 14943
rect 13219 14940 13231 14943
rect 14826 14940 14832 14952
rect 13219 14912 14832 14940
rect 13219 14909 13231 14912
rect 13173 14903 13231 14909
rect 14826 14900 14832 14912
rect 14884 14940 14890 14952
rect 16316 14940 16344 14971
rect 17126 14968 17132 15020
rect 17184 14968 17190 15020
rect 17328 15017 17356 15048
rect 18138 15036 18144 15048
rect 18196 15036 18202 15088
rect 18690 15036 18696 15088
rect 18748 15036 18754 15088
rect 19426 15076 19432 15088
rect 19168 15048 19432 15076
rect 17313 15011 17371 15017
rect 17313 14977 17325 15011
rect 17359 14977 17371 15011
rect 18049 15011 18107 15017
rect 18049 15008 18061 15011
rect 17313 14971 17371 14977
rect 17420 14980 18061 15008
rect 17034 14940 17040 14952
rect 14884 14912 17040 14940
rect 14884 14900 14890 14912
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 17144 14940 17172 14968
rect 17420 14940 17448 14980
rect 18049 14977 18061 14980
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18233 15011 18291 15017
rect 18233 14977 18245 15011
rect 18279 15008 18291 15011
rect 18414 15008 18420 15020
rect 18279 14980 18420 15008
rect 18279 14977 18291 14980
rect 18233 14971 18291 14977
rect 17144 14912 17448 14940
rect 17494 14900 17500 14952
rect 17552 14900 17558 14952
rect 17678 14900 17684 14952
rect 17736 14900 17742 14952
rect 17310 14872 17316 14884
rect 12544 14844 17316 14872
rect 12544 14816 12572 14844
rect 17310 14832 17316 14844
rect 17368 14832 17374 14884
rect 3326 14764 3332 14816
rect 3384 14804 3390 14816
rect 3878 14804 3884 14816
rect 3384 14776 3884 14804
rect 3384 14764 3390 14776
rect 3878 14764 3884 14776
rect 3936 14804 3942 14816
rect 4065 14807 4123 14813
rect 4065 14804 4077 14807
rect 3936 14776 4077 14804
rect 3936 14764 3942 14776
rect 4065 14773 4077 14776
rect 4111 14773 4123 14807
rect 4065 14767 4123 14773
rect 5166 14764 5172 14816
rect 5224 14764 5230 14816
rect 11606 14764 11612 14816
rect 11664 14764 11670 14816
rect 12526 14764 12532 14816
rect 12584 14764 12590 14816
rect 15289 14807 15347 14813
rect 15289 14773 15301 14807
rect 15335 14804 15347 14807
rect 15746 14804 15752 14816
rect 15335 14776 15752 14804
rect 15335 14773 15347 14776
rect 15289 14767 15347 14773
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 16206 14764 16212 14816
rect 16264 14764 16270 14816
rect 18064 14804 18092 14971
rect 18414 14968 18420 14980
rect 18472 14968 18478 15020
rect 18509 15011 18567 15017
rect 18509 14977 18521 15011
rect 18555 15008 18567 15011
rect 18708 15008 18736 15036
rect 19168 15017 19196 15048
rect 19426 15036 19432 15048
rect 19484 15076 19490 15088
rect 20070 15076 20076 15088
rect 19484 15048 20076 15076
rect 19484 15036 19490 15048
rect 20070 15036 20076 15048
rect 20128 15036 20134 15088
rect 20254 15036 20260 15088
rect 20312 15076 20318 15088
rect 21450 15076 21456 15088
rect 20312 15048 21456 15076
rect 20312 15036 20318 15048
rect 21450 15036 21456 15048
rect 21508 15076 21514 15088
rect 22097 15079 22155 15085
rect 22097 15076 22109 15079
rect 21508 15048 22109 15076
rect 21508 15036 21514 15048
rect 22097 15045 22109 15048
rect 22143 15045 22155 15079
rect 22097 15039 22155 15045
rect 18555 14980 18736 15008
rect 19153 15011 19211 15017
rect 18555 14977 18567 14980
rect 18509 14971 18567 14977
rect 19153 14977 19165 15011
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 19242 14968 19248 15020
rect 19300 15008 19306 15020
rect 19337 15011 19395 15017
rect 19337 15008 19349 15011
rect 19300 14980 19349 15008
rect 19300 14968 19306 14980
rect 19337 14977 19349 14980
rect 19383 15008 19395 15011
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 19383 14980 20453 15008
rect 19383 14977 19395 14980
rect 19337 14971 19395 14977
rect 20441 14977 20453 14980
rect 20487 15008 20499 15011
rect 20530 15008 20536 15020
rect 20487 14980 20536 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 20530 14968 20536 14980
rect 20588 14968 20594 15020
rect 20809 15011 20867 15017
rect 20809 14977 20821 15011
rect 20855 15008 20867 15011
rect 21358 15008 21364 15020
rect 20855 14980 21364 15008
rect 20855 14977 20867 14980
rect 20809 14971 20867 14977
rect 21358 14968 21364 14980
rect 21416 14968 21422 15020
rect 22112 15008 22140 15039
rect 22186 15036 22192 15088
rect 22244 15076 22250 15088
rect 23768 15076 23796 15104
rect 22244 15048 23796 15076
rect 22244 15036 22250 15048
rect 25130 15036 25136 15088
rect 25188 15076 25194 15088
rect 25593 15079 25651 15085
rect 25593 15076 25605 15079
rect 25188 15048 25605 15076
rect 25188 15036 25194 15048
rect 25593 15045 25605 15048
rect 25639 15045 25651 15079
rect 25593 15039 25651 15045
rect 25700 15048 26464 15076
rect 23290 15008 23296 15020
rect 22112 14980 23296 15008
rect 23290 14968 23296 14980
rect 23348 15008 23354 15020
rect 24026 15008 24032 15020
rect 23348 14980 24032 15008
rect 23348 14968 23354 14980
rect 24026 14968 24032 14980
rect 24084 14968 24090 15020
rect 25038 14968 25044 15020
rect 25096 15008 25102 15020
rect 25225 15011 25283 15017
rect 25225 15008 25237 15011
rect 25096 14980 25237 15008
rect 25096 14968 25102 14980
rect 25225 14977 25237 14980
rect 25271 14977 25283 15011
rect 25225 14971 25283 14977
rect 25317 15011 25375 15017
rect 25317 14977 25329 15011
rect 25363 14977 25375 15011
rect 25317 14971 25375 14977
rect 18601 14943 18659 14949
rect 18601 14909 18613 14943
rect 18647 14909 18659 14943
rect 18601 14903 18659 14909
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 18785 14943 18843 14949
rect 18785 14909 18797 14943
rect 18831 14940 18843 14943
rect 19610 14940 19616 14952
rect 18831 14912 19616 14940
rect 18831 14909 18843 14912
rect 18785 14903 18843 14909
rect 18138 14832 18144 14884
rect 18196 14872 18202 14884
rect 18616 14872 18644 14903
rect 18196 14844 18644 14872
rect 18708 14872 18736 14903
rect 19610 14900 19616 14912
rect 19668 14900 19674 14952
rect 19153 14875 19211 14881
rect 19153 14872 19165 14875
rect 18708 14844 19165 14872
rect 18196 14832 18202 14844
rect 18708 14804 18736 14844
rect 19153 14841 19165 14844
rect 19199 14841 19211 14875
rect 19153 14835 19211 14841
rect 18064 14776 18736 14804
rect 19168 14804 19196 14835
rect 19334 14832 19340 14884
rect 19392 14872 19398 14884
rect 21545 14875 21603 14881
rect 21545 14872 21557 14875
rect 19392 14844 21557 14872
rect 19392 14832 19398 14844
rect 21545 14841 21557 14844
rect 21591 14841 21603 14875
rect 25240 14872 25268 14971
rect 25332 14940 25360 14971
rect 25498 14968 25504 15020
rect 25556 14968 25562 15020
rect 25700 15017 25728 15048
rect 25685 15011 25743 15017
rect 25685 14977 25697 15011
rect 25731 14977 25743 15011
rect 25685 14971 25743 14977
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 14977 26019 15011
rect 25961 14971 26019 14977
rect 25976 14940 26004 14971
rect 26050 14968 26056 15020
rect 26108 14968 26114 15020
rect 26237 15011 26295 15017
rect 26237 15008 26249 15011
rect 26160 14980 26249 15008
rect 26160 14952 26188 14980
rect 26237 14977 26249 14980
rect 26283 14977 26295 15011
rect 26237 14971 26295 14977
rect 26326 14968 26332 15020
rect 26384 14968 26390 15020
rect 26436 15017 26464 15048
rect 27080 15048 27936 15076
rect 27080 15020 27108 15048
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 14977 26479 15011
rect 26421 14971 26479 14977
rect 25332 14912 25636 14940
rect 25608 14884 25636 14912
rect 25700 14912 26004 14940
rect 25406 14872 25412 14884
rect 25240 14844 25412 14872
rect 21545 14835 21603 14841
rect 25406 14832 25412 14844
rect 25464 14832 25470 14884
rect 25590 14832 25596 14884
rect 25648 14832 25654 14884
rect 25700 14816 25728 14912
rect 26142 14900 26148 14952
rect 26200 14900 26206 14952
rect 26436 14940 26464 14971
rect 27062 14968 27068 15020
rect 27120 14968 27126 15020
rect 27908 15017 27936 15048
rect 28184 15048 28580 15076
rect 27801 15011 27859 15017
rect 27801 14977 27813 15011
rect 27847 14977 27859 15011
rect 27801 14971 27859 14977
rect 27893 15011 27951 15017
rect 27893 14977 27905 15011
rect 27939 14977 27951 15011
rect 27893 14971 27951 14977
rect 26344 14912 26464 14940
rect 25869 14875 25927 14881
rect 25869 14841 25881 14875
rect 25915 14872 25927 14875
rect 26234 14872 26240 14884
rect 25915 14844 26240 14872
rect 25915 14841 25927 14844
rect 25869 14835 25927 14841
rect 26234 14832 26240 14844
rect 26292 14832 26298 14884
rect 26344 14816 26372 14912
rect 27154 14900 27160 14952
rect 27212 14940 27218 14952
rect 27816 14940 27844 14971
rect 27982 14968 27988 15020
rect 28040 15008 28046 15020
rect 28184 15017 28212 15048
rect 28552 15020 28580 15048
rect 28077 15011 28135 15017
rect 28077 15008 28089 15011
rect 28040 14980 28089 15008
rect 28040 14968 28046 14980
rect 28077 14977 28089 14980
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 28169 15011 28227 15017
rect 28169 14977 28181 15011
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28261 15011 28319 15017
rect 28261 14977 28273 15011
rect 28307 14977 28319 15011
rect 28261 14971 28319 14977
rect 27212 14912 27844 14940
rect 28092 14940 28120 14971
rect 28276 14940 28304 14971
rect 28534 14968 28540 15020
rect 28592 14968 28598 15020
rect 29840 15008 29868 15107
rect 30190 15036 30196 15088
rect 30248 15076 30254 15088
rect 30285 15079 30343 15085
rect 30285 15076 30297 15079
rect 30248 15048 30297 15076
rect 30248 15036 30254 15048
rect 30285 15045 30297 15048
rect 30331 15045 30343 15079
rect 30285 15039 30343 15045
rect 30926 15036 30932 15088
rect 30984 15036 30990 15088
rect 30009 15011 30067 15017
rect 30009 15008 30021 15011
rect 29840 14980 30021 15008
rect 30009 14977 30021 14980
rect 30055 14977 30067 15011
rect 30009 14971 30067 14977
rect 28092 14912 28304 14940
rect 30024 14940 30052 14971
rect 32766 14940 32772 14952
rect 30024 14912 32772 14940
rect 27212 14900 27218 14912
rect 32766 14900 32772 14912
rect 32824 14900 32830 14952
rect 19426 14804 19432 14816
rect 19168 14776 19432 14804
rect 19426 14764 19432 14776
rect 19484 14764 19490 14816
rect 20070 14764 20076 14816
rect 20128 14764 20134 14816
rect 25682 14764 25688 14816
rect 25740 14764 25746 14816
rect 26326 14764 26332 14816
rect 26384 14764 26390 14816
rect 31754 14764 31760 14816
rect 31812 14764 31818 14816
rect 1104 14714 35248 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 35248 14714
rect 1104 14640 35248 14662
rect 3234 14560 3240 14612
rect 3292 14560 3298 14612
rect 3602 14560 3608 14612
rect 3660 14560 3666 14612
rect 3786 14560 3792 14612
rect 3844 14600 3850 14612
rect 4617 14603 4675 14609
rect 4617 14600 4629 14603
rect 3844 14572 4629 14600
rect 3844 14560 3850 14572
rect 4617 14569 4629 14572
rect 4663 14569 4675 14603
rect 4617 14563 4675 14569
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 1857 14467 1915 14473
rect 1857 14464 1869 14467
rect 1544 14436 1869 14464
rect 1544 14424 1550 14436
rect 1857 14433 1869 14436
rect 1903 14433 1915 14467
rect 1857 14427 1915 14433
rect 2866 14424 2872 14476
rect 2924 14464 2930 14476
rect 3252 14464 3280 14560
rect 4249 14467 4307 14473
rect 4249 14464 4261 14467
rect 2924 14436 4261 14464
rect 2924 14424 2930 14436
rect 3988 14405 4016 14436
rect 4249 14433 4261 14436
rect 4295 14433 4307 14467
rect 4249 14427 4307 14433
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 4632 14396 4660 14563
rect 5166 14560 5172 14612
rect 5224 14560 5230 14612
rect 8294 14560 8300 14612
rect 8352 14560 8358 14612
rect 10873 14603 10931 14609
rect 10873 14569 10885 14603
rect 10919 14600 10931 14603
rect 10962 14600 10968 14612
rect 10919 14572 10968 14600
rect 10919 14569 10931 14572
rect 10873 14563 10931 14569
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11606 14560 11612 14612
rect 11664 14560 11670 14612
rect 15657 14603 15715 14609
rect 15657 14569 15669 14603
rect 15703 14600 15715 14603
rect 15930 14600 15936 14612
rect 15703 14572 15936 14600
rect 15703 14569 15715 14572
rect 15657 14563 15715 14569
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 16117 14603 16175 14609
rect 16117 14569 16129 14603
rect 16163 14600 16175 14603
rect 16206 14600 16212 14612
rect 16163 14572 16212 14600
rect 16163 14569 16175 14572
rect 16117 14563 16175 14569
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 16669 14603 16727 14609
rect 16669 14569 16681 14603
rect 16715 14569 16727 14603
rect 16669 14563 16727 14569
rect 5184 14464 5212 14560
rect 6457 14467 6515 14473
rect 6457 14464 6469 14467
rect 5184 14436 6469 14464
rect 6457 14433 6469 14436
rect 6503 14433 6515 14467
rect 6457 14427 6515 14433
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9640 14436 9689 14464
rect 9640 14424 9646 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 10980 14464 11008 14560
rect 10980 14436 11192 14464
rect 9677 14427 9735 14433
rect 6178 14396 6184 14408
rect 4632 14368 6184 14396
rect 3973 14359 4031 14365
rect 6178 14356 6184 14368
rect 6236 14356 6242 14408
rect 7466 14356 7472 14408
rect 7524 14396 7530 14408
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 7524 14368 7590 14396
rect 10520 14368 10977 14396
rect 7524 14356 7530 14368
rect 1486 14288 1492 14340
rect 1544 14328 1550 14340
rect 2133 14331 2191 14337
rect 2133 14328 2145 14331
rect 1544 14300 2145 14328
rect 1544 14288 1550 14300
rect 2133 14297 2145 14300
rect 2179 14297 2191 14331
rect 3881 14331 3939 14337
rect 3881 14328 3893 14331
rect 3358 14300 3893 14328
rect 2133 14291 2191 14297
rect 3881 14297 3893 14300
rect 3927 14297 3939 14331
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 3881 14291 3939 14297
rect 7944 14300 8953 14328
rect 7944 14269 7972 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 10520 14272 10548 14368
rect 10965 14365 10977 14368
rect 11011 14396 11023 14399
rect 11054 14396 11060 14408
rect 11011 14368 11060 14396
rect 11011 14365 11023 14368
rect 10965 14359 11023 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11164 14405 11192 14436
rect 11624 14405 11652 14560
rect 16684 14532 16712 14563
rect 17218 14560 17224 14612
rect 17276 14600 17282 14612
rect 17586 14600 17592 14612
rect 17276 14572 17592 14600
rect 17276 14560 17282 14572
rect 17586 14560 17592 14572
rect 17644 14600 17650 14612
rect 17681 14603 17739 14609
rect 17681 14600 17693 14603
rect 17644 14572 17693 14600
rect 17644 14560 17650 14572
rect 17681 14569 17693 14572
rect 17727 14569 17739 14603
rect 17681 14563 17739 14569
rect 18138 14560 18144 14612
rect 18196 14560 18202 14612
rect 19610 14560 19616 14612
rect 19668 14600 19674 14612
rect 20438 14600 20444 14612
rect 19668 14572 20444 14600
rect 19668 14560 19674 14572
rect 20438 14560 20444 14572
rect 20496 14560 20502 14612
rect 20990 14560 20996 14612
rect 21048 14560 21054 14612
rect 25038 14560 25044 14612
rect 25096 14600 25102 14612
rect 25225 14603 25283 14609
rect 25225 14600 25237 14603
rect 25096 14572 25237 14600
rect 25096 14560 25102 14572
rect 25225 14569 25237 14572
rect 25271 14569 25283 14603
rect 25225 14563 25283 14569
rect 25406 14560 25412 14612
rect 25464 14560 25470 14612
rect 30650 14560 30656 14612
rect 30708 14560 30714 14612
rect 30926 14560 30932 14612
rect 30984 14560 30990 14612
rect 16758 14532 16764 14544
rect 15580 14504 16764 14532
rect 14366 14464 14372 14476
rect 13004 14436 14372 14464
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14365 12127 14399
rect 12069 14359 12127 14365
rect 11333 14331 11391 14337
rect 11333 14297 11345 14331
rect 11379 14328 11391 14331
rect 11882 14328 11888 14340
rect 11379 14300 11888 14328
rect 11379 14297 11391 14300
rect 11333 14291 11391 14297
rect 11882 14288 11888 14300
rect 11940 14328 11946 14340
rect 12084 14328 12112 14359
rect 11940 14300 12112 14328
rect 13004 14314 13032 14436
rect 14366 14424 14372 14436
rect 14424 14464 14430 14476
rect 15194 14464 15200 14476
rect 14424 14436 15200 14464
rect 14424 14424 14430 14436
rect 15194 14424 15200 14436
rect 15252 14464 15258 14476
rect 15580 14473 15608 14504
rect 16758 14492 16764 14504
rect 16816 14492 16822 14544
rect 19797 14535 19855 14541
rect 19797 14501 19809 14535
rect 19843 14532 19855 14535
rect 20901 14535 20959 14541
rect 20901 14532 20913 14535
rect 19843 14504 20913 14532
rect 19843 14501 19855 14504
rect 19797 14495 19855 14501
rect 20901 14501 20913 14504
rect 20947 14501 20959 14535
rect 20901 14495 20959 14501
rect 21450 14492 21456 14544
rect 21508 14492 21514 14544
rect 25682 14492 25688 14544
rect 25740 14532 25746 14544
rect 27525 14535 27583 14541
rect 27525 14532 27537 14535
rect 25740 14504 27537 14532
rect 25740 14492 25746 14504
rect 27525 14501 27537 14504
rect 27571 14501 27583 14535
rect 27525 14495 27583 14501
rect 15565 14467 15623 14473
rect 15565 14464 15577 14467
rect 15252 14436 15577 14464
rect 15252 14424 15258 14436
rect 15565 14433 15577 14436
rect 15611 14433 15623 14467
rect 15565 14427 15623 14433
rect 16209 14467 16267 14473
rect 16209 14433 16221 14467
rect 16255 14464 16267 14467
rect 17494 14464 17500 14476
rect 16255 14436 17500 14464
rect 16255 14433 16267 14436
rect 16209 14427 16267 14433
rect 17494 14424 17500 14436
rect 17552 14464 17558 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 17552 14436 18429 14464
rect 17552 14424 17558 14436
rect 18417 14433 18429 14436
rect 18463 14464 18475 14467
rect 18690 14464 18696 14476
rect 18463 14436 18696 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 18690 14424 18696 14436
rect 18748 14424 18754 14476
rect 18877 14467 18935 14473
rect 18877 14433 18889 14467
rect 18923 14464 18935 14467
rect 20070 14464 20076 14476
rect 18923 14436 20076 14464
rect 18923 14433 18935 14436
rect 18877 14427 18935 14433
rect 14918 14356 14924 14408
rect 14976 14405 14982 14408
rect 15654 14405 15660 14408
rect 14976 14396 14985 14405
rect 15105 14399 15163 14405
rect 14976 14368 15021 14396
rect 14976 14359 14985 14368
rect 15105 14365 15117 14399
rect 15151 14396 15163 14399
rect 15651 14396 15660 14405
rect 15151 14368 15660 14396
rect 15151 14365 15163 14368
rect 15105 14359 15163 14365
rect 15651 14359 15660 14368
rect 14976 14356 14982 14359
rect 15654 14356 15660 14359
rect 15712 14356 15718 14408
rect 15746 14356 15752 14408
rect 15804 14396 15810 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15804 14368 15853 14396
rect 15804 14356 15810 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15841 14359 15899 14365
rect 15930 14356 15936 14408
rect 15988 14396 15994 14408
rect 15988 14368 16436 14396
rect 15988 14356 15994 14368
rect 11940 14288 11946 14300
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 15948 14328 15976 14356
rect 15620 14300 15976 14328
rect 15620 14288 15626 14300
rect 16022 14288 16028 14340
rect 16080 14328 16086 14340
rect 16301 14331 16359 14337
rect 16301 14328 16313 14331
rect 16080 14300 16313 14328
rect 16080 14288 16086 14300
rect 16301 14297 16313 14300
rect 16347 14297 16359 14331
rect 16408 14328 16436 14368
rect 16666 14356 16672 14408
rect 16724 14356 16730 14408
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14396 16819 14399
rect 17678 14396 17684 14408
rect 16807 14368 17684 14396
rect 16807 14365 16819 14368
rect 16761 14359 16819 14365
rect 16776 14328 16804 14359
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 17954 14356 17960 14408
rect 18012 14356 18018 14408
rect 18138 14356 18144 14408
rect 18196 14356 18202 14408
rect 18230 14356 18236 14408
rect 18288 14396 18294 14408
rect 18325 14399 18383 14405
rect 18325 14396 18337 14399
rect 18288 14368 18337 14396
rect 18288 14356 18294 14368
rect 18325 14365 18337 14368
rect 18371 14365 18383 14399
rect 18325 14359 18383 14365
rect 18506 14356 18512 14408
rect 18564 14356 18570 14408
rect 19242 14356 19248 14408
rect 19300 14356 19306 14408
rect 19996 14405 20024 14436
rect 20070 14424 20076 14436
rect 20128 14424 20134 14476
rect 22005 14467 22063 14473
rect 22005 14433 22017 14467
rect 22051 14464 22063 14467
rect 22051 14436 22416 14464
rect 22051 14433 22063 14436
rect 22005 14427 22063 14433
rect 19981 14399 20039 14405
rect 19981 14365 19993 14399
rect 20027 14396 20039 14399
rect 20027 14368 20061 14396
rect 20027 14365 20039 14368
rect 19981 14359 20039 14365
rect 20162 14356 20168 14408
rect 20220 14356 20226 14408
rect 20254 14356 20260 14408
rect 20312 14356 20318 14408
rect 20346 14356 20352 14408
rect 20404 14356 20410 14408
rect 20530 14356 20536 14408
rect 20588 14356 20594 14408
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14396 20775 14399
rect 20809 14399 20867 14405
rect 20809 14396 20821 14399
rect 20763 14368 20821 14396
rect 20763 14365 20775 14368
rect 20717 14359 20775 14365
rect 20809 14365 20821 14368
rect 20855 14365 20867 14399
rect 20809 14359 20867 14365
rect 21358 14356 21364 14408
rect 21416 14396 21422 14408
rect 21729 14399 21787 14405
rect 21729 14396 21741 14399
rect 21416 14368 21741 14396
rect 21416 14356 21422 14368
rect 21729 14365 21741 14368
rect 21775 14365 21787 14399
rect 21729 14359 21787 14365
rect 21818 14356 21824 14408
rect 21876 14356 21882 14408
rect 22388 14405 22416 14436
rect 22462 14424 22468 14476
rect 22520 14424 22526 14476
rect 23201 14467 23259 14473
rect 23201 14433 23213 14467
rect 23247 14464 23259 14467
rect 24857 14467 24915 14473
rect 24857 14464 24869 14467
rect 23247 14436 24869 14464
rect 23247 14433 23259 14436
rect 23201 14427 23259 14433
rect 24857 14433 24869 14436
rect 24903 14464 24915 14467
rect 25498 14464 25504 14476
rect 24903 14436 25504 14464
rect 24903 14433 24915 14436
rect 24857 14427 24915 14433
rect 25498 14424 25504 14436
rect 25556 14464 25562 14476
rect 26142 14464 26148 14476
rect 25556 14436 26148 14464
rect 25556 14424 25562 14436
rect 26142 14424 26148 14436
rect 26200 14464 26206 14476
rect 26200 14436 26832 14464
rect 26200 14424 26206 14436
rect 22373 14399 22431 14405
rect 22373 14365 22385 14399
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 23382 14356 23388 14408
rect 23440 14356 23446 14408
rect 23477 14399 23535 14405
rect 23477 14365 23489 14399
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 23661 14399 23719 14405
rect 23661 14365 23673 14399
rect 23707 14396 23719 14399
rect 23753 14399 23811 14405
rect 23753 14396 23765 14399
rect 23707 14368 23765 14396
rect 23707 14365 23719 14368
rect 23661 14359 23719 14365
rect 23753 14365 23765 14368
rect 23799 14365 23811 14399
rect 23753 14359 23811 14365
rect 16408 14300 16804 14328
rect 16301 14291 16359 14297
rect 16942 14288 16948 14340
rect 17000 14288 17006 14340
rect 18046 14328 18052 14340
rect 17328 14300 18052 14328
rect 7929 14263 7987 14269
rect 7929 14229 7941 14263
rect 7975 14229 7987 14263
rect 7929 14223 7987 14229
rect 10502 14220 10508 14272
rect 10560 14220 10566 14272
rect 15010 14220 15016 14272
rect 15068 14220 15074 14272
rect 15289 14263 15347 14269
rect 15289 14229 15301 14263
rect 15335 14260 15347 14263
rect 15378 14260 15384 14272
rect 15335 14232 15384 14260
rect 15335 14229 15347 14232
rect 15289 14223 15347 14229
rect 15378 14220 15384 14232
rect 15436 14260 15442 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15436 14232 15945 14260
rect 15436 14220 15442 14232
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 15933 14223 15991 14229
rect 16482 14220 16488 14272
rect 16540 14220 16546 14272
rect 16574 14220 16580 14272
rect 16632 14260 16638 14272
rect 17328 14269 17356 14300
rect 18046 14288 18052 14300
rect 18104 14328 18110 14340
rect 18524 14328 18552 14356
rect 18104 14300 18552 14328
rect 18104 14288 18110 14300
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 19613 14331 19671 14337
rect 19613 14328 19625 14331
rect 19484 14300 19625 14328
rect 19484 14288 19490 14300
rect 19613 14297 19625 14300
rect 19659 14297 19671 14331
rect 19613 14291 19671 14297
rect 21082 14288 21088 14340
rect 21140 14288 21146 14340
rect 21836 14328 21864 14356
rect 22738 14328 22744 14340
rect 21836 14300 22744 14328
rect 22738 14288 22744 14300
rect 22796 14328 22802 14340
rect 23492 14328 23520 14359
rect 25130 14356 25136 14408
rect 25188 14356 25194 14408
rect 25590 14356 25596 14408
rect 25648 14356 25654 14408
rect 26050 14356 26056 14408
rect 26108 14356 26114 14408
rect 26329 14399 26387 14405
rect 26329 14396 26341 14399
rect 26160 14368 26341 14396
rect 22796 14300 23520 14328
rect 25148 14328 25176 14356
rect 26160 14328 26188 14368
rect 26329 14365 26341 14368
rect 26375 14396 26387 14399
rect 26418 14396 26424 14408
rect 26375 14368 26424 14396
rect 26375 14365 26387 14368
rect 26329 14359 26387 14365
rect 26418 14356 26424 14368
rect 26476 14356 26482 14408
rect 26804 14405 26832 14436
rect 27154 14424 27160 14476
rect 27212 14424 27218 14476
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14365 26847 14399
rect 30668 14396 30696 14560
rect 34057 14467 34115 14473
rect 34057 14433 34069 14467
rect 34103 14433 34115 14467
rect 34057 14427 34115 14433
rect 30837 14399 30895 14405
rect 30837 14396 30849 14399
rect 30668 14368 30849 14396
rect 26789 14359 26847 14365
rect 30837 14365 30849 14368
rect 30883 14365 30895 14399
rect 30837 14359 30895 14365
rect 25148 14300 26188 14328
rect 34072 14328 34100 14427
rect 34517 14399 34575 14405
rect 34517 14365 34529 14399
rect 34563 14396 34575 14399
rect 34563 14368 35296 14396
rect 34563 14365 34575 14368
rect 34517 14359 34575 14365
rect 34606 14328 34612 14340
rect 34072 14300 34612 14328
rect 22796 14288 22802 14300
rect 34606 14288 34612 14300
rect 34664 14288 34670 14340
rect 17313 14263 17371 14269
rect 17313 14260 17325 14263
rect 16632 14232 17325 14260
rect 16632 14220 16638 14232
rect 17313 14229 17325 14232
rect 17359 14229 17371 14263
rect 17313 14223 17371 14229
rect 21266 14220 21272 14272
rect 21324 14260 21330 14272
rect 21637 14263 21695 14269
rect 21637 14260 21649 14263
rect 21324 14232 21649 14260
rect 21324 14220 21330 14232
rect 21637 14229 21649 14232
rect 21683 14229 21695 14263
rect 21637 14223 21695 14229
rect 23474 14220 23480 14272
rect 23532 14260 23538 14272
rect 23937 14263 23995 14269
rect 23937 14260 23949 14263
rect 23532 14232 23949 14260
rect 23532 14220 23538 14232
rect 23937 14229 23949 14232
rect 23983 14260 23995 14263
rect 24670 14260 24676 14272
rect 23983 14232 24676 14260
rect 23983 14229 23995 14232
rect 23937 14223 23995 14229
rect 24670 14220 24676 14232
rect 24728 14220 24734 14272
rect 25222 14220 25228 14272
rect 25280 14220 25286 14272
rect 1104 14170 35236 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 35236 14170
rect 1104 14096 35236 14118
rect 2314 14016 2320 14068
rect 2372 14016 2378 14068
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8720 14028 9045 14056
rect 8720 14016 8726 14028
rect 9033 14025 9045 14028
rect 9079 14056 9091 14059
rect 11057 14059 11115 14065
rect 11057 14056 11069 14059
rect 9079 14028 11069 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 11057 14025 11069 14028
rect 11103 14025 11115 14059
rect 11057 14019 11115 14025
rect 11606 14016 11612 14068
rect 11664 14016 11670 14068
rect 14918 14016 14924 14068
rect 14976 14016 14982 14068
rect 15562 14016 15568 14068
rect 15620 14016 15626 14068
rect 15654 14016 15660 14068
rect 15712 14016 15718 14068
rect 16206 14016 16212 14068
rect 16264 14056 16270 14068
rect 16301 14059 16359 14065
rect 16301 14056 16313 14059
rect 16264 14028 16313 14056
rect 16264 14016 16270 14028
rect 16301 14025 16313 14028
rect 16347 14025 16359 14059
rect 16301 14019 16359 14025
rect 16482 14016 16488 14068
rect 16540 14016 16546 14068
rect 16758 14016 16764 14068
rect 16816 14016 16822 14068
rect 16850 14016 16856 14068
rect 16908 14056 16914 14068
rect 16945 14059 17003 14065
rect 16945 14056 16957 14059
rect 16908 14028 16957 14056
rect 16908 14016 16914 14028
rect 16945 14025 16957 14028
rect 16991 14025 17003 14059
rect 16945 14019 17003 14025
rect 17310 14016 17316 14068
rect 17368 14056 17374 14068
rect 17589 14059 17647 14065
rect 17589 14056 17601 14059
rect 17368 14028 17601 14056
rect 17368 14016 17374 14028
rect 17589 14025 17601 14028
rect 17635 14056 17647 14059
rect 17954 14056 17960 14068
rect 17635 14028 17960 14056
rect 17635 14025 17647 14028
rect 17589 14019 17647 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 18230 14016 18236 14068
rect 18288 14056 18294 14068
rect 19518 14056 19524 14068
rect 18288 14028 19524 14056
rect 18288 14016 18294 14028
rect 19518 14016 19524 14028
rect 19576 14056 19582 14068
rect 19797 14059 19855 14065
rect 19797 14056 19809 14059
rect 19576 14028 19809 14056
rect 19576 14016 19582 14028
rect 19797 14025 19809 14028
rect 19843 14025 19855 14059
rect 19797 14019 19855 14025
rect 19981 14059 20039 14065
rect 19981 14025 19993 14059
rect 20027 14025 20039 14059
rect 19981 14019 20039 14025
rect 20073 14059 20131 14065
rect 20073 14025 20085 14059
rect 20119 14056 20131 14059
rect 20162 14056 20168 14068
rect 20119 14028 20168 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 5460 13960 6653 13988
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13920 2283 13923
rect 2271 13892 2820 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 2792 13725 2820 13892
rect 3142 13880 3148 13932
rect 3200 13920 3206 13932
rect 3970 13920 3976 13932
rect 3200 13892 3976 13920
rect 3200 13880 3206 13892
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 4065 13855 4123 13861
rect 4065 13821 4077 13855
rect 4111 13852 4123 13855
rect 4614 13852 4620 13864
rect 4111 13824 4620 13852
rect 4111 13821 4123 13824
rect 4065 13815 4123 13821
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 5460 13852 5488 13960
rect 6641 13957 6653 13960
rect 6687 13957 6699 13991
rect 8297 13991 8355 13997
rect 8297 13988 8309 13991
rect 7866 13960 8309 13988
rect 6641 13951 6699 13957
rect 8297 13957 8309 13960
rect 8343 13957 8355 13991
rect 8297 13951 8355 13957
rect 6178 13880 6184 13932
rect 6236 13920 6242 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 6236 13892 6377 13920
rect 6236 13880 6242 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 8389 13923 8447 13929
rect 8389 13889 8401 13923
rect 8435 13920 8447 13923
rect 8754 13920 8760 13932
rect 8435 13892 8760 13920
rect 8435 13889 8447 13892
rect 8389 13883 8447 13889
rect 8754 13880 8760 13892
rect 8812 13880 8818 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 11624 13920 11652 14016
rect 14936 13988 14964 14016
rect 15580 13988 15608 14016
rect 14844 13960 15608 13988
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11624 13892 11805 13920
rect 10137 13883 10195 13889
rect 11793 13889 11805 13892
rect 11839 13889 11851 13923
rect 11793 13883 11851 13889
rect 4724 13824 5488 13852
rect 8113 13855 8171 13861
rect 4341 13787 4399 13793
rect 4341 13753 4353 13787
rect 4387 13784 4399 13787
rect 4724 13784 4752 13824
rect 8113 13821 8125 13855
rect 8159 13852 8171 13855
rect 10152 13852 10180 13883
rect 11882 13880 11888 13932
rect 11940 13920 11946 13932
rect 12069 13923 12127 13929
rect 12069 13920 12081 13923
rect 11940 13892 12081 13920
rect 11940 13880 11946 13892
rect 12069 13889 12081 13892
rect 12115 13889 12127 13923
rect 12069 13883 12127 13889
rect 12989 13923 13047 13929
rect 12989 13889 13001 13923
rect 13035 13920 13047 13923
rect 13630 13920 13636 13932
rect 13035 13892 13636 13920
rect 13035 13889 13047 13892
rect 12989 13883 13047 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 13906 13880 13912 13932
rect 13964 13920 13970 13932
rect 14844 13929 14872 13960
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 13964 13892 14657 13920
rect 13964 13880 13970 13892
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13920 14979 13923
rect 15672 13920 15700 14016
rect 14967 13892 15700 13920
rect 16117 13923 16175 13929
rect 14967 13889 14979 13892
rect 14921 13883 14979 13889
rect 16117 13889 16129 13923
rect 16163 13889 16175 13923
rect 16117 13883 16175 13889
rect 16393 13923 16451 13929
rect 16393 13889 16405 13923
rect 16439 13920 16451 13923
rect 16500 13920 16528 14016
rect 17972 13988 18000 14016
rect 18325 13991 18383 13997
rect 18325 13988 18337 13991
rect 16439 13892 16528 13920
rect 16592 13960 16785 13988
rect 17972 13960 18337 13988
rect 16439 13889 16451 13892
rect 16393 13883 16451 13889
rect 8159 13824 10180 13852
rect 10689 13855 10747 13861
rect 8159 13821 8171 13824
rect 8113 13815 8171 13821
rect 10689 13821 10701 13855
rect 10735 13852 10747 13855
rect 11514 13852 11520 13864
rect 10735 13824 11520 13852
rect 10735 13821 10747 13824
rect 10689 13815 10747 13821
rect 11514 13812 11520 13824
rect 11572 13812 11578 13864
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 13081 13855 13139 13861
rect 13081 13852 13093 13855
rect 12667 13824 13093 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 13081 13821 13093 13824
rect 13127 13852 13139 13855
rect 14550 13852 14556 13864
rect 13127 13824 14556 13852
rect 13127 13821 13139 13824
rect 13081 13815 13139 13821
rect 14550 13812 14556 13824
rect 14608 13812 14614 13864
rect 14660 13852 14688 13883
rect 16132 13852 16160 13883
rect 16592 13864 16620 13960
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16574 13852 16580 13864
rect 14660 13824 16580 13852
rect 16574 13812 16580 13824
rect 16632 13812 16638 13864
rect 4387 13756 4752 13784
rect 13357 13787 13415 13793
rect 4387 13753 4399 13756
rect 4341 13747 4399 13753
rect 13357 13753 13369 13787
rect 13403 13784 13415 13787
rect 14182 13784 14188 13796
rect 13403 13756 14188 13784
rect 13403 13753 13415 13756
rect 13357 13747 13415 13753
rect 14182 13744 14188 13756
rect 14240 13744 14246 13796
rect 15010 13744 15016 13796
rect 15068 13784 15074 13796
rect 16684 13784 16712 13883
rect 16757 13852 16785 13960
rect 18325 13957 18337 13960
rect 18371 13988 18383 13991
rect 18414 13988 18420 14000
rect 18371 13960 18420 13988
rect 18371 13957 18383 13960
rect 18325 13951 18383 13957
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 19337 13991 19395 13997
rect 19337 13957 19349 13991
rect 19383 13988 19395 13991
rect 19996 13988 20024 14019
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20809 14059 20867 14065
rect 20809 14056 20821 14059
rect 20404 14028 20821 14056
rect 20404 14016 20410 14028
rect 20809 14025 20821 14028
rect 20855 14025 20867 14059
rect 20809 14019 20867 14025
rect 21634 14016 21640 14068
rect 21692 14056 21698 14068
rect 22186 14056 22192 14068
rect 21692 14028 22192 14056
rect 21692 14016 21698 14028
rect 22186 14016 22192 14028
rect 22244 14016 22250 14068
rect 22278 14016 22284 14068
rect 22336 14016 22342 14068
rect 22462 14016 22468 14068
rect 22520 14016 22526 14068
rect 23106 14016 23112 14068
rect 23164 14016 23170 14068
rect 24857 14059 24915 14065
rect 24857 14025 24869 14059
rect 24903 14056 24915 14059
rect 24946 14056 24952 14068
rect 24903 14028 24952 14056
rect 24903 14025 24915 14028
rect 24857 14019 24915 14025
rect 24946 14016 24952 14028
rect 25004 14056 25010 14068
rect 25517 14059 25575 14065
rect 25517 14056 25529 14059
rect 25004 14028 25529 14056
rect 25004 14016 25010 14028
rect 25517 14025 25529 14028
rect 25563 14025 25575 14059
rect 25517 14019 25575 14025
rect 25682 14016 25688 14068
rect 25740 14016 25746 14068
rect 31938 14016 31944 14068
rect 31996 14016 32002 14068
rect 34885 14059 34943 14065
rect 34885 14025 34897 14059
rect 34931 14056 34943 14059
rect 35268 14056 35296 14368
rect 34931 14028 35296 14056
rect 34931 14025 34943 14028
rect 34885 14019 34943 14025
rect 20272 13988 20300 14016
rect 19383 13960 19564 13988
rect 19996 13960 20300 13988
rect 19383 13957 19395 13960
rect 19337 13951 19395 13957
rect 16942 13880 16948 13932
rect 17000 13920 17006 13932
rect 17037 13923 17095 13929
rect 17037 13920 17049 13923
rect 17000 13892 17049 13920
rect 17000 13880 17006 13892
rect 17037 13889 17049 13892
rect 17083 13889 17095 13923
rect 18432 13920 18460 13948
rect 19426 13920 19432 13932
rect 18432 13892 19432 13920
rect 17037 13883 17095 13889
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 19536 13920 19564 13960
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 20717 13991 20775 13997
rect 20717 13988 20729 13991
rect 20588 13960 20729 13988
rect 20588 13948 20594 13960
rect 20717 13957 20729 13960
rect 20763 13988 20775 13991
rect 21545 13991 21603 13997
rect 21545 13988 21557 13991
rect 20763 13960 21557 13988
rect 20763 13957 20775 13960
rect 20717 13951 20775 13957
rect 21545 13957 21557 13960
rect 21591 13957 21603 13991
rect 21545 13951 21603 13957
rect 22097 13991 22155 13997
rect 22097 13957 22109 13991
rect 22143 13988 22155 13991
rect 22143 13960 22600 13988
rect 22143 13957 22155 13960
rect 22097 13951 22155 13957
rect 22572 13932 22600 13960
rect 24118 13948 24124 14000
rect 24176 13988 24182 14000
rect 24176 13960 24992 13988
rect 24176 13948 24182 13960
rect 21266 13920 21272 13932
rect 19536 13892 20116 13920
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 16757 13824 16865 13852
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 18785 13855 18843 13861
rect 18785 13821 18797 13855
rect 18831 13852 18843 13855
rect 19536 13852 19564 13892
rect 20088 13864 20116 13892
rect 20272 13892 21272 13920
rect 20272 13864 20300 13892
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 22278 13880 22284 13932
rect 22336 13880 22342 13932
rect 22554 13880 22560 13932
rect 22612 13880 22618 13932
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13889 23811 13923
rect 23753 13883 23811 13889
rect 18831 13824 19564 13852
rect 18831 13821 18843 13824
rect 18785 13815 18843 13821
rect 20070 13812 20076 13864
rect 20128 13812 20134 13864
rect 20254 13812 20260 13864
rect 20312 13812 20318 13864
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20438 13852 20444 13864
rect 20395 13824 20444 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20438 13812 20444 13824
rect 20496 13852 20502 13864
rect 22296 13852 22324 13880
rect 22741 13855 22799 13861
rect 22741 13852 22753 13855
rect 20496 13824 20944 13852
rect 20496 13812 20502 13824
rect 20916 13793 20944 13824
rect 22066 13824 22753 13852
rect 15068 13756 16712 13784
rect 20901 13787 20959 13793
rect 15068 13744 15074 13756
rect 20901 13753 20913 13787
rect 20947 13753 20959 13787
rect 20901 13747 20959 13753
rect 21910 13744 21916 13796
rect 21968 13744 21974 13796
rect 2777 13719 2835 13725
rect 2777 13685 2789 13719
rect 2823 13716 2835 13719
rect 3234 13716 3240 13728
rect 2823 13688 3240 13716
rect 2823 13685 2835 13688
rect 2777 13679 2835 13685
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 4062 13676 4068 13728
rect 4120 13716 4126 13728
rect 4801 13719 4859 13725
rect 4801 13716 4813 13719
rect 4120 13688 4813 13716
rect 4120 13676 4126 13688
rect 4801 13685 4813 13688
rect 4847 13716 4859 13719
rect 4890 13716 4896 13728
rect 4847 13688 4896 13716
rect 4847 13685 4859 13688
rect 4801 13679 4859 13685
rect 4890 13676 4896 13688
rect 4948 13676 4954 13728
rect 8754 13676 8760 13728
rect 8812 13676 8818 13728
rect 12342 13676 12348 13728
rect 12400 13716 12406 13728
rect 14642 13716 14648 13728
rect 12400 13688 14648 13716
rect 12400 13676 12406 13688
rect 14642 13676 14648 13688
rect 14700 13676 14706 13728
rect 14734 13676 14740 13728
rect 14792 13676 14798 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 16117 13719 16175 13725
rect 16117 13716 16129 13719
rect 15252 13688 16129 13716
rect 15252 13676 15258 13688
rect 16117 13685 16129 13688
rect 16163 13685 16175 13719
rect 16117 13679 16175 13685
rect 19150 13676 19156 13728
rect 19208 13716 19214 13728
rect 19797 13719 19855 13725
rect 19797 13716 19809 13719
rect 19208 13688 19809 13716
rect 19208 13676 19214 13688
rect 19797 13685 19809 13688
rect 19843 13685 19855 13719
rect 19797 13679 19855 13685
rect 20346 13676 20352 13728
rect 20404 13716 20410 13728
rect 22066 13716 22094 13824
rect 22741 13821 22753 13824
rect 22787 13852 22799 13855
rect 23658 13852 23664 13864
rect 22787 13824 23664 13852
rect 22787 13821 22799 13824
rect 22741 13815 22799 13821
rect 23658 13812 23664 13824
rect 23716 13852 23722 13864
rect 23768 13852 23796 13883
rect 23934 13880 23940 13932
rect 23992 13880 23998 13932
rect 24670 13880 24676 13932
rect 24728 13880 24734 13932
rect 24964 13920 24992 13960
rect 25038 13948 25044 14000
rect 25096 13988 25102 14000
rect 25317 13991 25375 13997
rect 25317 13988 25329 13991
rect 25096 13960 25329 13988
rect 25096 13948 25102 13960
rect 25317 13957 25329 13960
rect 25363 13957 25375 13991
rect 25317 13951 25375 13957
rect 34146 13948 34152 14000
rect 34204 13948 34210 14000
rect 27798 13920 27804 13932
rect 24964 13892 27804 13920
rect 27798 13880 27804 13892
rect 27856 13920 27862 13932
rect 28353 13923 28411 13929
rect 28353 13920 28365 13923
rect 27856 13892 28365 13920
rect 27856 13880 27862 13892
rect 28353 13889 28365 13892
rect 28399 13889 28411 13923
rect 28353 13883 28411 13889
rect 28460 13892 29868 13920
rect 23716 13824 23796 13852
rect 23716 13812 23722 13824
rect 24486 13812 24492 13864
rect 24544 13812 24550 13864
rect 24688 13852 24716 13880
rect 24688 13824 27936 13852
rect 27908 13784 27936 13824
rect 27982 13812 27988 13864
rect 28040 13852 28046 13864
rect 28261 13855 28319 13861
rect 28261 13852 28273 13855
rect 28040 13824 28273 13852
rect 28040 13812 28046 13824
rect 28261 13821 28273 13824
rect 28307 13821 28319 13855
rect 28460 13852 28488 13892
rect 29840 13864 29868 13892
rect 31570 13880 31576 13932
rect 31628 13880 31634 13932
rect 32309 13923 32367 13929
rect 32309 13920 32321 13923
rect 31772 13892 32321 13920
rect 28261 13815 28319 13821
rect 28368 13824 28488 13852
rect 28721 13855 28779 13861
rect 28368 13784 28396 13824
rect 28721 13821 28733 13855
rect 28767 13852 28779 13855
rect 28767 13824 29132 13852
rect 28767 13821 28779 13824
rect 28721 13815 28779 13821
rect 27908 13756 28396 13784
rect 29104 13728 29132 13824
rect 29822 13812 29828 13864
rect 29880 13812 29886 13864
rect 31478 13812 31484 13864
rect 31536 13852 31542 13864
rect 31665 13855 31723 13861
rect 31665 13852 31677 13855
rect 31536 13824 31677 13852
rect 31536 13812 31542 13824
rect 31665 13821 31677 13824
rect 31711 13821 31723 13855
rect 31665 13815 31723 13821
rect 31772 13728 31800 13892
rect 32309 13889 32321 13892
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 32214 13812 32220 13864
rect 32272 13812 32278 13864
rect 32766 13812 32772 13864
rect 32824 13852 32830 13864
rect 32953 13855 33011 13861
rect 32953 13852 32965 13855
rect 32824 13824 32965 13852
rect 32824 13812 32830 13824
rect 32953 13821 32965 13824
rect 32999 13852 33011 13855
rect 33137 13855 33195 13861
rect 33137 13852 33149 13855
rect 32999 13824 33149 13852
rect 32999 13821 33011 13824
rect 32953 13815 33011 13821
rect 33137 13821 33149 13824
rect 33183 13821 33195 13855
rect 33413 13855 33471 13861
rect 33413 13852 33425 13855
rect 33137 13815 33195 13821
rect 33244 13824 33425 13852
rect 32677 13787 32735 13793
rect 32677 13753 32689 13787
rect 32723 13784 32735 13787
rect 33244 13784 33272 13824
rect 33413 13821 33425 13824
rect 33459 13821 33471 13855
rect 33413 13815 33471 13821
rect 32723 13756 33272 13784
rect 32723 13753 32735 13756
rect 32677 13747 32735 13753
rect 20404 13688 22094 13716
rect 20404 13676 20410 13688
rect 22554 13676 22560 13728
rect 22612 13716 22618 13728
rect 23382 13716 23388 13728
rect 22612 13688 23388 13716
rect 22612 13676 22618 13688
rect 23382 13676 23388 13688
rect 23440 13716 23446 13728
rect 23477 13719 23535 13725
rect 23477 13716 23489 13719
rect 23440 13688 23489 13716
rect 23440 13676 23446 13688
rect 23477 13685 23489 13688
rect 23523 13685 23535 13719
rect 23477 13679 23535 13685
rect 25222 13676 25228 13728
rect 25280 13716 25286 13728
rect 25501 13719 25559 13725
rect 25501 13716 25513 13719
rect 25280 13688 25513 13716
rect 25280 13676 25286 13688
rect 25501 13685 25513 13688
rect 25547 13685 25559 13719
rect 25501 13679 25559 13685
rect 29086 13676 29092 13728
rect 29144 13676 29150 13728
rect 31665 13719 31723 13725
rect 31665 13685 31677 13719
rect 31711 13716 31723 13719
rect 31754 13716 31760 13728
rect 31711 13688 31760 13716
rect 31711 13685 31723 13688
rect 31665 13679 31723 13685
rect 31754 13676 31760 13688
rect 31812 13676 31818 13728
rect 1104 13626 35248 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 35248 13626
rect 1104 13552 35248 13574
rect 4249 13515 4307 13521
rect 4249 13481 4261 13515
rect 4295 13512 4307 13515
rect 4614 13512 4620 13524
rect 4295 13484 4620 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4724 13484 5948 13512
rect 4724 13444 4752 13484
rect 4264 13416 4752 13444
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 1452 13348 3556 13376
rect 1452 13336 1458 13348
rect 1670 13200 1676 13252
rect 1728 13200 1734 13252
rect 2406 13200 2412 13252
rect 2464 13200 2470 13252
rect 3142 13132 3148 13184
rect 3200 13132 3206 13184
rect 3528 13181 3556 13348
rect 4264 13320 4292 13416
rect 4632 13385 4660 13416
rect 4798 13404 4804 13456
rect 4856 13404 4862 13456
rect 4890 13404 4896 13456
rect 4948 13404 4954 13456
rect 4525 13379 4583 13385
rect 4525 13376 4537 13379
rect 4356 13348 4537 13376
rect 4356 13320 4384 13348
rect 4525 13345 4537 13348
rect 4571 13345 4583 13379
rect 4525 13339 4583 13345
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13345 4675 13379
rect 4816 13376 4844 13404
rect 4617 13339 4675 13345
rect 4724 13348 4844 13376
rect 4908 13376 4936 13404
rect 5629 13379 5687 13385
rect 4908 13348 5212 13376
rect 4246 13268 4252 13320
rect 4304 13268 4310 13320
rect 4338 13268 4344 13320
rect 4396 13268 4402 13320
rect 4724 13317 4752 13348
rect 4908 13317 4936 13348
rect 5184 13320 5212 13348
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 5813 13379 5871 13385
rect 5813 13376 5825 13379
rect 5675 13348 5825 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 5813 13345 5825 13348
rect 5859 13345 5871 13379
rect 5813 13339 5871 13345
rect 4433 13311 4491 13317
rect 4433 13277 4445 13311
rect 4479 13277 4491 13311
rect 4433 13271 4491 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 4893 13311 4951 13317
rect 4893 13277 4905 13311
rect 4939 13277 4951 13311
rect 4893 13271 4951 13277
rect 4985 13311 5043 13317
rect 4985 13277 4997 13311
rect 5031 13302 5043 13311
rect 5074 13302 5080 13320
rect 5031 13277 5080 13302
rect 4985 13274 5080 13277
rect 4985 13271 5043 13274
rect 3602 13200 3608 13252
rect 3660 13240 3666 13252
rect 4062 13240 4068 13252
rect 3660 13212 4068 13240
rect 3660 13200 3666 13212
rect 4062 13200 4068 13212
rect 4120 13200 4126 13252
rect 3513 13175 3571 13181
rect 3513 13141 3525 13175
rect 3559 13172 3571 13175
rect 3878 13172 3884 13184
rect 3559 13144 3884 13172
rect 3559 13141 3571 13144
rect 3513 13135 3571 13141
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 4356 13172 4384 13268
rect 4448 13240 4476 13271
rect 5074 13268 5080 13274
rect 5132 13268 5138 13320
rect 5166 13268 5172 13320
rect 5224 13268 5230 13320
rect 5258 13268 5264 13320
rect 5316 13268 5322 13320
rect 5350 13268 5356 13320
rect 5408 13268 5414 13320
rect 5920 13317 5948 13484
rect 14642 13472 14648 13524
rect 14700 13472 14706 13524
rect 14734 13472 14740 13524
rect 14792 13512 14798 13524
rect 14829 13515 14887 13521
rect 14829 13512 14841 13515
rect 14792 13484 14841 13512
rect 14792 13472 14798 13484
rect 14829 13481 14841 13484
rect 14875 13481 14887 13515
rect 14829 13475 14887 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 16114 13512 16120 13524
rect 15795 13484 16120 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16390 13472 16396 13524
rect 16448 13472 16454 13524
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 16942 13512 16948 13524
rect 16623 13484 16948 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17034 13472 17040 13524
rect 17092 13472 17098 13524
rect 17586 13472 17592 13524
rect 17644 13512 17650 13524
rect 18141 13515 18199 13521
rect 18141 13512 18153 13515
rect 17644 13484 18153 13512
rect 17644 13472 17650 13484
rect 18141 13481 18153 13484
rect 18187 13512 18199 13515
rect 18230 13512 18236 13524
rect 18187 13484 18236 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 18230 13472 18236 13484
rect 18288 13472 18294 13524
rect 18877 13515 18935 13521
rect 18877 13481 18889 13515
rect 18923 13512 18935 13515
rect 19242 13512 19248 13524
rect 18923 13484 19248 13512
rect 18923 13481 18935 13484
rect 18877 13475 18935 13481
rect 19242 13472 19248 13484
rect 19300 13472 19306 13524
rect 19518 13472 19524 13524
rect 19576 13472 19582 13524
rect 20438 13472 20444 13524
rect 20496 13512 20502 13524
rect 20533 13515 20591 13521
rect 20533 13512 20545 13515
rect 20496 13484 20545 13512
rect 20496 13472 20502 13484
rect 20533 13481 20545 13484
rect 20579 13512 20591 13515
rect 20990 13512 20996 13524
rect 20579 13484 20996 13512
rect 20579 13481 20591 13484
rect 20533 13475 20591 13481
rect 20990 13472 20996 13484
rect 21048 13512 21054 13524
rect 21269 13515 21327 13521
rect 21269 13512 21281 13515
rect 21048 13484 21281 13512
rect 21048 13472 21054 13484
rect 21269 13481 21281 13484
rect 21315 13481 21327 13515
rect 21269 13475 21327 13481
rect 21634 13472 21640 13524
rect 21692 13472 21698 13524
rect 21910 13512 21916 13524
rect 21836 13484 21916 13512
rect 14660 13444 14688 13472
rect 15930 13444 15936 13456
rect 14660 13416 15936 13444
rect 15930 13404 15936 13416
rect 15988 13404 15994 13456
rect 17052 13444 17080 13472
rect 17052 13416 17172 13444
rect 6273 13379 6331 13385
rect 6273 13345 6285 13379
rect 6319 13376 6331 13379
rect 9217 13379 9275 13385
rect 9217 13376 9229 13379
rect 6319 13348 9229 13376
rect 6319 13345 6331 13348
rect 6273 13339 6331 13345
rect 9217 13345 9229 13348
rect 9263 13345 9275 13379
rect 9217 13339 9275 13345
rect 10689 13379 10747 13385
rect 10689 13345 10701 13379
rect 10735 13345 10747 13379
rect 10689 13339 10747 13345
rect 11885 13379 11943 13385
rect 11885 13345 11897 13379
rect 11931 13376 11943 13379
rect 12158 13376 12164 13388
rect 11931 13348 12164 13376
rect 11931 13345 11943 13348
rect 11885 13339 11943 13345
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 8662 13268 8668 13320
rect 8720 13308 8726 13320
rect 8938 13308 8944 13320
rect 8720 13280 8944 13308
rect 8720 13268 8726 13280
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 10704 13308 10732 13339
rect 12158 13336 12164 13348
rect 12216 13376 12222 13388
rect 15378 13376 15384 13388
rect 12216 13348 12572 13376
rect 12216 13336 12222 13348
rect 10873 13311 10931 13317
rect 10873 13308 10885 13311
rect 10704 13280 10885 13308
rect 10873 13277 10885 13280
rect 10919 13277 10931 13311
rect 10873 13271 10931 13277
rect 11422 13268 11428 13320
rect 11480 13308 11486 13320
rect 12253 13311 12311 13317
rect 12253 13308 12265 13311
rect 11480 13280 12265 13308
rect 11480 13268 11486 13280
rect 12253 13277 12265 13280
rect 12299 13277 12311 13311
rect 12253 13271 12311 13277
rect 12345 13311 12403 13317
rect 12345 13277 12357 13311
rect 12391 13308 12403 13311
rect 12434 13308 12440 13320
rect 12391 13280 12440 13308
rect 12391 13277 12403 13280
rect 12345 13271 12403 13277
rect 4614 13240 4620 13252
rect 4448 13212 4620 13240
rect 4614 13200 4620 13212
rect 4672 13200 4678 13252
rect 9674 13200 9680 13252
rect 9732 13200 9738 13252
rect 12268 13240 12296 13271
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12544 13317 12572 13348
rect 15028 13348 15384 13376
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13277 12587 13311
rect 12529 13271 12587 13277
rect 14550 13268 14556 13320
rect 14608 13268 14614 13320
rect 14642 13268 14648 13320
rect 14700 13317 14706 13320
rect 15028 13317 15056 13348
rect 15378 13336 15384 13348
rect 15436 13376 15442 13388
rect 17037 13379 17095 13385
rect 17037 13376 17049 13379
rect 15436 13348 16804 13376
rect 15436 13336 15442 13348
rect 14700 13311 14749 13317
rect 14700 13277 14703 13311
rect 14737 13277 14749 13311
rect 14700 13271 14749 13277
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13277 15071 13311
rect 15013 13271 15071 13277
rect 14700 13268 14706 13271
rect 15194 13268 15200 13320
rect 15252 13268 15258 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 15565 13311 15623 13317
rect 15565 13277 15577 13311
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 14921 13243 14979 13249
rect 12268 13212 13124 13240
rect 13096 13184 13124 13212
rect 14921 13209 14933 13243
rect 14967 13240 14979 13243
rect 15580 13240 15608 13271
rect 16574 13268 16580 13320
rect 16632 13268 16638 13320
rect 16776 13317 16804 13348
rect 16868 13348 17049 13376
rect 16868 13317 16896 13348
rect 17037 13345 17049 13348
rect 17083 13345 17095 13379
rect 17037 13339 17095 13345
rect 17144 13320 17172 13416
rect 19426 13404 19432 13456
rect 19484 13444 19490 13456
rect 20456 13444 20484 13472
rect 19484 13416 20484 13444
rect 19484 13404 19490 13416
rect 17862 13336 17868 13388
rect 17920 13376 17926 13388
rect 17920 13348 18828 13376
rect 17920 13336 17926 13348
rect 16761 13311 16819 13317
rect 16761 13277 16773 13311
rect 16807 13277 16819 13311
rect 16761 13271 16819 13277
rect 16849 13311 16907 13317
rect 16849 13277 16861 13311
rect 16895 13277 16907 13311
rect 16849 13271 16907 13277
rect 16942 13268 16948 13320
rect 17000 13268 17006 13320
rect 17126 13268 17132 13320
rect 17184 13268 17190 13320
rect 18046 13268 18052 13320
rect 18104 13268 18110 13320
rect 18230 13268 18236 13320
rect 18288 13308 18294 13320
rect 18325 13311 18383 13317
rect 18325 13308 18337 13311
rect 18288 13280 18337 13308
rect 18288 13268 18294 13280
rect 18325 13277 18337 13280
rect 18371 13277 18383 13311
rect 18325 13271 18383 13277
rect 18414 13268 18420 13320
rect 18472 13308 18478 13320
rect 18601 13311 18659 13317
rect 18601 13308 18613 13311
rect 18472 13280 18613 13308
rect 18472 13268 18478 13280
rect 18601 13277 18613 13280
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 18693 13311 18751 13317
rect 18693 13277 18705 13311
rect 18739 13277 18751 13311
rect 18800 13308 18828 13348
rect 19150 13336 19156 13388
rect 19208 13376 19214 13388
rect 21836 13385 21864 13484
rect 21910 13472 21916 13484
rect 21968 13512 21974 13524
rect 22646 13512 22652 13524
rect 21968 13484 22652 13512
rect 21968 13472 21974 13484
rect 22646 13472 22652 13484
rect 22704 13512 22710 13524
rect 23017 13515 23075 13521
rect 23017 13512 23029 13515
rect 22704 13484 23029 13512
rect 22704 13472 22710 13484
rect 23017 13481 23029 13484
rect 23063 13512 23075 13515
rect 23106 13512 23112 13524
rect 23063 13484 23112 13512
rect 23063 13481 23075 13484
rect 23017 13475 23075 13481
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 23658 13472 23664 13524
rect 23716 13472 23722 13524
rect 27246 13472 27252 13524
rect 27304 13472 27310 13524
rect 28534 13472 28540 13524
rect 28592 13472 28598 13524
rect 31478 13472 31484 13524
rect 31536 13472 31542 13524
rect 31941 13515 31999 13521
rect 31941 13481 31953 13515
rect 31987 13512 31999 13515
rect 32214 13512 32220 13524
rect 31987 13484 32220 13512
rect 31987 13481 31999 13484
rect 31941 13475 31999 13481
rect 32214 13472 32220 13484
rect 32272 13472 32278 13524
rect 34146 13472 34152 13524
rect 34204 13472 34210 13524
rect 22002 13404 22008 13456
rect 22060 13444 22066 13456
rect 22189 13447 22247 13453
rect 22189 13444 22201 13447
rect 22060 13416 22201 13444
rect 22060 13404 22066 13416
rect 22189 13413 22201 13416
rect 22235 13444 22247 13447
rect 24486 13444 24492 13456
rect 22235 13416 24492 13444
rect 22235 13413 22247 13416
rect 22189 13407 22247 13413
rect 24486 13404 24492 13416
rect 24544 13404 24550 13456
rect 21821 13379 21879 13385
rect 21821 13376 21833 13379
rect 19208 13348 21833 13376
rect 19208 13336 19214 13348
rect 21821 13345 21833 13348
rect 21867 13345 21879 13379
rect 21821 13339 21879 13345
rect 29086 13336 29092 13388
rect 29144 13336 29150 13388
rect 29362 13336 29368 13388
rect 29420 13336 29426 13388
rect 19889 13311 19947 13317
rect 19889 13308 19901 13311
rect 18800 13280 19901 13308
rect 18693 13271 18751 13277
rect 19889 13277 19901 13280
rect 19935 13308 19947 13311
rect 20530 13308 20536 13320
rect 19935 13280 20536 13308
rect 19935 13277 19947 13280
rect 19889 13271 19947 13277
rect 14967 13212 15608 13240
rect 18064 13240 18092 13268
rect 18506 13240 18512 13252
rect 18064 13212 18512 13240
rect 14967 13209 14979 13212
rect 14921 13203 14979 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 18708 13240 18736 13271
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20901 13311 20959 13317
rect 20901 13277 20913 13311
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 19334 13240 19340 13252
rect 18708 13212 19340 13240
rect 5258 13172 5264 13184
rect 4356 13144 5264 13172
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 17034 13172 17040 13184
rect 13136 13144 17040 13172
rect 13136 13132 13142 13144
rect 17034 13132 17040 13144
rect 17092 13172 17098 13184
rect 17589 13175 17647 13181
rect 17589 13172 17601 13175
rect 17092 13144 17601 13172
rect 17092 13132 17098 13144
rect 17589 13141 17601 13144
rect 17635 13172 17647 13175
rect 18138 13172 18144 13184
rect 17635 13144 18144 13172
rect 17635 13141 17647 13144
rect 17589 13135 17647 13141
rect 18138 13132 18144 13144
rect 18196 13172 18202 13184
rect 18708 13172 18736 13212
rect 19334 13200 19340 13212
rect 19392 13240 19398 13252
rect 20254 13240 20260 13252
rect 19392 13212 20260 13240
rect 19392 13200 19398 13212
rect 20254 13200 20260 13212
rect 20312 13240 20318 13252
rect 20916 13240 20944 13271
rect 21358 13268 21364 13320
rect 21416 13308 21422 13320
rect 22005 13311 22063 13317
rect 22005 13308 22017 13311
rect 21416 13280 22017 13308
rect 21416 13268 21422 13280
rect 22005 13277 22017 13280
rect 22051 13308 22063 13311
rect 23566 13308 23572 13320
rect 22051 13280 23572 13308
rect 22051 13277 22063 13280
rect 22005 13271 22063 13277
rect 23566 13268 23572 13280
rect 23624 13268 23630 13320
rect 27430 13268 27436 13320
rect 27488 13268 27494 13320
rect 27525 13311 27583 13317
rect 27525 13277 27537 13311
rect 27571 13277 27583 13311
rect 27525 13271 27583 13277
rect 27709 13311 27767 13317
rect 27709 13277 27721 13311
rect 27755 13277 27767 13311
rect 27709 13271 27767 13277
rect 23934 13240 23940 13252
rect 20312 13212 20944 13240
rect 23308 13212 23940 13240
rect 20312 13200 20318 13212
rect 23308 13184 23336 13212
rect 23934 13200 23940 13212
rect 23992 13240 23998 13252
rect 24029 13243 24087 13249
rect 24029 13240 24041 13243
rect 23992 13212 24041 13240
rect 23992 13200 23998 13212
rect 24029 13209 24041 13212
rect 24075 13209 24087 13243
rect 27540 13240 27568 13271
rect 24029 13203 24087 13209
rect 27264 13212 27568 13240
rect 27724 13240 27752 13271
rect 27798 13268 27804 13320
rect 27856 13308 27862 13320
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 27856 13280 28089 13308
rect 27856 13268 27862 13280
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 28169 13311 28227 13317
rect 28169 13277 28181 13311
rect 28215 13277 28227 13311
rect 28169 13271 28227 13277
rect 27982 13240 27988 13252
rect 27724 13212 27988 13240
rect 27264 13184 27292 13212
rect 27982 13200 27988 13212
rect 28040 13200 28046 13252
rect 28184 13240 28212 13271
rect 28258 13268 28264 13320
rect 28316 13268 28322 13320
rect 28350 13268 28356 13320
rect 28408 13268 28414 13320
rect 28994 13268 29000 13320
rect 29052 13268 29058 13320
rect 29380 13308 29408 13336
rect 29733 13311 29791 13317
rect 29733 13308 29745 13311
rect 29380 13280 29745 13308
rect 29733 13277 29745 13280
rect 29779 13277 29791 13311
rect 31496 13308 31524 13472
rect 31754 13404 31760 13456
rect 31812 13444 31818 13456
rect 31849 13447 31907 13453
rect 31849 13444 31861 13447
rect 31812 13416 31861 13444
rect 31812 13404 31818 13416
rect 31849 13413 31861 13416
rect 31895 13413 31907 13447
rect 31849 13407 31907 13413
rect 32033 13379 32091 13385
rect 32033 13345 32045 13379
rect 32079 13376 32091 13379
rect 32309 13379 32367 13385
rect 32309 13376 32321 13379
rect 32079 13348 32321 13376
rect 32079 13345 32091 13348
rect 32033 13339 32091 13345
rect 32309 13345 32321 13348
rect 32355 13345 32367 13379
rect 32309 13339 32367 13345
rect 31662 13308 31668 13320
rect 31496 13280 31668 13308
rect 29733 13271 29791 13277
rect 31662 13268 31668 13280
rect 31720 13308 31726 13320
rect 31757 13311 31815 13317
rect 31757 13308 31769 13311
rect 31720 13280 31769 13308
rect 31720 13268 31726 13280
rect 31757 13277 31769 13280
rect 31803 13277 31815 13311
rect 31757 13271 31815 13277
rect 30009 13243 30067 13249
rect 30009 13240 30021 13243
rect 28092 13212 28212 13240
rect 29380 13212 30021 13240
rect 28092 13184 28120 13212
rect 18196 13144 18736 13172
rect 18196 13132 18202 13144
rect 22554 13132 22560 13184
rect 22612 13132 22618 13184
rect 23290 13132 23296 13184
rect 23348 13132 23354 13184
rect 27246 13132 27252 13184
rect 27304 13132 27310 13184
rect 28074 13132 28080 13184
rect 28132 13132 28138 13184
rect 29380 13181 29408 13212
rect 30009 13209 30021 13212
rect 30055 13209 30067 13243
rect 30009 13203 30067 13209
rect 30742 13200 30748 13252
rect 30800 13200 30806 13252
rect 29365 13175 29423 13181
rect 29365 13141 29377 13175
rect 29411 13141 29423 13175
rect 29365 13135 29423 13141
rect 31386 13132 31392 13184
rect 31444 13172 31450 13184
rect 31938 13172 31944 13184
rect 31444 13144 31944 13172
rect 31444 13132 31450 13144
rect 31938 13132 31944 13144
rect 31996 13172 32002 13184
rect 32048 13172 32076 13339
rect 34057 13311 34115 13317
rect 34057 13277 34069 13311
rect 34103 13277 34115 13311
rect 34057 13271 34115 13277
rect 31996 13144 32076 13172
rect 33965 13175 34023 13181
rect 31996 13132 32002 13144
rect 33965 13141 33977 13175
rect 34011 13172 34023 13175
rect 34072 13172 34100 13271
rect 34698 13172 34704 13184
rect 34011 13144 34704 13172
rect 34011 13141 34023 13144
rect 33965 13135 34023 13141
rect 34698 13132 34704 13144
rect 34756 13132 34762 13184
rect 1104 13082 35236 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 35236 13082
rect 1104 13008 35236 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 1670 12968 1676 12980
rect 1627 12940 1676 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 2406 12928 2412 12980
rect 2464 12928 2470 12980
rect 2866 12968 2872 12980
rect 2746 12940 2872 12968
rect 934 12792 940 12844
rect 992 12832 998 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 992 12804 1409 12832
rect 992 12792 998 12804
rect 1397 12801 1409 12804
rect 1443 12801 1455 12835
rect 1397 12795 1455 12801
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2746 12832 2774 12940
rect 2866 12928 2872 12940
rect 2924 12968 2930 12980
rect 3326 12968 3332 12980
rect 2924 12940 3332 12968
rect 2924 12928 2930 12940
rect 3326 12928 3332 12940
rect 3384 12968 3390 12980
rect 3513 12971 3571 12977
rect 3513 12968 3525 12971
rect 3384 12940 3525 12968
rect 3384 12928 3390 12940
rect 3513 12937 3525 12940
rect 3559 12937 3571 12971
rect 3513 12931 3571 12937
rect 3878 12928 3884 12980
rect 3936 12928 3942 12980
rect 5350 12968 5356 12980
rect 4632 12940 5356 12968
rect 3970 12860 3976 12912
rect 4028 12900 4034 12912
rect 4065 12903 4123 12909
rect 4065 12900 4077 12903
rect 4028 12872 4077 12900
rect 4028 12860 4034 12872
rect 4065 12869 4077 12872
rect 4111 12869 4123 12903
rect 4065 12863 4123 12869
rect 4632 12844 4660 12940
rect 5350 12928 5356 12940
rect 5408 12968 5414 12980
rect 6523 12971 6581 12977
rect 6523 12968 6535 12971
rect 5408 12940 6535 12968
rect 5408 12928 5414 12940
rect 6523 12937 6535 12940
rect 6569 12937 6581 12971
rect 6523 12931 6581 12937
rect 8849 12971 8907 12977
rect 8849 12937 8861 12971
rect 8895 12937 8907 12971
rect 8849 12931 8907 12937
rect 5166 12860 5172 12912
rect 5224 12900 5230 12912
rect 5445 12903 5503 12909
rect 5445 12900 5457 12903
rect 5224 12872 5457 12900
rect 5224 12860 5230 12872
rect 5445 12869 5457 12872
rect 5491 12900 5503 12903
rect 6733 12903 6791 12909
rect 6733 12900 6745 12903
rect 5491 12872 6745 12900
rect 5491 12869 5503 12872
rect 5445 12863 5503 12869
rect 6733 12869 6745 12872
rect 6779 12869 6791 12903
rect 7377 12903 7435 12909
rect 7377 12900 7389 12903
rect 6733 12863 6791 12869
rect 6840 12872 7389 12900
rect 2547 12804 2774 12832
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 3142 12792 3148 12844
rect 3200 12832 3206 12844
rect 4246 12832 4252 12844
rect 3200 12804 4252 12832
rect 3200 12792 3206 12804
rect 4246 12792 4252 12804
rect 4304 12792 4310 12844
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12832 4399 12835
rect 4614 12832 4620 12844
rect 4387 12804 4620 12832
rect 4387 12801 4399 12804
rect 4341 12795 4399 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5258 12792 5264 12844
rect 5316 12832 5322 12844
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5316 12804 5825 12832
rect 5316 12792 5322 12804
rect 5813 12801 5825 12804
rect 5859 12801 5871 12835
rect 5813 12795 5871 12801
rect 5905 12767 5963 12773
rect 5905 12733 5917 12767
rect 5951 12733 5963 12767
rect 5905 12727 5963 12733
rect 6181 12767 6239 12773
rect 6181 12733 6193 12767
rect 6227 12764 6239 12767
rect 6840 12764 6868 12872
rect 7377 12869 7389 12872
rect 7423 12869 7435 12903
rect 7377 12863 7435 12869
rect 8386 12860 8392 12912
rect 8444 12860 8450 12912
rect 8864 12900 8892 12931
rect 8938 12928 8944 12980
rect 8996 12968 9002 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 8996 12940 9137 12968
rect 8996 12928 9002 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 9125 12931 9183 12937
rect 9401 12971 9459 12977
rect 9401 12937 9413 12971
rect 9447 12968 9459 12971
rect 9674 12968 9680 12980
rect 9447 12940 9680 12968
rect 9447 12937 9459 12940
rect 9401 12931 9459 12937
rect 9674 12928 9680 12940
rect 9732 12928 9738 12980
rect 12526 12968 12532 12980
rect 12406 12940 12532 12968
rect 8864 12872 10180 12900
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 10152 12841 10180 12872
rect 10502 12860 10508 12912
rect 10560 12860 10566 12912
rect 11333 12903 11391 12909
rect 11333 12869 11345 12903
rect 11379 12900 11391 12903
rect 12406 12900 12434 12940
rect 12526 12928 12532 12940
rect 12584 12928 12590 12980
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12937 14427 12971
rect 14369 12931 14427 12937
rect 11379 12872 12434 12900
rect 13791 12903 13849 12909
rect 11379 12869 11391 12872
rect 11333 12863 11391 12869
rect 9309 12835 9367 12841
rect 9309 12801 9321 12835
rect 9355 12832 9367 12835
rect 10137 12835 10195 12841
rect 9355 12804 9904 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 6227 12736 6868 12764
rect 7101 12767 7159 12773
rect 6227 12733 6239 12736
rect 6181 12727 6239 12733
rect 7101 12733 7113 12767
rect 7147 12764 7159 12767
rect 8956 12764 8984 12792
rect 9582 12764 9588 12776
rect 7147 12736 9588 12764
rect 7147 12733 7159 12736
rect 7101 12727 7159 12733
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 4706 12696 4712 12708
rect 4571 12668 4712 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 4706 12656 4712 12668
rect 4764 12656 4770 12708
rect 5920 12696 5948 12727
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 6365 12699 6423 12705
rect 6365 12696 6377 12699
rect 5920 12668 6377 12696
rect 6365 12665 6377 12668
rect 6411 12665 6423 12699
rect 6365 12659 6423 12665
rect 4062 12588 4068 12640
rect 4120 12628 4126 12640
rect 4157 12631 4215 12637
rect 4157 12628 4169 12631
rect 4120 12600 4169 12628
rect 4120 12588 4126 12600
rect 4157 12597 4169 12600
rect 4203 12628 4215 12631
rect 4338 12628 4344 12640
rect 4203 12600 4344 12628
rect 4203 12597 4215 12600
rect 4157 12591 4215 12597
rect 4338 12588 4344 12600
rect 4396 12588 4402 12640
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 9876 12637 9904 12804
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 11900 12841 11928 12872
rect 13791 12869 13803 12903
rect 13837 12900 13849 12903
rect 14384 12900 14412 12931
rect 14642 12928 14648 12980
rect 14700 12968 14706 12980
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14700 12940 15117 12968
rect 14700 12928 14706 12940
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15105 12931 15163 12937
rect 15286 12928 15292 12980
rect 15344 12928 15350 12980
rect 15930 12928 15936 12980
rect 15988 12928 15994 12980
rect 16301 12971 16359 12977
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 17494 12968 17500 12980
rect 16347 12940 17500 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 17681 12971 17739 12977
rect 17681 12968 17693 12971
rect 17644 12940 17693 12968
rect 17644 12928 17650 12940
rect 17681 12937 17693 12940
rect 17727 12937 17739 12971
rect 17681 12931 17739 12937
rect 18506 12928 18512 12980
rect 18564 12968 18570 12980
rect 19150 12968 19156 12980
rect 18564 12940 19156 12968
rect 18564 12928 18570 12940
rect 19150 12928 19156 12940
rect 19208 12928 19214 12980
rect 19242 12928 19248 12980
rect 19300 12928 19306 12980
rect 19337 12971 19395 12977
rect 19337 12937 19349 12971
rect 19383 12968 19395 12971
rect 19426 12968 19432 12980
rect 19383 12940 19432 12968
rect 19383 12937 19395 12940
rect 19337 12931 19395 12937
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19794 12928 19800 12980
rect 19852 12968 19858 12980
rect 20073 12971 20131 12977
rect 20073 12968 20085 12971
rect 19852 12940 20085 12968
rect 19852 12928 19858 12940
rect 20073 12937 20085 12940
rect 20119 12937 20131 12971
rect 20073 12931 20131 12937
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 21082 12968 21088 12980
rect 20303 12940 21088 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 21358 12928 21364 12980
rect 21416 12968 21422 12980
rect 21453 12971 21511 12977
rect 21453 12968 21465 12971
rect 21416 12940 21465 12968
rect 21416 12928 21422 12940
rect 21453 12937 21465 12940
rect 21499 12937 21511 12971
rect 22738 12968 22744 12980
rect 21453 12931 21511 12937
rect 22204 12940 22744 12968
rect 15304 12900 15332 12928
rect 13837 12872 14412 12900
rect 14660 12872 15332 12900
rect 15948 12900 15976 12928
rect 19260 12900 19288 12928
rect 15948 12872 18092 12900
rect 13837 12869 13849 12872
rect 13791 12863 13849 12869
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 11572 12804 11621 12832
rect 11572 12792 11578 12804
rect 11609 12801 11621 12804
rect 11655 12801 11667 12835
rect 11609 12795 11667 12801
rect 11885 12835 11943 12841
rect 11885 12801 11897 12835
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 12434 12792 12440 12844
rect 12492 12792 12498 12844
rect 13630 12792 13636 12844
rect 13688 12792 13694 12844
rect 13906 12792 13912 12844
rect 13964 12792 13970 12844
rect 14001 12835 14059 12841
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12764 12035 12767
rect 12526 12764 12532 12776
rect 12023 12736 12532 12764
rect 12023 12733 12035 12736
rect 11977 12727 12035 12733
rect 12526 12724 12532 12736
rect 12584 12724 12590 12776
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 13924 12764 13952 12792
rect 13219 12736 13952 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 5132 12600 6561 12628
rect 5132 12588 5138 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 9861 12631 9919 12637
rect 9861 12597 9873 12631
rect 9907 12628 9919 12631
rect 10042 12628 10048 12640
rect 9907 12600 10048 12628
rect 9907 12597 9919 12600
rect 9861 12591 9919 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 14016 12628 14044 12795
rect 14090 12792 14096 12844
rect 14148 12792 14154 12844
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 14660 12832 14688 12872
rect 14323 12804 14688 12832
rect 14737 12835 14795 12841
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 14737 12801 14749 12835
rect 14783 12832 14795 12835
rect 15013 12835 15071 12841
rect 15013 12832 15025 12835
rect 14783 12804 15025 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 15013 12801 15025 12804
rect 15059 12832 15071 12835
rect 15102 12832 15108 12844
rect 15059 12804 15108 12832
rect 15059 12801 15071 12804
rect 15013 12795 15071 12801
rect 15102 12792 15108 12804
rect 15160 12792 15166 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15930 12832 15936 12844
rect 15243 12804 15936 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 14553 12767 14611 12773
rect 14553 12733 14565 12767
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 14458 12656 14464 12708
rect 14516 12696 14522 12708
rect 14568 12696 14596 12727
rect 14642 12724 14648 12776
rect 14700 12724 14706 12776
rect 14826 12724 14832 12776
rect 14884 12724 14890 12776
rect 15746 12724 15752 12776
rect 15804 12764 15810 12776
rect 16132 12764 16160 12795
rect 16390 12792 16396 12844
rect 16448 12792 16454 12844
rect 17034 12792 17040 12844
rect 17092 12792 17098 12844
rect 17310 12792 17316 12844
rect 17368 12792 17374 12844
rect 17862 12792 17868 12844
rect 17920 12792 17926 12844
rect 18064 12841 18092 12872
rect 18524 12872 19288 12900
rect 19444 12900 19472 12928
rect 19705 12903 19763 12909
rect 19705 12900 19717 12903
rect 19444 12872 19717 12900
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18414 12832 18420 12844
rect 18095 12804 18420 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 18524 12841 18552 12872
rect 19705 12869 19717 12872
rect 19751 12869 19763 12903
rect 19705 12863 19763 12869
rect 20990 12860 20996 12912
rect 21048 12860 21054 12912
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12801 18567 12835
rect 18509 12795 18567 12801
rect 18601 12835 18659 12841
rect 18601 12801 18613 12835
rect 18647 12801 18659 12835
rect 18601 12795 18659 12801
rect 18785 12835 18843 12841
rect 18785 12801 18797 12835
rect 18831 12801 18843 12835
rect 18785 12795 18843 12801
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12832 18935 12835
rect 19058 12832 19064 12844
rect 18923 12804 19064 12832
rect 18923 12801 18935 12804
rect 18877 12795 18935 12801
rect 15804 12736 16160 12764
rect 18233 12767 18291 12773
rect 15804 12724 15810 12736
rect 18233 12733 18245 12767
rect 18279 12764 18291 12767
rect 18616 12764 18644 12795
rect 18690 12764 18696 12776
rect 18279 12736 18696 12764
rect 18279 12733 18291 12736
rect 18233 12727 18291 12733
rect 18690 12724 18696 12736
rect 18748 12724 18754 12776
rect 18800 12764 18828 12795
rect 19058 12792 19064 12804
rect 19116 12792 19122 12844
rect 19245 12835 19303 12841
rect 19245 12801 19257 12835
rect 19291 12832 19303 12835
rect 19334 12832 19340 12844
rect 19291 12804 19340 12832
rect 19291 12801 19303 12804
rect 19245 12795 19303 12801
rect 19334 12792 19340 12804
rect 19392 12832 19398 12844
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19392 12804 19901 12832
rect 19392 12792 19398 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 18969 12767 19027 12773
rect 18969 12764 18981 12767
rect 18800 12736 18981 12764
rect 18969 12733 18981 12736
rect 19015 12733 19027 12767
rect 19904 12764 19932 12795
rect 19978 12792 19984 12844
rect 20036 12792 20042 12844
rect 22204 12841 22232 12940
rect 22738 12928 22744 12940
rect 22796 12968 22802 12980
rect 23198 12968 23204 12980
rect 22796 12940 23204 12968
rect 22796 12928 22802 12940
rect 23198 12928 23204 12940
rect 23256 12968 23262 12980
rect 23293 12971 23351 12977
rect 23293 12968 23305 12971
rect 23256 12940 23305 12968
rect 23256 12928 23262 12940
rect 23293 12937 23305 12940
rect 23339 12937 23351 12971
rect 23293 12931 23351 12937
rect 25222 12928 25228 12980
rect 25280 12928 25286 12980
rect 27062 12928 27068 12980
rect 27120 12968 27126 12980
rect 27985 12971 28043 12977
rect 27120 12940 27660 12968
rect 27120 12928 27126 12940
rect 23109 12903 23167 12909
rect 23109 12900 23121 12903
rect 22841 12872 23121 12900
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 20548 12804 22017 12832
rect 20548 12776 20576 12804
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 20530 12764 20536 12776
rect 19904 12736 20536 12764
rect 18969 12727 19027 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 21913 12767 21971 12773
rect 21913 12733 21925 12767
rect 21959 12733 21971 12767
rect 21913 12727 21971 12733
rect 15470 12696 15476 12708
rect 14516 12668 15476 12696
rect 14516 12656 14522 12668
rect 15470 12656 15476 12668
rect 15528 12696 15534 12708
rect 16482 12696 16488 12708
rect 15528 12668 16488 12696
rect 15528 12656 15534 12668
rect 16482 12656 16488 12668
rect 16540 12656 16546 12708
rect 19426 12696 19432 12708
rect 18248 12668 19432 12696
rect 18248 12640 18276 12668
rect 19426 12656 19432 12668
rect 19484 12696 19490 12708
rect 19521 12699 19579 12705
rect 19521 12696 19533 12699
rect 19484 12668 19533 12696
rect 19484 12656 19490 12668
rect 19521 12665 19533 12668
rect 19567 12665 19579 12699
rect 19521 12659 19579 12665
rect 15010 12628 15016 12640
rect 14016 12600 15016 12628
rect 15010 12588 15016 12600
rect 15068 12628 15074 12640
rect 15746 12628 15752 12640
rect 15068 12600 15752 12628
rect 15068 12588 15074 12600
rect 15746 12588 15752 12600
rect 15804 12588 15810 12640
rect 16114 12588 16120 12640
rect 16172 12588 16178 12640
rect 18230 12588 18236 12640
rect 18288 12588 18294 12640
rect 18322 12588 18328 12640
rect 18380 12588 18386 12640
rect 21928 12628 21956 12727
rect 22020 12696 22048 12795
rect 22554 12792 22560 12844
rect 22612 12832 22618 12844
rect 22841 12832 22869 12872
rect 23109 12869 23121 12872
rect 23155 12869 23167 12903
rect 25240 12900 25268 12928
rect 26878 12900 26884 12912
rect 25240 12872 25636 12900
rect 23109 12863 23167 12869
rect 22612 12804 22869 12832
rect 23201 12835 23259 12841
rect 22612 12792 22618 12804
rect 23201 12801 23213 12835
rect 23247 12832 23259 12835
rect 23658 12832 23664 12844
rect 23247 12804 23664 12832
rect 23247 12801 23259 12804
rect 23201 12795 23259 12801
rect 23658 12792 23664 12804
rect 23716 12832 23722 12844
rect 23845 12835 23903 12841
rect 23845 12832 23857 12835
rect 23716 12804 23857 12832
rect 23716 12792 23722 12804
rect 23845 12801 23857 12804
rect 23891 12801 23903 12835
rect 23845 12795 23903 12801
rect 24121 12835 24179 12841
rect 24121 12801 24133 12835
rect 24167 12801 24179 12835
rect 24121 12795 24179 12801
rect 22094 12724 22100 12776
rect 22152 12724 22158 12776
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12764 22431 12767
rect 24136 12764 24164 12795
rect 24486 12792 24492 12844
rect 24544 12792 24550 12844
rect 25038 12792 25044 12844
rect 25096 12792 25102 12844
rect 25608 12841 25636 12872
rect 26528 12872 26884 12900
rect 25225 12835 25283 12841
rect 25225 12801 25237 12835
rect 25271 12801 25283 12835
rect 25225 12795 25283 12801
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 26145 12835 26203 12841
rect 26145 12801 26157 12835
rect 26191 12801 26203 12835
rect 26145 12795 26203 12801
rect 22419 12736 24164 12764
rect 22419 12733 22431 12736
rect 22373 12727 22431 12733
rect 25130 12724 25136 12776
rect 25188 12724 25194 12776
rect 25240 12764 25268 12795
rect 25866 12764 25872 12776
rect 25240 12736 25872 12764
rect 22830 12696 22836 12708
rect 22020 12668 22836 12696
rect 22830 12656 22836 12668
rect 22888 12696 22894 12708
rect 22925 12699 22983 12705
rect 22925 12696 22937 12699
rect 22888 12668 22937 12696
rect 22888 12656 22894 12668
rect 22925 12665 22937 12668
rect 22971 12665 22983 12699
rect 25240 12696 25268 12736
rect 25866 12724 25872 12736
rect 25924 12764 25930 12776
rect 26053 12767 26111 12773
rect 26053 12764 26065 12767
rect 25924 12736 26065 12764
rect 25924 12724 25930 12736
rect 26053 12733 26065 12736
rect 26099 12733 26111 12767
rect 26053 12727 26111 12733
rect 26160 12696 26188 12795
rect 26528 12773 26556 12872
rect 26878 12860 26884 12872
rect 26936 12900 26942 12912
rect 27632 12909 27660 12940
rect 27985 12937 27997 12971
rect 28031 12968 28043 12971
rect 28258 12968 28264 12980
rect 28031 12940 28264 12968
rect 28031 12937 28043 12940
rect 27985 12931 28043 12937
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 28629 12971 28687 12977
rect 28629 12937 28641 12971
rect 28675 12968 28687 12971
rect 28994 12968 29000 12980
rect 28675 12940 29000 12968
rect 28675 12937 28687 12940
rect 28629 12931 28687 12937
rect 28994 12928 29000 12940
rect 29052 12928 29058 12980
rect 29362 12928 29368 12980
rect 29420 12968 29426 12980
rect 29549 12971 29607 12977
rect 29549 12968 29561 12971
rect 29420 12940 29561 12968
rect 29420 12928 29426 12940
rect 29549 12937 29561 12940
rect 29595 12968 29607 12971
rect 29730 12968 29736 12980
rect 29595 12940 29736 12968
rect 29595 12937 29607 12940
rect 29549 12931 29607 12937
rect 29730 12928 29736 12940
rect 29788 12928 29794 12980
rect 30561 12971 30619 12977
rect 30561 12937 30573 12971
rect 30607 12968 30619 12971
rect 30650 12968 30656 12980
rect 30607 12940 30656 12968
rect 30607 12937 30619 12940
rect 30561 12931 30619 12937
rect 30650 12928 30656 12940
rect 30708 12928 30714 12980
rect 30742 12928 30748 12980
rect 30800 12928 30806 12980
rect 31386 12928 31392 12980
rect 31444 12968 31450 12980
rect 31573 12971 31631 12977
rect 31573 12968 31585 12971
rect 31444 12940 31585 12968
rect 31444 12928 31450 12940
rect 31573 12937 31585 12940
rect 31619 12937 31631 12971
rect 31573 12931 31631 12937
rect 27617 12903 27675 12909
rect 26936 12872 27384 12900
rect 26936 12860 26942 12872
rect 27157 12835 27215 12841
rect 27157 12832 27169 12835
rect 26804 12804 27169 12832
rect 26804 12776 26832 12804
rect 27157 12801 27169 12804
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 27246 12792 27252 12844
rect 27304 12792 27310 12844
rect 27356 12841 27384 12872
rect 27617 12869 27629 12903
rect 27663 12869 27675 12903
rect 27617 12863 27675 12869
rect 27706 12860 27712 12912
rect 27764 12900 27770 12912
rect 27817 12903 27875 12909
rect 27817 12900 27829 12903
rect 27764 12872 27829 12900
rect 27764 12860 27770 12872
rect 27817 12869 27829 12872
rect 27863 12869 27875 12903
rect 28276 12900 28304 12928
rect 28276 12872 28488 12900
rect 27817 12863 27875 12869
rect 27341 12835 27399 12841
rect 27341 12801 27353 12835
rect 27387 12801 27399 12835
rect 27341 12795 27399 12801
rect 28261 12835 28319 12841
rect 28261 12801 28273 12835
rect 28307 12801 28319 12835
rect 28261 12795 28319 12801
rect 26513 12767 26571 12773
rect 26513 12733 26525 12767
rect 26559 12733 26571 12767
rect 26513 12727 26571 12733
rect 26786 12724 26792 12776
rect 26844 12724 26850 12776
rect 27065 12767 27123 12773
rect 27065 12733 27077 12767
rect 27111 12733 27123 12767
rect 27065 12727 27123 12733
rect 27525 12767 27583 12773
rect 27525 12733 27537 12767
rect 27571 12764 27583 12767
rect 28074 12764 28080 12776
rect 27571 12736 28080 12764
rect 27571 12733 27583 12736
rect 27525 12727 27583 12733
rect 22925 12659 22983 12665
rect 23492 12668 25268 12696
rect 26068 12668 26188 12696
rect 27080 12696 27108 12727
rect 28074 12724 28080 12736
rect 28132 12764 28138 12776
rect 28276 12764 28304 12795
rect 28132 12736 28304 12764
rect 28132 12724 28138 12736
rect 28350 12724 28356 12776
rect 28408 12724 28414 12776
rect 27614 12696 27620 12708
rect 27080 12668 27620 12696
rect 23492 12640 23520 12668
rect 26068 12640 26096 12668
rect 27614 12656 27620 12668
rect 27672 12656 27678 12708
rect 22186 12628 22192 12640
rect 21928 12600 22192 12628
rect 22186 12588 22192 12600
rect 22244 12588 22250 12640
rect 22646 12588 22652 12640
rect 22704 12628 22710 12640
rect 23382 12628 23388 12640
rect 22704 12600 23388 12628
rect 22704 12588 22710 12600
rect 23382 12588 23388 12600
rect 23440 12588 23446 12640
rect 23474 12588 23480 12640
rect 23532 12588 23538 12640
rect 26050 12588 26056 12640
rect 26108 12588 26114 12640
rect 26694 12588 26700 12640
rect 26752 12628 26758 12640
rect 27246 12628 27252 12640
rect 26752 12600 27252 12628
rect 26752 12588 26758 12600
rect 27246 12588 27252 12600
rect 27304 12628 27310 12640
rect 28460 12637 28488 12872
rect 30668 12841 30696 12928
rect 31662 12860 31668 12912
rect 31720 12900 31726 12912
rect 31720 12872 32352 12900
rect 31720 12860 31726 12872
rect 30653 12835 30711 12841
rect 30653 12801 30665 12835
rect 30699 12801 30711 12835
rect 30653 12795 30711 12801
rect 31754 12792 31760 12844
rect 31812 12792 31818 12844
rect 31938 12792 31944 12844
rect 31996 12792 32002 12844
rect 32324 12841 32352 12872
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12801 32367 12835
rect 32309 12795 32367 12801
rect 31849 12767 31907 12773
rect 31849 12733 31861 12767
rect 31895 12764 31907 12767
rect 32217 12767 32275 12773
rect 32217 12764 32229 12767
rect 31895 12736 32229 12764
rect 31895 12733 31907 12736
rect 31849 12727 31907 12733
rect 32217 12733 32229 12736
rect 32263 12733 32275 12767
rect 32217 12727 32275 12733
rect 32674 12656 32680 12708
rect 32732 12656 32738 12708
rect 27801 12631 27859 12637
rect 27801 12628 27813 12631
rect 27304 12600 27813 12628
rect 27304 12588 27310 12600
rect 27801 12597 27813 12600
rect 27847 12597 27859 12631
rect 27801 12591 27859 12597
rect 28445 12631 28503 12637
rect 28445 12597 28457 12631
rect 28491 12597 28503 12631
rect 28445 12591 28503 12597
rect 34609 12631 34667 12637
rect 34609 12597 34621 12631
rect 34655 12628 34667 12631
rect 34698 12628 34704 12640
rect 34655 12600 34704 12628
rect 34655 12597 34667 12600
rect 34609 12591 34667 12597
rect 34698 12588 34704 12600
rect 34756 12588 34762 12640
rect 1104 12538 35248 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 35248 12538
rect 1104 12464 35248 12486
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 4062 12424 4068 12436
rect 3191 12396 4068 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 8205 12427 8263 12433
rect 8205 12393 8217 12427
rect 8251 12424 8263 12427
rect 8386 12424 8392 12436
rect 8251 12396 8392 12424
rect 8251 12393 8263 12396
rect 8205 12387 8263 12393
rect 8386 12384 8392 12396
rect 8444 12384 8450 12436
rect 8665 12427 8723 12433
rect 8665 12393 8677 12427
rect 8711 12424 8723 12427
rect 8754 12424 8760 12436
rect 8711 12396 8760 12424
rect 8711 12393 8723 12396
rect 8665 12387 8723 12393
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 4249 12359 4307 12365
rect 4249 12356 4261 12359
rect 3384 12328 4261 12356
rect 3384 12316 3390 12328
rect 1394 12248 1400 12300
rect 1452 12248 1458 12300
rect 3436 12229 3464 12328
rect 3988 12229 4016 12328
rect 4249 12325 4261 12328
rect 4295 12325 4307 12359
rect 4249 12319 4307 12325
rect 3421 12223 3479 12229
rect 3421 12189 3433 12223
rect 3467 12189 3479 12223
rect 3421 12183 3479 12189
rect 3973 12223 4031 12229
rect 3973 12189 3985 12223
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 4672 12192 6285 12220
rect 4672 12180 4678 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6273 12183 6331 12189
rect 6886 12192 7021 12220
rect 1670 12112 1676 12164
rect 1728 12112 1734 12164
rect 3329 12155 3387 12161
rect 3329 12152 3341 12155
rect 2898 12124 3341 12152
rect 3329 12121 3341 12124
rect 3375 12121 3387 12155
rect 3329 12115 3387 12121
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 6457 12087 6515 12093
rect 6457 12053 6469 12087
rect 6503 12084 6515 12087
rect 6886 12084 6914 12192
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8680 12220 8708 12387
rect 8754 12384 8760 12396
rect 8812 12424 8818 12436
rect 10042 12424 10048 12436
rect 8812 12396 10048 12424
rect 8812 12384 8818 12396
rect 10042 12384 10048 12396
rect 10100 12384 10106 12436
rect 11514 12384 11520 12436
rect 11572 12384 11578 12436
rect 14090 12384 14096 12436
rect 14148 12384 14154 12436
rect 15102 12424 15108 12436
rect 14200 12396 15108 12424
rect 14200 12288 14228 12396
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 16206 12384 16212 12436
rect 16264 12424 16270 12436
rect 16393 12427 16451 12433
rect 16393 12424 16405 12427
rect 16264 12396 16405 12424
rect 16264 12384 16270 12396
rect 16393 12393 16405 12396
rect 16439 12393 16451 12427
rect 16393 12387 16451 12393
rect 16684 12396 17356 12424
rect 14366 12316 14372 12368
rect 14424 12356 14430 12368
rect 15120 12356 15148 12384
rect 16574 12356 16580 12368
rect 14424 12328 15056 12356
rect 15120 12328 16580 12356
rect 14424 12316 14430 12328
rect 13556 12260 14228 12288
rect 14384 12288 14412 12316
rect 14384 12260 14596 12288
rect 8159 12192 8708 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 12434 12180 12440 12232
rect 12492 12180 12498 12232
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 13556 12138 13584 12260
rect 13906 12180 13912 12232
rect 13964 12220 13970 12232
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 13964 12192 14289 12220
rect 13964 12180 13970 12192
rect 14277 12189 14289 12192
rect 14323 12220 14335 12223
rect 14458 12220 14464 12232
rect 14323 12192 14464 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 14458 12180 14464 12192
rect 14516 12180 14522 12232
rect 14568 12229 14596 12260
rect 14918 12248 14924 12300
rect 14976 12248 14982 12300
rect 15028 12288 15056 12328
rect 16574 12316 16580 12328
rect 16632 12316 16638 12368
rect 15028 12260 15332 12288
rect 14553 12223 14611 12229
rect 14553 12189 14565 12223
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14734 12180 14740 12232
rect 14792 12220 14798 12232
rect 15304 12229 15332 12260
rect 15562 12248 15568 12300
rect 15620 12248 15626 12300
rect 15654 12248 15660 12300
rect 15712 12248 15718 12300
rect 15059 12223 15117 12229
rect 14792 12198 14872 12220
rect 15059 12198 15071 12223
rect 14792 12192 15071 12198
rect 14792 12180 14798 12192
rect 14844 12189 15071 12192
rect 15105 12189 15117 12223
rect 14844 12183 15117 12189
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 15381 12223 15439 12229
rect 15381 12189 15393 12223
rect 15427 12222 15439 12223
rect 15427 12220 15516 12222
rect 15746 12220 15752 12232
rect 15427 12194 15752 12220
rect 15427 12189 15439 12194
rect 15488 12192 15752 12194
rect 15381 12183 15439 12189
rect 14844 12170 15102 12183
rect 15197 12155 15255 12161
rect 15197 12121 15209 12155
rect 15243 12121 15255 12155
rect 15304 12152 15332 12183
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 16684 12229 16712 12396
rect 17328 12356 17356 12396
rect 17494 12384 17500 12436
rect 17552 12384 17558 12436
rect 17954 12384 17960 12436
rect 18012 12424 18018 12436
rect 18141 12427 18199 12433
rect 18141 12424 18153 12427
rect 18012 12396 18153 12424
rect 18012 12384 18018 12396
rect 18141 12393 18153 12396
rect 18187 12393 18199 12427
rect 18141 12387 18199 12393
rect 18414 12384 18420 12436
rect 18472 12424 18478 12436
rect 18472 12396 19334 12424
rect 18472 12384 18478 12396
rect 19306 12356 19334 12396
rect 19978 12384 19984 12436
rect 20036 12424 20042 12436
rect 20073 12427 20131 12433
rect 20073 12424 20085 12427
rect 20036 12396 20085 12424
rect 20036 12384 20042 12396
rect 20073 12393 20085 12396
rect 20119 12424 20131 12427
rect 20257 12427 20315 12433
rect 20257 12424 20269 12427
rect 20119 12396 20269 12424
rect 20119 12393 20131 12396
rect 20073 12387 20131 12393
rect 20257 12393 20269 12396
rect 20303 12424 20315 12427
rect 22281 12427 22339 12433
rect 20303 12396 21864 12424
rect 20303 12393 20315 12396
rect 20257 12387 20315 12393
rect 17328 12328 19012 12356
rect 19306 12328 20116 12356
rect 16868 12260 17080 12288
rect 16868 12232 16896 12260
rect 16025 12223 16083 12229
rect 16025 12220 16037 12223
rect 15988 12192 16037 12220
rect 15988 12180 15994 12192
rect 16025 12189 16037 12192
rect 16071 12189 16083 12223
rect 16669 12223 16727 12229
rect 16025 12183 16083 12189
rect 16580 12201 16638 12207
rect 16580 12167 16592 12201
rect 16626 12167 16638 12201
rect 16669 12189 16681 12223
rect 16715 12189 16727 12223
rect 16669 12183 16727 12189
rect 16850 12180 16856 12232
rect 16908 12180 16914 12232
rect 17052 12229 17080 12260
rect 17954 12248 17960 12300
rect 18012 12288 18018 12300
rect 18984 12288 19012 12328
rect 20088 12300 20116 12328
rect 19794 12288 19800 12300
rect 18012 12260 18644 12288
rect 18012 12248 18018 12260
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 17037 12223 17095 12229
rect 17037 12189 17049 12223
rect 17083 12189 17095 12223
rect 17037 12183 17095 12189
rect 16580 12164 16638 12167
rect 15841 12155 15899 12161
rect 15841 12152 15853 12155
rect 15304 12124 15853 12152
rect 15197 12115 15255 12121
rect 15841 12121 15853 12124
rect 15887 12121 15899 12155
rect 15841 12115 15899 12121
rect 6503 12056 6914 12084
rect 6503 12053 6515 12056
rect 6457 12047 6515 12053
rect 7190 12044 7196 12096
rect 7248 12044 7254 12096
rect 13630 12044 13636 12096
rect 13688 12084 13694 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 13688 12056 14473 12084
rect 13688 12044 13694 12056
rect 14461 12053 14473 12056
rect 14507 12084 14519 12087
rect 15212 12084 15240 12115
rect 16574 12112 16580 12164
rect 16632 12112 16638 12164
rect 16758 12112 16764 12164
rect 16816 12152 16822 12164
rect 16960 12152 16988 12183
rect 17218 12180 17224 12232
rect 17276 12220 17282 12232
rect 17313 12223 17371 12229
rect 17313 12220 17325 12223
rect 17276 12192 17325 12220
rect 17276 12180 17282 12192
rect 17313 12189 17325 12192
rect 17359 12189 17371 12223
rect 17313 12183 17371 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12220 17923 12223
rect 18506 12220 18512 12232
rect 17911 12192 18512 12220
rect 17911 12189 17923 12192
rect 17865 12183 17923 12189
rect 17129 12155 17187 12161
rect 17129 12152 17141 12155
rect 16816 12124 17141 12152
rect 16816 12112 16822 12124
rect 17129 12121 17141 12124
rect 17175 12121 17187 12155
rect 17328 12152 17356 12183
rect 18506 12180 18512 12192
rect 18564 12180 18570 12232
rect 18616 12229 18644 12260
rect 18984 12260 19800 12288
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18690 12180 18696 12232
rect 18748 12180 18754 12232
rect 18984 12229 19012 12260
rect 19794 12248 19800 12260
rect 19852 12248 19858 12300
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 18785 12223 18843 12229
rect 18785 12189 18797 12223
rect 18831 12189 18843 12223
rect 18785 12183 18843 12189
rect 18969 12223 19027 12229
rect 18969 12189 18981 12223
rect 19015 12189 19027 12223
rect 18969 12183 19027 12189
rect 18230 12152 18236 12164
rect 17328 12124 18236 12152
rect 17129 12115 17187 12121
rect 18230 12112 18236 12124
rect 18288 12112 18294 12164
rect 18800 12096 18828 12183
rect 19426 12180 19432 12232
rect 19484 12180 19490 12232
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19981 12223 20039 12229
rect 19981 12189 19993 12223
rect 20027 12220 20039 12223
rect 20088 12220 20116 12248
rect 20027 12192 20116 12220
rect 20257 12223 20315 12229
rect 20027 12189 20039 12192
rect 19981 12183 20039 12189
rect 20257 12189 20269 12223
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 19628 12152 19656 12183
rect 19352 12124 19656 12152
rect 19352 12096 19380 12124
rect 20272 12096 20300 12183
rect 20346 12180 20352 12232
rect 20404 12220 20410 12232
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 20404 12192 21097 12220
rect 20404 12180 20410 12192
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 21177 12223 21235 12229
rect 21177 12189 21189 12223
rect 21223 12220 21235 12223
rect 21453 12223 21511 12229
rect 21453 12220 21465 12223
rect 21223 12192 21465 12220
rect 21223 12189 21235 12192
rect 21177 12183 21235 12189
rect 21453 12189 21465 12192
rect 21499 12189 21511 12223
rect 21453 12183 21511 12189
rect 21637 12223 21695 12229
rect 21637 12189 21649 12223
rect 21683 12220 21695 12223
rect 21726 12220 21732 12232
rect 21683 12192 21732 12220
rect 21683 12189 21695 12192
rect 21637 12183 21695 12189
rect 21726 12180 21732 12192
rect 21784 12180 21790 12232
rect 21836 12229 21864 12396
rect 22281 12393 22293 12427
rect 22327 12424 22339 12427
rect 22830 12424 22836 12436
rect 22327 12396 22836 12424
rect 22327 12393 22339 12396
rect 22281 12387 22339 12393
rect 22830 12384 22836 12396
rect 22888 12424 22894 12436
rect 23290 12424 23296 12436
rect 22888 12396 23296 12424
rect 22888 12384 22894 12396
rect 23290 12384 23296 12396
rect 23348 12384 23354 12436
rect 23382 12384 23388 12436
rect 23440 12424 23446 12436
rect 25041 12427 25099 12433
rect 23440 12396 24716 12424
rect 23440 12384 23446 12396
rect 22741 12359 22799 12365
rect 22741 12325 22753 12359
rect 22787 12356 22799 12359
rect 24581 12359 24639 12365
rect 24581 12356 24593 12359
rect 22787 12328 23336 12356
rect 22787 12325 22799 12328
rect 22741 12319 22799 12325
rect 22020 12260 22968 12288
rect 22020 12232 22048 12260
rect 21821 12223 21879 12229
rect 21821 12189 21833 12223
rect 21867 12189 21879 12223
rect 21821 12183 21879 12189
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22002 12220 22008 12232
rect 21959 12192 22008 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 21836 12152 21864 12183
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 22520 12192 22569 12220
rect 22520 12180 22526 12192
rect 22557 12189 22569 12192
rect 22603 12189 22615 12223
rect 22557 12183 22615 12189
rect 22738 12180 22744 12232
rect 22796 12180 22802 12232
rect 22940 12220 22968 12260
rect 23017 12223 23075 12229
rect 23017 12220 23029 12223
rect 22940 12192 23029 12220
rect 23017 12189 23029 12192
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 23198 12180 23204 12232
rect 23256 12180 23262 12232
rect 22094 12152 22100 12164
rect 21836 12124 22100 12152
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 23109 12155 23167 12161
rect 23109 12121 23121 12155
rect 23155 12121 23167 12155
rect 23308 12152 23336 12328
rect 23860 12328 24593 12356
rect 23860 12300 23888 12328
rect 24581 12325 24593 12328
rect 24627 12325 24639 12359
rect 24581 12319 24639 12325
rect 23842 12248 23848 12300
rect 23900 12248 23906 12300
rect 23382 12180 23388 12232
rect 23440 12180 23446 12232
rect 23477 12223 23535 12229
rect 23477 12189 23489 12223
rect 23523 12220 23535 12223
rect 23569 12223 23627 12229
rect 23569 12220 23581 12223
rect 23523 12192 23581 12220
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 23569 12189 23581 12192
rect 23615 12189 23627 12223
rect 23569 12183 23627 12189
rect 24121 12223 24179 12229
rect 24121 12189 24133 12223
rect 24167 12220 24179 12223
rect 24688 12220 24716 12396
rect 25041 12393 25053 12427
rect 25087 12424 25099 12427
rect 25222 12424 25228 12436
rect 25087 12396 25228 12424
rect 25087 12393 25099 12396
rect 25041 12387 25099 12393
rect 25222 12384 25228 12396
rect 25280 12424 25286 12436
rect 27249 12427 27307 12433
rect 25280 12396 26280 12424
rect 25280 12384 25286 12396
rect 25593 12359 25651 12365
rect 25593 12356 25605 12359
rect 25056 12328 25605 12356
rect 25056 12220 25084 12328
rect 25593 12325 25605 12328
rect 25639 12325 25651 12359
rect 25593 12319 25651 12325
rect 25866 12316 25872 12368
rect 25924 12316 25930 12368
rect 25884 12288 25912 12316
rect 25884 12260 26188 12288
rect 25682 12220 25688 12232
rect 24167 12192 25084 12220
rect 25148 12192 25688 12220
rect 24167 12189 24179 12192
rect 24121 12183 24179 12189
rect 23308 12124 24164 12152
rect 23109 12115 23167 12121
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 14507 12056 18337 12084
rect 14507 12053 14519 12056
rect 14461 12047 14519 12053
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18325 12047 18383 12053
rect 18782 12044 18788 12096
rect 18840 12044 18846 12096
rect 19334 12044 19340 12096
rect 19392 12044 19398 12096
rect 20254 12044 20260 12096
rect 20312 12044 20318 12096
rect 20625 12087 20683 12093
rect 20625 12053 20637 12087
rect 20671 12084 20683 12087
rect 20717 12087 20775 12093
rect 20717 12084 20729 12087
rect 20671 12056 20729 12084
rect 20671 12053 20683 12056
rect 20625 12047 20683 12053
rect 20717 12053 20729 12056
rect 20763 12053 20775 12087
rect 20717 12047 20775 12053
rect 21082 12044 21088 12096
rect 21140 12084 21146 12096
rect 21361 12087 21419 12093
rect 21361 12084 21373 12087
rect 21140 12056 21373 12084
rect 21140 12044 21146 12056
rect 21361 12053 21373 12056
rect 21407 12053 21419 12087
rect 21361 12047 21419 12053
rect 22830 12044 22836 12096
rect 22888 12044 22894 12096
rect 22922 12044 22928 12096
rect 22980 12084 22986 12096
rect 23124 12084 23152 12115
rect 22980 12056 23152 12084
rect 22980 12044 22986 12056
rect 23566 12044 23572 12096
rect 23624 12084 23630 12096
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 23624 12056 23765 12084
rect 23624 12044 23630 12056
rect 23753 12053 23765 12056
rect 23799 12053 23811 12087
rect 23753 12047 23811 12053
rect 23842 12044 23848 12096
rect 23900 12044 23906 12096
rect 23934 12044 23940 12096
rect 23992 12044 23998 12096
rect 24136 12084 24164 12124
rect 24210 12112 24216 12164
rect 24268 12152 24274 12164
rect 25148 12161 25176 12192
rect 25682 12180 25688 12192
rect 25740 12222 25746 12232
rect 25777 12223 25835 12229
rect 25777 12222 25789 12223
rect 25740 12194 25789 12222
rect 25740 12180 25746 12194
rect 25777 12189 25789 12194
rect 25823 12189 25835 12223
rect 25883 12223 25941 12229
rect 25883 12222 25895 12223
rect 25777 12183 25835 12189
rect 25880 12189 25895 12222
rect 25929 12189 25941 12223
rect 25880 12183 25941 12189
rect 25133 12155 25191 12161
rect 25133 12152 25145 12155
rect 24268 12124 25145 12152
rect 24268 12112 24274 12124
rect 25133 12121 25145 12124
rect 25179 12121 25191 12155
rect 25133 12115 25191 12121
rect 25314 12112 25320 12164
rect 25372 12152 25378 12164
rect 25880 12152 25908 12183
rect 26050 12180 26056 12232
rect 26108 12180 26114 12232
rect 26160 12229 26188 12260
rect 26145 12223 26203 12229
rect 26145 12189 26157 12223
rect 26191 12189 26203 12223
rect 26252 12220 26280 12396
rect 27249 12393 27261 12427
rect 27295 12424 27307 12427
rect 27430 12424 27436 12436
rect 27295 12396 27436 12424
rect 27295 12393 27307 12396
rect 27249 12387 27307 12393
rect 27430 12384 27436 12396
rect 27488 12384 27494 12436
rect 32674 12384 32680 12436
rect 32732 12384 32738 12436
rect 26329 12291 26387 12297
rect 26329 12257 26341 12291
rect 26375 12288 26387 12291
rect 26375 12260 27568 12288
rect 26375 12257 26387 12260
rect 26329 12251 26387 12257
rect 26697 12223 26755 12229
rect 26697 12220 26709 12223
rect 26252 12192 26709 12220
rect 26145 12183 26203 12189
rect 26697 12189 26709 12192
rect 26743 12220 26755 12223
rect 26786 12220 26792 12232
rect 26743 12192 26792 12220
rect 26743 12189 26755 12192
rect 26697 12183 26755 12189
rect 26786 12180 26792 12192
rect 26844 12180 26850 12232
rect 26878 12180 26884 12232
rect 26936 12180 26942 12232
rect 27080 12229 27108 12260
rect 27540 12232 27568 12260
rect 29822 12248 29828 12300
rect 29880 12248 29886 12300
rect 32692 12288 32720 12384
rect 33045 12291 33103 12297
rect 33045 12288 33057 12291
rect 32692 12260 33057 12288
rect 33045 12257 33057 12260
rect 33091 12257 33103 12291
rect 33045 12251 33103 12257
rect 27065 12223 27123 12229
rect 27065 12189 27077 12223
rect 27111 12189 27123 12223
rect 27065 12183 27123 12189
rect 27154 12180 27160 12232
rect 27212 12220 27218 12232
rect 27341 12223 27399 12229
rect 27341 12220 27353 12223
rect 27212 12192 27353 12220
rect 27212 12180 27218 12192
rect 27341 12189 27353 12192
rect 27387 12189 27399 12223
rect 27341 12183 27399 12189
rect 27522 12180 27528 12232
rect 27580 12180 27586 12232
rect 29549 12223 29607 12229
rect 29549 12189 29561 12223
rect 29595 12189 29607 12223
rect 29549 12183 29607 12189
rect 25372 12124 25908 12152
rect 26973 12155 27031 12161
rect 25372 12112 25378 12124
rect 26973 12121 26985 12155
rect 27019 12121 27031 12155
rect 26973 12115 27031 12121
rect 29365 12155 29423 12161
rect 29365 12121 29377 12155
rect 29411 12152 29423 12155
rect 29564 12152 29592 12183
rect 30926 12180 30932 12232
rect 30984 12180 30990 12232
rect 32677 12223 32735 12229
rect 32677 12189 32689 12223
rect 32723 12220 32735 12223
rect 32766 12220 32772 12232
rect 32723 12192 32772 12220
rect 32723 12189 32735 12192
rect 32677 12183 32735 12189
rect 32766 12180 32772 12192
rect 32824 12180 32830 12232
rect 34698 12180 34704 12232
rect 34756 12180 34762 12232
rect 29730 12152 29736 12164
rect 29411 12124 29736 12152
rect 29411 12121 29423 12124
rect 29365 12115 29423 12121
rect 26694 12084 26700 12096
rect 24136 12056 26700 12084
rect 26694 12044 26700 12056
rect 26752 12044 26758 12096
rect 26988 12084 27016 12115
rect 29730 12112 29736 12124
rect 29788 12112 29794 12164
rect 34793 12155 34851 12161
rect 34793 12152 34805 12155
rect 34270 12124 34805 12152
rect 34793 12121 34805 12124
rect 34839 12121 34851 12155
rect 34793 12115 34851 12121
rect 27062 12084 27068 12096
rect 26988 12056 27068 12084
rect 27062 12044 27068 12056
rect 27120 12044 27126 12096
rect 27433 12087 27491 12093
rect 27433 12053 27445 12087
rect 27479 12084 27491 12087
rect 27706 12084 27712 12096
rect 27479 12056 27712 12084
rect 27479 12053 27491 12056
rect 27433 12047 27491 12053
rect 27706 12044 27712 12056
rect 27764 12044 27770 12096
rect 31294 12044 31300 12096
rect 31352 12044 31358 12096
rect 34514 12044 34520 12096
rect 34572 12044 34578 12096
rect 1104 11994 35236 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 35236 11994
rect 1104 11920 35236 11942
rect 4249 11883 4307 11889
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 4614 11880 4620 11892
rect 4295 11852 4620 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 7190 11840 7196 11892
rect 7248 11880 7254 11892
rect 7248 11852 7972 11880
rect 7248 11840 7254 11852
rect 7944 11821 7972 11852
rect 13078 11840 13084 11892
rect 13136 11840 13142 11892
rect 13354 11840 13360 11892
rect 13412 11840 13418 11892
rect 13906 11840 13912 11892
rect 13964 11840 13970 11892
rect 17129 11883 17187 11889
rect 17129 11849 17141 11883
rect 17175 11849 17187 11883
rect 17129 11843 17187 11849
rect 17773 11883 17831 11889
rect 17773 11849 17785 11883
rect 17819 11880 17831 11883
rect 17862 11880 17868 11892
rect 17819 11852 17868 11880
rect 17819 11849 17831 11852
rect 17773 11843 17831 11849
rect 7929 11815 7987 11821
rect 7929 11781 7941 11815
rect 7975 11781 7987 11815
rect 9585 11815 9643 11821
rect 9585 11812 9597 11815
rect 9154 11784 9597 11812
rect 7929 11775 7987 11781
rect 9585 11781 9597 11784
rect 9631 11781 9643 11815
rect 9585 11775 9643 11781
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 12342 11812 12348 11824
rect 10827 11784 12348 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 12342 11772 12348 11784
rect 12400 11772 12406 11824
rect 1394 11704 1400 11756
rect 1452 11744 1458 11756
rect 2501 11747 2559 11753
rect 2501 11744 2513 11747
rect 1452 11716 2513 11744
rect 1452 11704 1458 11716
rect 2501 11713 2513 11716
rect 2547 11713 2559 11747
rect 2501 11707 2559 11713
rect 3878 11704 3884 11756
rect 3936 11704 3942 11756
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11744 9735 11747
rect 10042 11744 10048 11756
rect 9723 11716 10048 11744
rect 9723 11713 9735 11716
rect 9677 11707 9735 11713
rect 10042 11704 10048 11716
rect 10100 11704 10106 11756
rect 10229 11747 10287 11753
rect 10229 11713 10241 11747
rect 10275 11713 10287 11747
rect 10229 11707 10287 11713
rect 2774 11636 2780 11688
rect 2832 11636 2838 11688
rect 4614 11636 4620 11688
rect 4672 11676 4678 11688
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 4672 11648 7665 11676
rect 4672 11636 4678 11648
rect 7653 11645 7665 11648
rect 7699 11676 7711 11679
rect 9401 11679 9459 11685
rect 7699 11648 8984 11676
rect 7699 11645 7711 11648
rect 7653 11639 7711 11645
rect 8956 11608 8984 11648
rect 9401 11645 9413 11679
rect 9447 11676 9459 11679
rect 10244 11676 10272 11707
rect 9447 11648 10272 11676
rect 13096 11676 13124 11840
rect 13372 11744 13400 11840
rect 16669 11815 16727 11821
rect 16669 11812 16681 11815
rect 15580 11784 16681 11812
rect 15580 11756 15608 11784
rect 13541 11747 13599 11753
rect 13541 11744 13553 11747
rect 13372 11716 13553 11744
rect 13541 11713 13553 11716
rect 13587 11713 13599 11747
rect 13541 11707 13599 11713
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 13740 11676 13768 11707
rect 15562 11704 15568 11756
rect 15620 11704 15626 11756
rect 16022 11704 16028 11756
rect 16080 11704 16086 11756
rect 16316 11753 16344 11784
rect 16669 11781 16681 11784
rect 16715 11781 16727 11815
rect 16669 11775 16727 11781
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11713 16359 11747
rect 16301 11707 16359 11713
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16485 11747 16543 11753
rect 16485 11744 16497 11747
rect 16448 11716 16497 11744
rect 16448 11704 16454 11716
rect 16485 11713 16497 11716
rect 16531 11744 16543 11747
rect 16945 11747 17003 11753
rect 16945 11744 16957 11747
rect 16531 11716 16957 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 16945 11713 16957 11716
rect 16991 11713 17003 11747
rect 17144 11744 17172 11843
rect 17862 11840 17868 11852
rect 17920 11840 17926 11892
rect 19337 11883 19395 11889
rect 19337 11849 19349 11883
rect 19383 11880 19395 11883
rect 19426 11880 19432 11892
rect 19383 11852 19432 11880
rect 19383 11849 19395 11852
rect 19337 11843 19395 11849
rect 19426 11840 19432 11852
rect 19484 11840 19490 11892
rect 20622 11840 20628 11892
rect 20680 11840 20686 11892
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21376 11852 21833 11880
rect 17313 11815 17371 11821
rect 17313 11781 17325 11815
rect 17359 11812 17371 11815
rect 20640 11812 20668 11840
rect 17359 11784 20668 11812
rect 17359 11781 17371 11784
rect 17313 11775 17371 11781
rect 20990 11772 20996 11824
rect 21048 11812 21054 11824
rect 21376 11821 21404 11852
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 22186 11840 22192 11892
rect 22244 11840 22250 11892
rect 22278 11840 22284 11892
rect 22336 11840 22342 11892
rect 23198 11840 23204 11892
rect 23256 11880 23262 11892
rect 23293 11883 23351 11889
rect 23293 11880 23305 11883
rect 23256 11852 23305 11880
rect 23256 11840 23262 11852
rect 23293 11849 23305 11852
rect 23339 11849 23351 11883
rect 23293 11843 23351 11849
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 24673 11883 24731 11889
rect 24673 11880 24685 11883
rect 23624 11852 24685 11880
rect 23624 11840 23630 11852
rect 24673 11849 24685 11852
rect 24719 11880 24731 11883
rect 24762 11880 24768 11892
rect 24719 11852 24768 11880
rect 24719 11849 24731 11852
rect 24673 11843 24731 11849
rect 24762 11840 24768 11852
rect 24820 11880 24826 11892
rect 25409 11883 25467 11889
rect 25409 11880 25421 11883
rect 24820 11852 25421 11880
rect 24820 11840 24826 11852
rect 25409 11849 25421 11852
rect 25455 11849 25467 11883
rect 25409 11843 25467 11849
rect 26421 11883 26479 11889
rect 26421 11849 26433 11883
rect 26467 11880 26479 11883
rect 26510 11880 26516 11892
rect 26467 11852 26516 11880
rect 26467 11849 26479 11852
rect 26421 11843 26479 11849
rect 26510 11840 26516 11852
rect 26568 11880 26574 11892
rect 27062 11880 27068 11892
rect 26568 11852 27068 11880
rect 26568 11840 26574 11852
rect 27062 11840 27068 11852
rect 27120 11840 27126 11892
rect 27614 11840 27620 11892
rect 27672 11840 27678 11892
rect 27706 11840 27712 11892
rect 27764 11840 27770 11892
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 28353 11883 28411 11889
rect 28353 11880 28365 11883
rect 28040 11852 28365 11880
rect 28040 11840 28046 11852
rect 28353 11849 28365 11852
rect 28399 11849 28411 11883
rect 28994 11880 29000 11892
rect 28353 11843 28411 11849
rect 28736 11852 29000 11880
rect 21177 11815 21235 11821
rect 21177 11812 21189 11815
rect 21048 11784 21189 11812
rect 21048 11772 21054 11784
rect 21177 11781 21189 11784
rect 21223 11781 21235 11815
rect 21177 11775 21235 11781
rect 21361 11815 21419 11821
rect 21361 11781 21373 11815
rect 21407 11781 21419 11815
rect 22833 11815 22891 11821
rect 22833 11812 22845 11815
rect 21361 11775 21419 11781
rect 21652 11784 22845 11812
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 17144 11716 17233 11744
rect 16945 11707 17003 11713
rect 17221 11713 17233 11716
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11713 17463 11747
rect 17405 11707 17463 11713
rect 13096 11648 13768 11676
rect 9447 11645 9459 11648
rect 9401 11639 9459 11645
rect 9582 11608 9588 11620
rect 8956 11580 9588 11608
rect 9582 11568 9588 11580
rect 9640 11568 9646 11620
rect 10042 11500 10048 11552
rect 10100 11500 10106 11552
rect 16040 11540 16068 11704
rect 16761 11679 16819 11685
rect 16761 11676 16773 11679
rect 16316 11648 16773 11676
rect 16114 11568 16120 11620
rect 16172 11617 16178 11620
rect 16172 11611 16221 11617
rect 16172 11577 16175 11611
rect 16209 11608 16221 11611
rect 16316 11608 16344 11648
rect 16761 11645 16773 11648
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 16209 11580 16344 11608
rect 16393 11611 16451 11617
rect 16209 11577 16221 11580
rect 16172 11571 16221 11577
rect 16393 11577 16405 11611
rect 16439 11608 16451 11611
rect 17420 11608 17448 11707
rect 18414 11704 18420 11756
rect 18472 11704 18478 11756
rect 18506 11704 18512 11756
rect 18564 11744 18570 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18564 11716 18613 11744
rect 18564 11704 18570 11716
rect 18601 11713 18613 11716
rect 18647 11744 18659 11747
rect 20346 11744 20352 11756
rect 18647 11716 20352 11744
rect 18647 11713 18659 11716
rect 18601 11707 18659 11713
rect 20346 11704 20352 11716
rect 20404 11744 20410 11756
rect 20717 11747 20775 11753
rect 20717 11744 20729 11747
rect 20404 11716 20729 11744
rect 20404 11704 20410 11716
rect 20717 11713 20729 11716
rect 20763 11713 20775 11747
rect 20717 11707 20775 11713
rect 21082 11704 21088 11756
rect 21140 11704 21146 11756
rect 21192 11744 21220 11775
rect 21652 11744 21680 11784
rect 22833 11781 22845 11784
rect 22879 11812 22891 11815
rect 23216 11812 23244 11840
rect 22879 11784 23244 11812
rect 22879 11781 22891 11784
rect 22833 11775 22891 11781
rect 21192 11716 21680 11744
rect 21726 11704 21732 11756
rect 21784 11744 21790 11756
rect 22649 11747 22707 11753
rect 22649 11744 22661 11747
rect 21784 11716 22661 11744
rect 21784 11704 21790 11716
rect 22649 11713 22661 11716
rect 22695 11713 22707 11747
rect 23216 11744 23244 11784
rect 23934 11772 23940 11824
rect 23992 11812 23998 11824
rect 25041 11815 25099 11821
rect 25041 11812 25053 11815
rect 23992 11784 25053 11812
rect 23992 11772 23998 11784
rect 25041 11781 25053 11784
rect 25087 11781 25099 11815
rect 25041 11775 25099 11781
rect 26694 11772 26700 11824
rect 26752 11812 26758 11824
rect 26752 11784 27384 11812
rect 26752 11772 26758 11784
rect 24029 11747 24087 11753
rect 24029 11744 24041 11747
rect 22649 11707 22707 11713
rect 22925 11737 22983 11743
rect 18782 11636 18788 11688
rect 18840 11676 18846 11688
rect 18840 11648 22416 11676
rect 18840 11636 18846 11648
rect 16439 11580 17448 11608
rect 19981 11611 20039 11617
rect 16439 11577 16451 11580
rect 16393 11571 16451 11577
rect 19981 11577 19993 11611
rect 20027 11608 20039 11611
rect 20070 11608 20076 11620
rect 20027 11580 20076 11608
rect 20027 11577 20039 11580
rect 19981 11571 20039 11577
rect 16172 11568 16178 11571
rect 20070 11568 20076 11580
rect 20128 11608 20134 11620
rect 20128 11580 21220 11608
rect 20128 11568 20134 11580
rect 21192 11552 21220 11580
rect 21358 11568 21364 11620
rect 21416 11568 21422 11620
rect 22388 11608 22416 11648
rect 22462 11636 22468 11688
rect 22520 11636 22526 11688
rect 22664 11676 22692 11707
rect 22925 11703 22937 11737
rect 22971 11703 22983 11737
rect 23216 11716 24041 11744
rect 24029 11713 24041 11716
rect 24075 11744 24087 11747
rect 24305 11747 24363 11753
rect 24305 11744 24317 11747
rect 24075 11716 24317 11744
rect 24075 11713 24087 11716
rect 24029 11707 24087 11713
rect 24305 11713 24317 11716
rect 24351 11713 24363 11747
rect 24305 11707 24363 11713
rect 25958 11704 25964 11756
rect 26016 11744 26022 11756
rect 26329 11747 26387 11753
rect 26973 11747 27031 11753
rect 26329 11744 26341 11747
rect 26016 11716 26341 11744
rect 26016 11704 26022 11716
rect 26329 11713 26341 11716
rect 26375 11744 26464 11747
rect 26973 11744 26985 11747
rect 26375 11719 26985 11744
rect 26375 11713 26387 11719
rect 26436 11716 26985 11719
rect 26329 11707 26387 11713
rect 26973 11713 26985 11716
rect 27019 11713 27031 11747
rect 26973 11707 27031 11713
rect 27062 11704 27068 11756
rect 27120 11744 27126 11756
rect 27356 11753 27384 11784
rect 27157 11747 27215 11753
rect 27157 11744 27169 11747
rect 27120 11716 27169 11744
rect 27120 11704 27126 11716
rect 27157 11713 27169 11716
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 27249 11747 27307 11753
rect 27249 11713 27261 11747
rect 27295 11713 27307 11747
rect 27249 11707 27307 11713
rect 27341 11747 27399 11753
rect 27341 11713 27353 11747
rect 27387 11713 27399 11747
rect 27632 11744 27660 11840
rect 27724 11812 27752 11840
rect 27724 11784 28028 11812
rect 28000 11753 28028 11784
rect 27709 11747 27767 11753
rect 27709 11744 27721 11747
rect 27632 11716 27721 11744
rect 27341 11707 27399 11713
rect 27709 11713 27721 11716
rect 27755 11713 27767 11747
rect 27709 11707 27767 11713
rect 27802 11747 27860 11753
rect 27802 11713 27814 11747
rect 27848 11713 27860 11747
rect 27802 11707 27860 11713
rect 27985 11747 28043 11753
rect 27985 11713 27997 11747
rect 28031 11713 28043 11747
rect 27985 11707 28043 11713
rect 22925 11697 22983 11703
rect 22830 11676 22836 11688
rect 22664 11648 22836 11676
rect 22830 11636 22836 11648
rect 22888 11636 22894 11688
rect 22940 11620 22968 11697
rect 25314 11636 25320 11688
rect 25372 11676 25378 11688
rect 26697 11679 26755 11685
rect 26697 11676 26709 11679
rect 25372 11648 26709 11676
rect 25372 11636 25378 11648
rect 26697 11645 26709 11648
rect 26743 11676 26755 11679
rect 27264 11676 27292 11707
rect 27817 11676 27845 11707
rect 28074 11704 28080 11756
rect 28132 11704 28138 11756
rect 28736 11753 28764 11852
rect 28994 11840 29000 11852
rect 29052 11880 29058 11892
rect 29730 11880 29736 11892
rect 29052 11852 29736 11880
rect 29052 11840 29058 11852
rect 29730 11840 29736 11852
rect 29788 11840 29794 11892
rect 30926 11840 30932 11892
rect 30984 11840 30990 11892
rect 31938 11840 31944 11892
rect 31996 11880 32002 11892
rect 32309 11883 32367 11889
rect 32309 11880 32321 11883
rect 31996 11852 32321 11880
rect 31996 11840 32002 11852
rect 32309 11849 32321 11852
rect 32355 11849 32367 11883
rect 32309 11843 32367 11849
rect 34514 11840 34520 11892
rect 34572 11840 34578 11892
rect 30653 11815 30711 11821
rect 30653 11812 30665 11815
rect 30222 11784 30665 11812
rect 30653 11781 30665 11784
rect 30699 11781 30711 11815
rect 30653 11775 30711 11781
rect 31294 11772 31300 11824
rect 31352 11812 31358 11824
rect 31570 11812 31576 11824
rect 31352 11784 31576 11812
rect 31352 11772 31358 11784
rect 31570 11772 31576 11784
rect 31628 11812 31634 11824
rect 31628 11784 31708 11812
rect 31628 11772 31634 11784
rect 28174 11747 28232 11753
rect 28174 11713 28186 11747
rect 28220 11713 28232 11747
rect 28174 11707 28232 11713
rect 28721 11747 28779 11753
rect 28721 11713 28733 11747
rect 28767 11713 28779 11747
rect 28721 11707 28779 11713
rect 26743 11648 27292 11676
rect 27724 11648 27845 11676
rect 26743 11645 26755 11648
rect 26697 11639 26755 11645
rect 22922 11608 22928 11620
rect 22388 11580 22928 11608
rect 22922 11568 22928 11580
rect 22980 11568 22986 11620
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 16040 11512 16681 11540
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 16669 11503 16727 11509
rect 18322 11500 18328 11552
rect 18380 11540 18386 11552
rect 19334 11540 19340 11552
rect 18380 11512 19340 11540
rect 18380 11500 18386 11512
rect 19334 11500 19340 11512
rect 19392 11540 19398 11552
rect 19613 11543 19671 11549
rect 19613 11540 19625 11543
rect 19392 11512 19625 11540
rect 19392 11500 19398 11512
rect 19613 11509 19625 11512
rect 19659 11509 19671 11543
rect 19613 11503 19671 11509
rect 20346 11500 20352 11552
rect 20404 11500 20410 11552
rect 21174 11500 21180 11552
rect 21232 11500 21238 11552
rect 22278 11500 22284 11552
rect 22336 11540 22342 11552
rect 22649 11543 22707 11549
rect 22649 11540 22661 11543
rect 22336 11512 22661 11540
rect 22336 11500 22342 11512
rect 22649 11509 22661 11512
rect 22695 11540 22707 11543
rect 22738 11540 22744 11552
rect 22695 11512 22744 11540
rect 22695 11509 22707 11512
rect 22649 11503 22707 11509
rect 22738 11500 22744 11512
rect 22796 11500 22802 11552
rect 23290 11500 23296 11552
rect 23348 11540 23354 11552
rect 23569 11543 23627 11549
rect 23569 11540 23581 11543
rect 23348 11512 23581 11540
rect 23348 11500 23354 11512
rect 23569 11509 23581 11512
rect 23615 11509 23627 11543
rect 23569 11503 23627 11509
rect 25682 11500 25688 11552
rect 25740 11540 25746 11552
rect 26605 11543 26663 11549
rect 26605 11540 26617 11543
rect 25740 11512 26617 11540
rect 25740 11500 25746 11512
rect 26605 11509 26617 11512
rect 26651 11540 26663 11543
rect 26694 11540 26700 11552
rect 26651 11512 26700 11540
rect 26651 11509 26663 11512
rect 26605 11503 26663 11509
rect 26694 11500 26700 11512
rect 26752 11500 26758 11552
rect 26789 11543 26847 11549
rect 26789 11509 26801 11543
rect 26835 11540 26847 11543
rect 27246 11540 27252 11552
rect 26835 11512 27252 11540
rect 26835 11509 26847 11512
rect 26789 11503 26847 11509
rect 27246 11500 27252 11512
rect 27304 11540 27310 11552
rect 27724 11540 27752 11648
rect 27890 11636 27896 11688
rect 27948 11676 27954 11688
rect 28184 11676 28212 11707
rect 30374 11704 30380 11756
rect 30432 11744 30438 11756
rect 31680 11753 31708 11784
rect 30745 11747 30803 11753
rect 30745 11744 30757 11747
rect 30432 11716 30757 11744
rect 30432 11704 30438 11716
rect 30745 11713 30757 11716
rect 30791 11744 30803 11747
rect 31021 11747 31079 11753
rect 31021 11744 31033 11747
rect 30791 11716 31033 11744
rect 30791 11713 30803 11716
rect 30745 11707 30803 11713
rect 31021 11713 31033 11716
rect 31067 11744 31079 11747
rect 31389 11747 31447 11753
rect 31389 11744 31401 11747
rect 31067 11716 31401 11744
rect 31067 11713 31079 11716
rect 31021 11707 31079 11713
rect 31389 11713 31401 11716
rect 31435 11713 31447 11747
rect 31389 11707 31447 11713
rect 31665 11747 31723 11753
rect 31665 11713 31677 11747
rect 31711 11713 31723 11747
rect 31665 11707 31723 11713
rect 28997 11679 29055 11685
rect 28997 11676 29009 11679
rect 27948 11648 28212 11676
rect 28276 11648 29009 11676
rect 27948 11636 27954 11648
rect 27798 11568 27804 11620
rect 27856 11608 27862 11620
rect 28276 11608 28304 11648
rect 28997 11645 29009 11648
rect 29043 11645 29055 11679
rect 28997 11639 29055 11645
rect 31478 11636 31484 11688
rect 31536 11676 31542 11688
rect 31956 11685 31984 11840
rect 34532 11744 34560 11840
rect 34701 11747 34759 11753
rect 34701 11744 34713 11747
rect 34532 11716 34713 11744
rect 34701 11713 34713 11716
rect 34747 11713 34759 11747
rect 34701 11707 34759 11713
rect 34790 11704 34796 11756
rect 34848 11704 34854 11756
rect 31757 11679 31815 11685
rect 31757 11676 31769 11679
rect 31536 11648 31769 11676
rect 31536 11636 31542 11648
rect 31757 11645 31769 11648
rect 31803 11645 31815 11679
rect 31757 11639 31815 11645
rect 31941 11679 31999 11685
rect 31941 11645 31953 11679
rect 31987 11645 31999 11679
rect 31941 11639 31999 11645
rect 34425 11679 34483 11685
rect 34425 11645 34437 11679
rect 34471 11676 34483 11679
rect 34808 11676 34836 11704
rect 34471 11648 34836 11676
rect 34471 11645 34483 11648
rect 34425 11639 34483 11645
rect 27856 11580 28304 11608
rect 27856 11568 27862 11580
rect 27304 11512 27752 11540
rect 27304 11500 27310 11512
rect 30466 11500 30472 11552
rect 30524 11500 30530 11552
rect 31846 11500 31852 11552
rect 31904 11500 31910 11552
rect 1104 11450 35248 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 35248 11450
rect 1104 11376 35248 11398
rect 1578 11296 1584 11348
rect 1636 11296 1642 11348
rect 17954 11296 17960 11348
rect 18012 11336 18018 11348
rect 18141 11339 18199 11345
rect 18141 11336 18153 11339
rect 18012 11308 18153 11336
rect 18012 11296 18018 11308
rect 18141 11305 18153 11308
rect 18187 11305 18199 11339
rect 18141 11299 18199 11305
rect 18414 11296 18420 11348
rect 18472 11296 18478 11348
rect 18506 11296 18512 11348
rect 18564 11296 18570 11348
rect 20165 11339 20223 11345
rect 20165 11305 20177 11339
rect 20211 11336 20223 11339
rect 20990 11336 20996 11348
rect 20211 11308 20996 11336
rect 20211 11305 20223 11308
rect 20165 11299 20223 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 22186 11296 22192 11348
rect 22244 11336 22250 11348
rect 22281 11339 22339 11345
rect 22281 11336 22293 11339
rect 22244 11308 22293 11336
rect 22244 11296 22250 11308
rect 22281 11305 22293 11308
rect 22327 11305 22339 11339
rect 22281 11299 22339 11305
rect 22554 11296 22560 11348
rect 22612 11336 22618 11348
rect 22649 11339 22707 11345
rect 22649 11336 22661 11339
rect 22612 11308 22661 11336
rect 22612 11296 22618 11308
rect 22649 11305 22661 11308
rect 22695 11336 22707 11339
rect 23934 11336 23940 11348
rect 22695 11308 23940 11336
rect 22695 11305 22707 11308
rect 22649 11299 22707 11305
rect 23934 11296 23940 11308
rect 23992 11296 23998 11348
rect 24210 11296 24216 11348
rect 24268 11296 24274 11348
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 27706 11296 27712 11348
rect 27764 11296 27770 11348
rect 27801 11339 27859 11345
rect 27801 11305 27813 11339
rect 27847 11336 27859 11339
rect 28350 11336 28356 11348
rect 27847 11308 28356 11336
rect 27847 11305 27859 11308
rect 27801 11299 27859 11305
rect 28350 11296 28356 11308
rect 28408 11296 28414 11348
rect 28629 11339 28687 11345
rect 28629 11305 28641 11339
rect 28675 11336 28687 11339
rect 28994 11336 29000 11348
rect 28675 11308 29000 11336
rect 28675 11305 28687 11308
rect 28629 11299 28687 11305
rect 28994 11296 29000 11308
rect 29052 11296 29058 11348
rect 30466 11296 30472 11348
rect 30524 11296 30530 11348
rect 31478 11296 31484 11348
rect 31536 11296 31542 11348
rect 31754 11296 31760 11348
rect 31812 11296 31818 11348
rect 31846 11296 31852 11348
rect 31904 11296 31910 11348
rect 18432 11268 18460 11296
rect 18877 11271 18935 11277
rect 18877 11268 18889 11271
rect 18432 11240 18889 11268
rect 18877 11237 18889 11240
rect 18923 11237 18935 11271
rect 18877 11231 18935 11237
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 21008 11132 21036 11296
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 21361 11271 21419 11277
rect 21361 11268 21373 11271
rect 21232 11240 21373 11268
rect 21232 11228 21238 11240
rect 21361 11237 21373 11240
rect 21407 11268 21419 11271
rect 21729 11271 21787 11277
rect 21729 11268 21741 11271
rect 21407 11240 21741 11268
rect 21407 11237 21419 11240
rect 21361 11231 21419 11237
rect 21729 11237 21741 11240
rect 21775 11268 21787 11271
rect 22094 11268 22100 11280
rect 21775 11240 22100 11268
rect 21775 11237 21787 11240
rect 21729 11231 21787 11237
rect 22094 11228 22100 11240
rect 22152 11268 22158 11280
rect 22572 11268 22600 11296
rect 22152 11240 22600 11268
rect 22152 11228 22158 11240
rect 22830 11228 22836 11280
rect 22888 11268 22894 11280
rect 24670 11268 24676 11280
rect 22888 11240 24676 11268
rect 22888 11228 22894 11240
rect 22002 11132 22008 11144
rect 21008 11104 22008 11132
rect 22002 11092 22008 11104
rect 22060 11132 22066 11144
rect 22097 11135 22155 11141
rect 22097 11132 22109 11135
rect 22060 11104 22109 11132
rect 22060 11092 22066 11104
rect 22097 11101 22109 11104
rect 22143 11101 22155 11135
rect 22097 11095 22155 11101
rect 22278 11092 22284 11144
rect 22336 11092 22342 11144
rect 22370 11092 22376 11144
rect 22428 11132 22434 11144
rect 22830 11132 22836 11144
rect 22428 11104 22836 11132
rect 22428 11092 22434 11104
rect 22830 11092 22836 11104
rect 22888 11132 22894 11144
rect 23017 11135 23075 11141
rect 23017 11132 23029 11135
rect 22888 11104 23029 11132
rect 22888 11092 22894 11104
rect 23017 11101 23029 11104
rect 23063 11101 23075 11135
rect 23017 11095 23075 11101
rect 23201 11135 23259 11141
rect 23201 11101 23213 11135
rect 23247 11101 23259 11135
rect 23308 11132 23336 11240
rect 24670 11228 24676 11240
rect 24728 11228 24734 11280
rect 25332 11268 25360 11296
rect 25869 11271 25927 11277
rect 25869 11268 25881 11271
rect 25332 11240 25881 11268
rect 25869 11237 25881 11240
rect 25915 11237 25927 11271
rect 25869 11231 25927 11237
rect 23385 11203 23443 11209
rect 23385 11169 23397 11203
rect 23431 11200 23443 11203
rect 23569 11203 23627 11209
rect 23569 11200 23581 11203
rect 23431 11172 23581 11200
rect 23431 11169 23443 11172
rect 23385 11163 23443 11169
rect 23569 11169 23581 11172
rect 23615 11200 23627 11203
rect 25884 11200 25912 11231
rect 27724 11200 27752 11296
rect 27890 11228 27896 11280
rect 27948 11228 27954 11280
rect 28074 11228 28080 11280
rect 28132 11228 28138 11280
rect 23615 11172 24532 11200
rect 23615 11169 23627 11172
rect 23569 11163 23627 11169
rect 24504 11144 24532 11172
rect 24596 11172 25176 11200
rect 25884 11172 27108 11200
rect 23477 11135 23535 11141
rect 23477 11132 23489 11135
rect 23308 11104 23489 11132
rect 23201 11095 23259 11101
rect 23477 11101 23489 11104
rect 23523 11101 23535 11135
rect 23477 11095 23535 11101
rect 9582 11024 9588 11076
rect 9640 11024 9646 11076
rect 19334 11024 19340 11076
rect 19392 11064 19398 11076
rect 20438 11064 20444 11076
rect 19392 11036 20444 11064
rect 19392 11024 19398 11036
rect 20438 11024 20444 11036
rect 20496 11064 20502 11076
rect 22646 11064 22652 11076
rect 20496 11036 22652 11064
rect 20496 11024 20502 11036
rect 22646 11024 22652 11036
rect 22704 11064 22710 11076
rect 23216 11064 23244 11095
rect 23658 11092 23664 11144
rect 23716 11132 23722 11144
rect 23937 11135 23995 11141
rect 23937 11132 23949 11135
rect 23716 11104 23949 11132
rect 23716 11092 23722 11104
rect 23937 11101 23949 11104
rect 23983 11101 23995 11135
rect 23937 11095 23995 11101
rect 24026 11092 24032 11144
rect 24084 11092 24090 11144
rect 24394 11092 24400 11144
rect 24452 11092 24458 11144
rect 24486 11092 24492 11144
rect 24544 11092 24550 11144
rect 22704 11036 23244 11064
rect 22704 11024 22710 11036
rect 23566 11024 23572 11076
rect 23624 11064 23630 11076
rect 23753 11067 23811 11073
rect 23753 11064 23765 11067
rect 23624 11036 23765 11064
rect 23624 11024 23630 11036
rect 23753 11033 23765 11036
rect 23799 11033 23811 11067
rect 23753 11027 23811 11033
rect 23845 11067 23903 11073
rect 23845 11033 23857 11067
rect 23891 11064 23903 11067
rect 24044 11064 24072 11092
rect 24596 11064 24624 11172
rect 24762 11092 24768 11144
rect 24820 11092 24826 11144
rect 25148 11141 25176 11172
rect 25133 11135 25191 11141
rect 25133 11101 25145 11135
rect 25179 11101 25191 11135
rect 25133 11095 25191 11101
rect 25498 11092 25504 11144
rect 25556 11092 25562 11144
rect 25961 11135 26019 11141
rect 25961 11101 25973 11135
rect 26007 11101 26019 11135
rect 25961 11095 26019 11101
rect 23891 11036 24624 11064
rect 23891 11033 23903 11036
rect 23845 11027 23903 11033
rect 24670 11024 24676 11076
rect 24728 11064 24734 11076
rect 25976 11064 26004 11095
rect 26694 11092 26700 11144
rect 26752 11132 26758 11144
rect 27080 11141 27108 11172
rect 27448 11172 27752 11200
rect 26881 11135 26939 11141
rect 26881 11132 26893 11135
rect 26752 11104 26893 11132
rect 26752 11092 26758 11104
rect 26881 11101 26893 11104
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 27065 11135 27123 11141
rect 27065 11101 27077 11135
rect 27111 11101 27123 11135
rect 27065 11095 27123 11101
rect 27246 11092 27252 11144
rect 27304 11092 27310 11144
rect 27448 11141 27476 11172
rect 27433 11135 27491 11141
rect 27433 11101 27445 11135
rect 27479 11101 27491 11135
rect 27433 11095 27491 11101
rect 27614 11092 27620 11144
rect 27672 11132 27678 11144
rect 27908 11132 27936 11228
rect 27672 11104 27936 11132
rect 27672 11092 27678 11104
rect 24728 11036 26004 11064
rect 26973 11067 27031 11073
rect 24728 11024 24734 11036
rect 26973 11033 26985 11067
rect 27019 11064 27031 11067
rect 27525 11067 27583 11073
rect 27525 11064 27537 11067
rect 27019 11036 27537 11064
rect 27019 11033 27031 11036
rect 26973 11027 27031 11033
rect 27525 11033 27537 11036
rect 27571 11064 27583 11067
rect 28092 11064 28120 11228
rect 30484 11200 30512 11296
rect 31389 11203 31447 11209
rect 31389 11200 31401 11203
rect 30484 11172 31401 11200
rect 31389 11169 31401 11172
rect 31435 11200 31447 11203
rect 31864 11200 31892 11296
rect 32401 11271 32459 11277
rect 32401 11237 32413 11271
rect 32447 11237 32459 11271
rect 32401 11231 32459 11237
rect 31941 11203 31999 11209
rect 31941 11200 31953 11203
rect 31435 11172 31754 11200
rect 31864 11172 31953 11200
rect 31435 11169 31447 11172
rect 31389 11163 31447 11169
rect 31726 11144 31754 11172
rect 31941 11169 31953 11172
rect 31987 11169 31999 11203
rect 32416 11200 32444 11231
rect 33045 11203 33103 11209
rect 33045 11200 33057 11203
rect 32416 11172 33057 11200
rect 31941 11163 31999 11169
rect 33045 11169 33057 11172
rect 33091 11169 33103 11203
rect 33045 11163 33103 11169
rect 34517 11203 34575 11209
rect 34517 11169 34529 11203
rect 34563 11200 34575 11203
rect 34606 11200 34612 11212
rect 34563 11172 34612 11200
rect 34563 11169 34575 11172
rect 34517 11163 34575 11169
rect 34606 11160 34612 11172
rect 34664 11160 34670 11212
rect 31570 11092 31576 11144
rect 31628 11092 31634 11144
rect 31726 11104 31760 11144
rect 31754 11092 31760 11104
rect 31812 11132 31818 11144
rect 32033 11135 32091 11141
rect 32033 11132 32045 11135
rect 31812 11104 32045 11132
rect 31812 11092 31818 11104
rect 32033 11101 32045 11104
rect 32079 11101 32091 11135
rect 32033 11095 32091 11101
rect 32766 11092 32772 11144
rect 32824 11092 32830 11144
rect 34698 11092 34704 11144
rect 34756 11092 34762 11144
rect 27571 11036 28120 11064
rect 27571 11033 27583 11036
rect 27525 11027 27583 11033
rect 30374 11024 30380 11076
rect 30432 11024 30438 11076
rect 31110 11024 31116 11076
rect 31168 11064 31174 11076
rect 31297 11067 31355 11073
rect 31297 11064 31309 11067
rect 31168 11036 31309 11064
rect 31168 11024 31174 11036
rect 31297 11033 31309 11036
rect 31343 11033 31355 11067
rect 34793 11067 34851 11073
rect 34793 11064 34805 11067
rect 34270 11036 34805 11064
rect 31297 11027 31355 11033
rect 34793 11033 34805 11036
rect 34839 11033 34851 11067
rect 34793 11027 34851 11033
rect 19426 10956 19432 11008
rect 19484 10996 19490 11008
rect 28902 10996 28908 11008
rect 19484 10968 28908 10996
rect 19484 10956 19490 10968
rect 28902 10956 28908 10968
rect 28960 10996 28966 11008
rect 30392 10996 30420 11024
rect 28960 10968 30420 10996
rect 28960 10956 28966 10968
rect 1104 10906 35236 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 35236 10906
rect 1104 10832 35236 10854
rect 10594 10752 10600 10804
rect 10652 10792 10658 10804
rect 19334 10792 19340 10804
rect 10652 10764 19340 10792
rect 10652 10752 10658 10764
rect 19334 10752 19340 10764
rect 19392 10752 19398 10804
rect 20990 10752 20996 10804
rect 21048 10752 21054 10804
rect 22094 10752 22100 10804
rect 22152 10752 22158 10804
rect 23569 10795 23627 10801
rect 22480 10764 23244 10792
rect 19984 10736 20036 10742
rect 21008 10724 21036 10752
rect 19984 10678 20036 10684
rect 20640 10696 21036 10724
rect 22112 10724 22140 10752
rect 22112 10696 22324 10724
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 9309 10659 9367 10665
rect 9309 10656 9321 10659
rect 3292 10628 9321 10656
rect 3292 10616 3298 10628
rect 9309 10625 9321 10628
rect 9355 10656 9367 10659
rect 9355 10628 11836 10656
rect 9355 10625 9367 10628
rect 9309 10619 9367 10625
rect 11808 10529 11836 10628
rect 18690 10616 18696 10668
rect 18748 10616 18754 10668
rect 19242 10616 19248 10668
rect 19300 10616 19306 10668
rect 20438 10616 20444 10668
rect 20496 10616 20502 10668
rect 20640 10665 20668 10696
rect 20625 10659 20683 10665
rect 20625 10625 20637 10659
rect 20671 10625 20683 10659
rect 20625 10619 20683 10625
rect 20717 10659 20775 10665
rect 20717 10625 20729 10659
rect 20763 10625 20775 10659
rect 20717 10619 20775 10625
rect 20901 10659 20959 10665
rect 20901 10625 20913 10659
rect 20947 10656 20959 10659
rect 20947 10628 21312 10656
rect 20947 10625 20959 10628
rect 20901 10619 20959 10625
rect 19978 10548 19984 10600
rect 20036 10588 20042 10600
rect 20732 10588 20760 10619
rect 21284 10600 21312 10628
rect 21358 10616 21364 10668
rect 21416 10656 21422 10668
rect 22296 10665 22324 10696
rect 22097 10659 22155 10665
rect 22097 10656 22109 10659
rect 21416 10628 22109 10656
rect 21416 10616 21422 10628
rect 22097 10625 22109 10628
rect 22143 10625 22155 10659
rect 22097 10619 22155 10625
rect 22281 10659 22339 10665
rect 22281 10625 22293 10659
rect 22327 10625 22339 10659
rect 22480 10656 22508 10764
rect 22646 10684 22652 10736
rect 22704 10724 22710 10736
rect 22704 10696 23060 10724
rect 22704 10684 22710 10696
rect 23032 10668 23060 10696
rect 22281 10619 22339 10625
rect 22388 10628 22508 10656
rect 21174 10588 21180 10600
rect 20036 10560 21180 10588
rect 20036 10548 20042 10560
rect 21174 10548 21180 10560
rect 21232 10548 21238 10600
rect 21266 10548 21272 10600
rect 21324 10588 21330 10600
rect 22388 10588 22416 10628
rect 22554 10616 22560 10668
rect 22612 10616 22618 10668
rect 23014 10616 23020 10668
rect 23072 10616 23078 10668
rect 23216 10665 23244 10764
rect 23569 10761 23581 10795
rect 23615 10792 23627 10795
rect 23842 10792 23848 10804
rect 23615 10764 23848 10792
rect 23615 10761 23627 10764
rect 23569 10755 23627 10761
rect 23842 10752 23848 10764
rect 23900 10752 23906 10804
rect 25498 10752 25504 10804
rect 25556 10752 25562 10804
rect 25774 10752 25780 10804
rect 25832 10752 25838 10804
rect 27433 10795 27491 10801
rect 27433 10761 27445 10795
rect 27479 10792 27491 10795
rect 27522 10792 27528 10804
rect 27479 10764 27528 10792
rect 27479 10761 27491 10764
rect 27433 10755 27491 10761
rect 27522 10752 27528 10764
rect 27580 10752 27586 10804
rect 28994 10752 29000 10804
rect 29052 10792 29058 10804
rect 29362 10792 29368 10804
rect 29052 10764 29368 10792
rect 29052 10752 29058 10764
rect 29362 10752 29368 10764
rect 29420 10752 29426 10804
rect 31297 10795 31355 10801
rect 31297 10761 31309 10795
rect 31343 10792 31355 10795
rect 31938 10792 31944 10804
rect 31343 10764 31944 10792
rect 31343 10761 31355 10764
rect 31297 10755 31355 10761
rect 24394 10684 24400 10736
rect 24452 10684 24458 10736
rect 24486 10684 24492 10736
rect 24544 10724 24550 10736
rect 25516 10724 25544 10752
rect 24544 10696 25544 10724
rect 25792 10724 25820 10752
rect 25869 10727 25927 10733
rect 25869 10724 25881 10727
rect 25792 10696 25881 10724
rect 24544 10684 24550 10696
rect 23201 10659 23259 10665
rect 23201 10625 23213 10659
rect 23247 10625 23259 10659
rect 23201 10619 23259 10625
rect 21324 10560 22416 10588
rect 21324 10548 21330 10560
rect 22462 10548 22468 10600
rect 22520 10588 22526 10600
rect 22649 10591 22707 10597
rect 22649 10588 22661 10591
rect 22520 10560 22661 10588
rect 22520 10548 22526 10560
rect 22649 10557 22661 10560
rect 22695 10588 22707 10591
rect 23109 10591 23167 10597
rect 23109 10588 23121 10591
rect 22695 10560 23121 10588
rect 22695 10557 22707 10560
rect 22649 10551 22707 10557
rect 23109 10557 23121 10560
rect 23155 10557 23167 10591
rect 23216 10588 23244 10619
rect 23566 10616 23572 10668
rect 23624 10656 23630 10668
rect 24412 10656 24440 10684
rect 23624 10628 24440 10656
rect 23624 10616 23630 10628
rect 24670 10616 24676 10668
rect 24728 10616 24734 10668
rect 24872 10665 24900 10696
rect 25869 10693 25881 10696
rect 25915 10724 25927 10727
rect 26510 10724 26516 10736
rect 25915 10696 26516 10724
rect 25915 10693 25927 10696
rect 25869 10687 25927 10693
rect 26510 10684 26516 10696
rect 26568 10724 26574 10736
rect 26568 10696 27200 10724
rect 26568 10684 26574 10696
rect 24857 10659 24915 10665
rect 24857 10625 24869 10659
rect 24903 10625 24915 10659
rect 24857 10619 24915 10625
rect 24949 10659 25007 10665
rect 24949 10625 24961 10659
rect 24995 10625 25007 10659
rect 24949 10619 25007 10625
rect 23658 10588 23664 10600
rect 23216 10560 23664 10588
rect 23109 10551 23167 10557
rect 23658 10548 23664 10560
rect 23716 10588 23722 10600
rect 23845 10591 23903 10597
rect 23845 10588 23857 10591
rect 23716 10560 23857 10588
rect 23716 10548 23722 10560
rect 23845 10557 23857 10560
rect 23891 10588 23903 10591
rect 24210 10588 24216 10600
rect 23891 10560 24216 10588
rect 23891 10557 23903 10560
rect 23845 10551 23903 10557
rect 24210 10548 24216 10560
rect 24268 10548 24274 10600
rect 11793 10523 11851 10529
rect 11793 10489 11805 10523
rect 11839 10520 11851 10523
rect 21545 10523 21603 10529
rect 11839 10492 12434 10520
rect 11839 10489 11851 10492
rect 11793 10483 11851 10489
rect 12406 10452 12434 10492
rect 21545 10489 21557 10523
rect 21591 10520 21603 10523
rect 22738 10520 22744 10532
rect 21591 10492 22744 10520
rect 21591 10489 21603 10492
rect 21545 10483 21603 10489
rect 22738 10480 22744 10492
rect 22796 10480 22802 10532
rect 22925 10523 22983 10529
rect 22925 10489 22937 10523
rect 22971 10520 22983 10523
rect 24964 10520 24992 10619
rect 25038 10616 25044 10668
rect 25096 10656 25102 10668
rect 25593 10659 25651 10665
rect 25593 10656 25605 10659
rect 25096 10628 25605 10656
rect 25096 10616 25102 10628
rect 25593 10625 25605 10628
rect 25639 10625 25651 10659
rect 25593 10619 25651 10625
rect 25777 10659 25835 10665
rect 25777 10625 25789 10659
rect 25823 10625 25835 10659
rect 25777 10619 25835 10625
rect 25222 10548 25228 10600
rect 25280 10588 25286 10600
rect 25792 10588 25820 10619
rect 25958 10616 25964 10668
rect 26016 10616 26022 10668
rect 27172 10665 27200 10696
rect 26237 10659 26295 10665
rect 26068 10654 26188 10656
rect 26237 10654 26249 10659
rect 26068 10628 26249 10654
rect 25280 10560 25820 10588
rect 25280 10548 25286 10560
rect 25501 10523 25559 10529
rect 22971 10492 25452 10520
rect 22971 10489 22983 10492
rect 22925 10483 22983 10489
rect 17218 10452 17224 10464
rect 12406 10424 17224 10452
rect 17218 10412 17224 10424
rect 17276 10412 17282 10464
rect 20530 10412 20536 10464
rect 20588 10412 20594 10464
rect 20806 10412 20812 10464
rect 20864 10412 20870 10464
rect 22189 10455 22247 10461
rect 22189 10421 22201 10455
rect 22235 10452 22247 10455
rect 22278 10452 22284 10464
rect 22235 10424 22284 10452
rect 22235 10421 22247 10424
rect 22189 10415 22247 10421
rect 22278 10412 22284 10424
rect 22336 10452 22342 10464
rect 22557 10455 22615 10461
rect 22557 10452 22569 10455
rect 22336 10424 22569 10452
rect 22336 10412 22342 10424
rect 22557 10421 22569 10424
rect 22603 10421 22615 10455
rect 22557 10415 22615 10421
rect 24857 10455 24915 10461
rect 24857 10421 24869 10455
rect 24903 10452 24915 10455
rect 25038 10452 25044 10464
rect 24903 10424 25044 10452
rect 24903 10421 24915 10424
rect 24857 10415 24915 10421
rect 25038 10412 25044 10424
rect 25096 10412 25102 10464
rect 25424 10452 25452 10492
rect 25501 10489 25513 10523
rect 25547 10520 25559 10523
rect 26068 10520 26096 10628
rect 26160 10626 26249 10628
rect 26237 10625 26249 10626
rect 26283 10625 26295 10659
rect 26237 10619 26295 10625
rect 26421 10659 26479 10665
rect 26421 10625 26433 10659
rect 26467 10625 26479 10659
rect 26421 10619 26479 10625
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 26436 10588 26464 10619
rect 28902 10616 28908 10668
rect 28960 10656 28966 10668
rect 29825 10659 29883 10665
rect 29825 10656 29837 10659
rect 28960 10628 29837 10656
rect 28960 10616 28966 10628
rect 29825 10625 29837 10628
rect 29871 10656 29883 10659
rect 30009 10659 30067 10665
rect 30009 10656 30021 10659
rect 29871 10628 30021 10656
rect 29871 10625 29883 10628
rect 29825 10619 29883 10625
rect 30009 10625 30021 10628
rect 30055 10625 30067 10659
rect 30009 10619 30067 10625
rect 31478 10616 31484 10668
rect 31536 10616 31542 10668
rect 31570 10616 31576 10668
rect 31628 10616 31634 10668
rect 31754 10616 31760 10668
rect 31812 10616 31818 10668
rect 31864 10665 31892 10764
rect 31938 10752 31944 10764
rect 31996 10752 32002 10804
rect 32677 10795 32735 10801
rect 32677 10761 32689 10795
rect 32723 10792 32735 10795
rect 32766 10792 32772 10804
rect 32723 10764 32772 10792
rect 32723 10761 32735 10764
rect 32677 10755 32735 10761
rect 32766 10752 32772 10764
rect 32824 10792 32830 10804
rect 32953 10795 33011 10801
rect 32953 10792 32965 10795
rect 32824 10764 32965 10792
rect 32824 10752 32830 10764
rect 32953 10761 32965 10764
rect 32999 10761 33011 10795
rect 32953 10755 33011 10761
rect 31849 10659 31907 10665
rect 31849 10625 31861 10659
rect 31895 10625 31907 10659
rect 31849 10619 31907 10625
rect 32214 10616 32220 10668
rect 32272 10616 32278 10668
rect 26160 10560 26464 10588
rect 27065 10591 27123 10597
rect 26160 10529 26188 10560
rect 27065 10557 27077 10591
rect 27111 10557 27123 10591
rect 27065 10551 27123 10557
rect 25547 10492 26096 10520
rect 26145 10523 26203 10529
rect 25547 10489 25559 10492
rect 25501 10483 25559 10489
rect 26145 10489 26157 10523
rect 26191 10489 26203 10523
rect 26145 10483 26203 10489
rect 26326 10480 26332 10532
rect 26384 10480 26390 10532
rect 27080 10452 27108 10551
rect 27246 10548 27252 10600
rect 27304 10548 27310 10600
rect 31294 10480 31300 10532
rect 31352 10520 31358 10532
rect 31496 10520 31524 10616
rect 31588 10588 31616 10616
rect 32232 10588 32260 10616
rect 31588 10560 32260 10588
rect 31665 10523 31723 10529
rect 31665 10520 31677 10523
rect 31352 10492 31677 10520
rect 31352 10480 31358 10492
rect 31665 10489 31677 10492
rect 31711 10489 31723 10523
rect 31665 10483 31723 10489
rect 27522 10452 27528 10464
rect 25424 10424 27528 10452
rect 27522 10412 27528 10424
rect 27580 10412 27586 10464
rect 30098 10412 30104 10464
rect 30156 10412 30162 10464
rect 31386 10412 31392 10464
rect 31444 10412 31450 10464
rect 34054 10412 34060 10464
rect 34112 10452 34118 10464
rect 34149 10455 34207 10461
rect 34149 10452 34161 10455
rect 34112 10424 34161 10452
rect 34112 10412 34118 10424
rect 34149 10421 34161 10424
rect 34195 10452 34207 10455
rect 34517 10455 34575 10461
rect 34517 10452 34529 10455
rect 34195 10424 34529 10452
rect 34195 10421 34207 10424
rect 34149 10415 34207 10421
rect 34517 10421 34529 10424
rect 34563 10452 34575 10455
rect 34698 10452 34704 10464
rect 34563 10424 34704 10452
rect 34563 10421 34575 10424
rect 34517 10415 34575 10421
rect 34698 10412 34704 10424
rect 34756 10412 34762 10464
rect 1104 10362 35248 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 35248 10362
rect 1104 10288 35248 10310
rect 4065 10251 4123 10257
rect 4065 10217 4077 10251
rect 4111 10248 4123 10251
rect 4614 10248 4620 10260
rect 4111 10220 4620 10248
rect 4111 10217 4123 10220
rect 4065 10211 4123 10217
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10112 1639 10115
rect 4080 10112 4108 10211
rect 4614 10208 4620 10220
rect 4672 10208 4678 10260
rect 18690 10208 18696 10260
rect 18748 10208 18754 10260
rect 19242 10208 19248 10260
rect 19300 10248 19306 10260
rect 19521 10251 19579 10257
rect 19521 10248 19533 10251
rect 19300 10220 19533 10248
rect 19300 10208 19306 10220
rect 19521 10217 19533 10220
rect 19567 10217 19579 10251
rect 19521 10211 19579 10217
rect 19978 10208 19984 10260
rect 20036 10208 20042 10260
rect 20530 10208 20536 10260
rect 20588 10208 20594 10260
rect 20806 10208 20812 10260
rect 20864 10208 20870 10260
rect 21266 10208 21272 10260
rect 21324 10208 21330 10260
rect 22002 10208 22008 10260
rect 22060 10208 22066 10260
rect 22830 10208 22836 10260
rect 22888 10208 22894 10260
rect 23014 10208 23020 10260
rect 23072 10248 23078 10260
rect 23201 10251 23259 10257
rect 23201 10248 23213 10251
rect 23072 10220 23213 10248
rect 23072 10208 23078 10220
rect 23201 10217 23213 10220
rect 23247 10217 23259 10251
rect 23201 10211 23259 10217
rect 23661 10251 23719 10257
rect 23661 10217 23673 10251
rect 23707 10248 23719 10251
rect 24026 10248 24032 10260
rect 23707 10220 24032 10248
rect 23707 10217 23719 10220
rect 23661 10211 23719 10217
rect 24026 10208 24032 10220
rect 24084 10208 24090 10260
rect 24210 10208 24216 10260
rect 24268 10248 24274 10260
rect 24581 10251 24639 10257
rect 24581 10248 24593 10251
rect 24268 10220 24593 10248
rect 24268 10208 24274 10220
rect 24581 10217 24593 10220
rect 24627 10217 24639 10251
rect 24581 10211 24639 10217
rect 24765 10251 24823 10257
rect 24765 10217 24777 10251
rect 24811 10248 24823 10251
rect 25222 10248 25228 10260
rect 24811 10220 25228 10248
rect 24811 10217 24823 10220
rect 24765 10211 24823 10217
rect 25222 10208 25228 10220
rect 25280 10208 25286 10260
rect 26142 10208 26148 10260
rect 26200 10248 26206 10260
rect 26200 10220 28212 10248
rect 26200 10208 26206 10220
rect 1627 10084 4108 10112
rect 18141 10115 18199 10121
rect 1627 10081 1639 10084
rect 1581 10075 1639 10081
rect 18141 10081 18153 10115
rect 18187 10112 18199 10115
rect 18322 10112 18328 10124
rect 18187 10084 18328 10112
rect 18187 10081 18199 10084
rect 18141 10075 18199 10081
rect 18322 10072 18328 10084
rect 18380 10112 18386 10124
rect 19996 10112 20024 10208
rect 18380 10084 18828 10112
rect 18380 10072 18386 10084
rect 3602 10004 3608 10056
rect 3660 10004 3666 10056
rect 18598 10004 18604 10056
rect 18656 10004 18662 10056
rect 18800 10053 18828 10084
rect 19444 10084 20024 10112
rect 19444 10053 19472 10084
rect 20548 10053 20576 10208
rect 20625 10115 20683 10121
rect 20625 10081 20637 10115
rect 20671 10112 20683 10115
rect 20824 10112 20852 10208
rect 20901 10183 20959 10189
rect 20901 10149 20913 10183
rect 20947 10180 20959 10183
rect 20947 10152 27660 10180
rect 20947 10149 20959 10152
rect 20901 10143 20959 10149
rect 20671 10084 20852 10112
rect 20671 10081 20683 10084
rect 20625 10075 20683 10081
rect 22554 10072 22560 10124
rect 22612 10112 22618 10124
rect 23566 10112 23572 10124
rect 22612 10084 23572 10112
rect 22612 10072 22618 10084
rect 23566 10072 23572 10084
rect 23624 10072 23630 10124
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10013 18843 10047
rect 18785 10007 18843 10013
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10013 19487 10047
rect 19429 10007 19487 10013
rect 19613 10047 19671 10053
rect 19613 10013 19625 10047
rect 19659 10013 19671 10047
rect 19613 10007 19671 10013
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 1394 9936 1400 9988
rect 1452 9976 1458 9988
rect 1857 9979 1915 9985
rect 1857 9976 1869 9979
rect 1452 9948 1869 9976
rect 1452 9936 1458 9948
rect 1857 9945 1869 9948
rect 1903 9945 1915 9979
rect 1857 9939 1915 9945
rect 2866 9936 2872 9988
rect 2924 9936 2930 9988
rect 18509 9979 18567 9985
rect 18509 9945 18521 9979
rect 18555 9976 18567 9979
rect 19628 9976 19656 10007
rect 22002 10004 22008 10056
rect 22060 10044 22066 10056
rect 22189 10047 22247 10053
rect 22189 10044 22201 10047
rect 22060 10016 22201 10044
rect 22060 10004 22066 10016
rect 22189 10013 22201 10016
rect 22235 10013 22247 10047
rect 22189 10007 22247 10013
rect 22462 10004 22468 10056
rect 22520 10004 22526 10056
rect 23658 10004 23664 10056
rect 23716 10044 23722 10056
rect 23845 10047 23903 10053
rect 23845 10044 23857 10047
rect 23716 10016 23857 10044
rect 23716 10004 23722 10016
rect 23845 10013 23857 10016
rect 23891 10044 23903 10047
rect 24026 10044 24032 10056
rect 23891 10016 24032 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 24118 10004 24124 10056
rect 24176 10004 24182 10056
rect 24213 10047 24271 10053
rect 24213 10013 24225 10047
rect 24259 10044 24271 10047
rect 25038 10044 25044 10056
rect 24259 10016 25044 10044
rect 24259 10013 24271 10016
rect 24213 10007 24271 10013
rect 25038 10004 25044 10016
rect 25096 10004 25102 10056
rect 25774 10004 25780 10056
rect 25832 10044 25838 10056
rect 26513 10047 26571 10053
rect 26513 10044 26525 10047
rect 25832 10016 26525 10044
rect 25832 10004 25838 10016
rect 26513 10013 26525 10016
rect 26559 10013 26571 10047
rect 26513 10007 26571 10013
rect 26973 10047 27031 10053
rect 26973 10013 26985 10047
rect 27019 10044 27031 10047
rect 27246 10044 27252 10056
rect 27019 10016 27252 10044
rect 27019 10013 27031 10016
rect 26973 10007 27031 10013
rect 18555 9948 21680 9976
rect 18555 9945 18567 9948
rect 18509 9939 18567 9945
rect 18598 9868 18604 9920
rect 18656 9908 18662 9920
rect 20346 9908 20352 9920
rect 18656 9880 20352 9908
rect 18656 9868 18662 9880
rect 20346 9868 20352 9880
rect 20404 9908 20410 9920
rect 21358 9908 21364 9920
rect 20404 9880 21364 9908
rect 20404 9868 20410 9880
rect 21358 9868 21364 9880
rect 21416 9908 21422 9920
rect 21545 9911 21603 9917
rect 21545 9908 21557 9911
rect 21416 9880 21557 9908
rect 21416 9868 21422 9880
rect 21545 9877 21557 9880
rect 21591 9877 21603 9911
rect 21652 9908 21680 9948
rect 23934 9936 23940 9988
rect 23992 9976 23998 9988
rect 24397 9979 24455 9985
rect 24397 9976 24409 9979
rect 23992 9948 24409 9976
rect 23992 9936 23998 9948
rect 24397 9945 24409 9948
rect 24443 9945 24455 9979
rect 24397 9939 24455 9945
rect 22830 9908 22836 9920
rect 21652 9880 22836 9908
rect 21545 9871 21603 9877
rect 22830 9868 22836 9880
rect 22888 9868 22894 9920
rect 22922 9868 22928 9920
rect 22980 9908 22986 9920
rect 24302 9908 24308 9920
rect 22980 9880 24308 9908
rect 22980 9868 22986 9880
rect 24302 9868 24308 9880
rect 24360 9868 24366 9920
rect 24412 9908 24440 9939
rect 24486 9936 24492 9988
rect 24544 9976 24550 9988
rect 24597 9979 24655 9985
rect 24597 9976 24609 9979
rect 24544 9948 24609 9976
rect 24544 9936 24550 9948
rect 24597 9945 24609 9948
rect 24643 9945 24655 9979
rect 24597 9939 24655 9945
rect 25130 9936 25136 9988
rect 25188 9976 25194 9988
rect 26142 9976 26148 9988
rect 25188 9948 26148 9976
rect 25188 9936 25194 9948
rect 26142 9936 26148 9948
rect 26200 9976 26206 9988
rect 26200 9948 26358 9976
rect 26200 9936 26206 9948
rect 25041 9911 25099 9917
rect 25041 9908 25053 9911
rect 24412 9880 25053 9908
rect 25041 9877 25053 9880
rect 25087 9908 25099 9911
rect 25409 9911 25467 9917
rect 25409 9908 25421 9911
rect 25087 9880 25421 9908
rect 25087 9877 25099 9880
rect 25041 9871 25099 9877
rect 25409 9877 25421 9880
rect 25455 9877 25467 9911
rect 25409 9871 25467 9877
rect 25958 9868 25964 9920
rect 26016 9908 26022 9920
rect 26988 9908 27016 10007
rect 27246 10004 27252 10016
rect 27304 10004 27310 10056
rect 27632 9976 27660 10152
rect 28074 10072 28080 10124
rect 28132 10072 28138 10124
rect 28184 10053 28212 10220
rect 28902 10208 28908 10260
rect 28960 10248 28966 10260
rect 28997 10251 29055 10257
rect 28997 10248 29009 10251
rect 28960 10220 29009 10248
rect 28960 10208 28966 10220
rect 28997 10217 29009 10220
rect 29043 10217 29055 10251
rect 28997 10211 29055 10217
rect 28169 10047 28227 10053
rect 28169 10013 28181 10047
rect 28215 10013 28227 10047
rect 29012 10044 29040 10211
rect 31294 10208 31300 10260
rect 31352 10208 31358 10260
rect 31386 10208 31392 10260
rect 31444 10208 31450 10260
rect 31938 10208 31944 10260
rect 31996 10248 32002 10260
rect 32493 10251 32551 10257
rect 32493 10248 32505 10251
rect 31996 10220 32505 10248
rect 31996 10208 32002 10220
rect 32493 10217 32505 10220
rect 32539 10217 32551 10251
rect 32493 10211 32551 10217
rect 31404 10112 31432 10208
rect 31956 10180 31984 10208
rect 31864 10152 31984 10180
rect 31481 10115 31539 10121
rect 31481 10112 31493 10115
rect 31404 10084 31493 10112
rect 31481 10081 31493 10084
rect 31527 10081 31539 10115
rect 31481 10075 31539 10081
rect 29181 10047 29239 10053
rect 29181 10044 29193 10047
rect 29012 10016 29193 10044
rect 28169 10007 28227 10013
rect 29181 10013 29193 10016
rect 29227 10013 29239 10047
rect 29181 10007 29239 10013
rect 29362 10004 29368 10056
rect 29420 10044 29426 10056
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 29420 10016 29561 10044
rect 29420 10004 29426 10016
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 31110 10004 31116 10056
rect 31168 10044 31174 10056
rect 31573 10047 31631 10053
rect 31573 10044 31585 10047
rect 31168 10016 31585 10044
rect 31168 10004 31174 10016
rect 31573 10013 31585 10016
rect 31619 10013 31631 10047
rect 31864 10044 31892 10152
rect 31941 10115 31999 10121
rect 31941 10081 31953 10115
rect 31987 10112 31999 10115
rect 33045 10115 33103 10121
rect 33045 10112 33057 10115
rect 31987 10084 33057 10112
rect 31987 10081 31999 10084
rect 31941 10075 31999 10081
rect 33045 10081 33057 10084
rect 33091 10081 33103 10115
rect 33045 10075 33103 10081
rect 34072 10084 34744 10112
rect 34072 10056 34100 10084
rect 32033 10047 32091 10053
rect 32033 10044 32045 10047
rect 31864 10016 32045 10044
rect 31573 10007 31631 10013
rect 32033 10013 32045 10016
rect 32079 10013 32091 10047
rect 32033 10007 32091 10013
rect 32214 10004 32220 10056
rect 32272 10004 32278 10056
rect 32766 10004 32772 10056
rect 32824 10004 32830 10056
rect 34054 10004 34060 10056
rect 34112 10004 34118 10056
rect 34716 10053 34744 10084
rect 34701 10047 34759 10053
rect 34701 10013 34713 10047
rect 34747 10013 34759 10047
rect 34701 10007 34759 10013
rect 29825 9979 29883 9985
rect 29825 9976 29837 9979
rect 27632 9948 29837 9976
rect 29825 9945 29837 9948
rect 29871 9945 29883 9979
rect 29825 9939 29883 9945
rect 30098 9936 30104 9988
rect 30156 9976 30162 9988
rect 32232 9976 32260 10004
rect 34793 9979 34851 9985
rect 34793 9976 34805 9979
rect 30156 9948 30314 9976
rect 32232 9948 32812 9976
rect 34270 9948 34805 9976
rect 30156 9936 30162 9948
rect 32784 9920 32812 9948
rect 34793 9945 34805 9948
rect 34839 9945 34851 9979
rect 34793 9939 34851 9945
rect 26016 9880 27016 9908
rect 26016 9868 26022 9880
rect 28534 9868 28540 9920
rect 28592 9868 28598 9920
rect 29270 9868 29276 9920
rect 29328 9868 29334 9920
rect 32214 9868 32220 9920
rect 32272 9868 32278 9920
rect 32766 9868 32772 9920
rect 32824 9868 32830 9920
rect 34514 9868 34520 9920
rect 34572 9868 34578 9920
rect 1104 9818 35236 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 35236 9818
rect 1104 9744 35236 9766
rect 2866 9664 2872 9716
rect 2924 9664 2930 9716
rect 3234 9704 3240 9716
rect 3195 9676 3240 9704
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 17218 9664 17224 9716
rect 17276 9704 17282 9716
rect 22922 9704 22928 9716
rect 17276 9676 22928 9704
rect 17276 9664 17282 9676
rect 22922 9664 22928 9676
rect 22980 9664 22986 9716
rect 23014 9664 23020 9716
rect 23072 9704 23078 9716
rect 23109 9707 23167 9713
rect 23109 9704 23121 9707
rect 23072 9676 23121 9704
rect 23072 9664 23078 9676
rect 23109 9673 23121 9676
rect 23155 9673 23167 9707
rect 23109 9667 23167 9673
rect 24026 9664 24032 9716
rect 24084 9664 24090 9716
rect 24118 9664 24124 9716
rect 24176 9704 24182 9716
rect 24397 9707 24455 9713
rect 24397 9704 24409 9707
rect 24176 9676 24409 9704
rect 24176 9664 24182 9676
rect 24397 9673 24409 9676
rect 24443 9673 24455 9707
rect 26234 9704 26240 9716
rect 24397 9667 24455 9673
rect 24872 9676 26240 9704
rect 2777 9639 2835 9645
rect 2777 9605 2789 9639
rect 2823 9636 2835 9639
rect 2884 9636 2912 9664
rect 2823 9608 2912 9636
rect 2823 9605 2835 9608
rect 2777 9599 2835 9605
rect 2869 9571 2927 9577
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3252 9568 3280 9664
rect 18325 9639 18383 9645
rect 18325 9605 18337 9639
rect 18371 9636 18383 9639
rect 18598 9636 18604 9648
rect 18371 9608 18604 9636
rect 18371 9605 18383 9608
rect 18325 9599 18383 9605
rect 18598 9596 18604 9608
rect 18656 9596 18662 9648
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 22373 9639 22431 9645
rect 22373 9636 22385 9639
rect 22152 9608 22385 9636
rect 22152 9596 22158 9608
rect 22373 9605 22385 9608
rect 22419 9605 22431 9639
rect 22373 9599 22431 9605
rect 2915 9540 3280 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 22186 9528 22192 9580
rect 22244 9528 22250 9580
rect 22388 9568 22416 9599
rect 22462 9596 22468 9648
rect 22520 9636 22526 9648
rect 22833 9639 22891 9645
rect 22833 9636 22845 9639
rect 22520 9608 22845 9636
rect 22520 9596 22526 9608
rect 22833 9605 22845 9608
rect 22879 9636 22891 9639
rect 23290 9636 23296 9648
rect 22879 9608 23296 9636
rect 22879 9605 22891 9608
rect 22833 9599 22891 9605
rect 23290 9596 23296 9608
rect 23348 9636 23354 9648
rect 24136 9636 24164 9664
rect 23348 9608 24164 9636
rect 23348 9596 23354 9608
rect 24302 9596 24308 9648
rect 24360 9636 24366 9648
rect 24872 9636 24900 9676
rect 26234 9664 26240 9676
rect 26292 9704 26298 9716
rect 26602 9704 26608 9716
rect 26292 9676 26608 9704
rect 26292 9664 26298 9676
rect 26602 9664 26608 9676
rect 26660 9664 26666 9716
rect 28074 9664 28080 9716
rect 28132 9664 28138 9716
rect 24360 9608 24900 9636
rect 24360 9596 24366 9608
rect 27154 9596 27160 9648
rect 27212 9636 27218 9648
rect 27433 9639 27491 9645
rect 27212 9608 27384 9636
rect 27212 9596 27218 9608
rect 23014 9568 23020 9580
rect 22388 9540 23020 9568
rect 23014 9528 23020 9540
rect 23072 9568 23078 9580
rect 23385 9571 23443 9577
rect 23385 9568 23397 9571
rect 23072 9540 23397 9568
rect 23072 9528 23078 9540
rect 23385 9537 23397 9540
rect 23431 9537 23443 9571
rect 23385 9531 23443 9537
rect 23661 9571 23719 9577
rect 23661 9537 23673 9571
rect 23707 9568 23719 9571
rect 23934 9568 23940 9580
rect 23707 9540 23940 9568
rect 23707 9537 23719 9540
rect 23661 9531 23719 9537
rect 23934 9528 23940 9540
rect 23992 9528 23998 9580
rect 24026 9528 24032 9580
rect 24084 9568 24090 9580
rect 27356 9577 27384 9608
rect 27433 9605 27445 9639
rect 27479 9636 27491 9639
rect 28092 9636 28120 9664
rect 27479 9608 28120 9636
rect 27479 9605 27491 9608
rect 27433 9599 27491 9605
rect 28534 9596 28540 9648
rect 28592 9636 28598 9648
rect 28813 9639 28871 9645
rect 28813 9636 28825 9639
rect 28592 9608 28825 9636
rect 28592 9596 28598 9608
rect 28813 9605 28825 9608
rect 28859 9605 28871 9639
rect 28813 9599 28871 9605
rect 29270 9596 29276 9648
rect 29328 9596 29334 9648
rect 24765 9571 24823 9577
rect 24765 9568 24777 9571
rect 24084 9540 24777 9568
rect 24084 9528 24090 9540
rect 24765 9537 24777 9540
rect 24811 9537 24823 9571
rect 24765 9531 24823 9537
rect 27341 9571 27399 9577
rect 27341 9537 27353 9571
rect 27387 9537 27399 9571
rect 27341 9531 27399 9537
rect 27522 9528 27528 9580
rect 27580 9528 27586 9580
rect 31294 9528 31300 9580
rect 31352 9568 31358 9580
rect 32309 9571 32367 9577
rect 32309 9568 32321 9571
rect 31352 9540 32321 9568
rect 31352 9528 31358 9540
rect 32309 9537 32321 9540
rect 32355 9537 32367 9571
rect 32309 9531 32367 9537
rect 32766 9528 32772 9580
rect 32824 9528 32830 9580
rect 34514 9528 34520 9580
rect 34572 9568 34578 9580
rect 34701 9571 34759 9577
rect 34701 9568 34713 9571
rect 34572 9540 34713 9568
rect 34572 9528 34578 9540
rect 34701 9537 34713 9540
rect 34747 9537 34759 9571
rect 34701 9531 34759 9537
rect 34790 9528 34796 9580
rect 34848 9528 34854 9580
rect 22097 9503 22155 9509
rect 22097 9469 22109 9503
rect 22143 9500 22155 9503
rect 22204 9500 22232 9528
rect 22143 9472 22232 9500
rect 28445 9503 28503 9509
rect 22143 9469 22155 9472
rect 22097 9463 22155 9469
rect 28445 9469 28457 9503
rect 28491 9500 28503 9503
rect 28537 9503 28595 9509
rect 28537 9500 28549 9503
rect 28491 9472 28549 9500
rect 28491 9469 28503 9472
rect 28445 9463 28503 9469
rect 28537 9469 28549 9472
rect 28583 9500 28595 9503
rect 29362 9500 29368 9512
rect 28583 9472 29368 9500
rect 28583 9469 28595 9472
rect 28537 9463 28595 9469
rect 29362 9460 29368 9472
rect 29420 9460 29426 9512
rect 30285 9503 30343 9509
rect 30285 9469 30297 9503
rect 30331 9500 30343 9503
rect 31110 9500 31116 9512
rect 30331 9472 31116 9500
rect 30331 9469 30343 9472
rect 30285 9463 30343 9469
rect 31110 9460 31116 9472
rect 31168 9460 31174 9512
rect 32214 9460 32220 9512
rect 32272 9460 32278 9512
rect 34425 9503 34483 9509
rect 34425 9469 34437 9503
rect 34471 9500 34483 9503
rect 34808 9500 34836 9528
rect 34471 9472 34836 9500
rect 34471 9469 34483 9472
rect 34425 9463 34483 9469
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 32582 9324 32588 9376
rect 32640 9324 32646 9376
rect 32950 9324 32956 9376
rect 33008 9324 33014 9376
rect 1104 9274 35248 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 35248 9274
rect 1104 9200 35248 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 1670 9160 1676 9172
rect 1627 9132 1676 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 1670 9120 1676 9132
rect 1728 9120 1734 9172
rect 23014 9120 23020 9172
rect 23072 9120 23078 9172
rect 23477 9163 23535 9169
rect 23477 9129 23489 9163
rect 23523 9160 23535 9163
rect 23934 9160 23940 9172
rect 23523 9132 23940 9160
rect 23523 9129 23535 9132
rect 23477 9123 23535 9129
rect 23934 9120 23940 9132
rect 23992 9120 23998 9172
rect 32950 9120 32956 9172
rect 33008 9120 33014 9172
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 27709 9095 27767 9101
rect 27709 9092 27721 9095
rect 10100 9064 27721 9092
rect 10100 9052 10106 9064
rect 27709 9061 27721 9064
rect 27755 9092 27767 9095
rect 27755 9064 31754 9092
rect 27755 9061 27767 9064
rect 27709 9055 27767 9061
rect 31726 9024 31754 9064
rect 31726 8996 32812 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 23750 8916 23756 8968
rect 23808 8956 23814 8968
rect 24489 8959 24547 8965
rect 24489 8956 24501 8959
rect 23808 8928 24501 8956
rect 23808 8916 23814 8928
rect 24489 8925 24501 8928
rect 24535 8925 24547 8959
rect 24489 8919 24547 8925
rect 25038 8916 25044 8968
rect 25096 8916 25102 8968
rect 26234 8916 26240 8968
rect 26292 8956 26298 8968
rect 26421 8959 26479 8965
rect 26421 8956 26433 8959
rect 26292 8928 26433 8956
rect 26292 8916 26298 8928
rect 26421 8925 26433 8928
rect 26467 8956 26479 8959
rect 28445 8959 28503 8965
rect 28445 8956 28457 8959
rect 26467 8928 28457 8956
rect 26467 8925 26479 8928
rect 26421 8919 26479 8925
rect 28445 8925 28457 8928
rect 28491 8925 28503 8959
rect 28445 8919 28503 8925
rect 25964 8900 26016 8906
rect 32784 8888 32812 8996
rect 32861 8959 32919 8965
rect 32861 8925 32873 8959
rect 32907 8956 32919 8959
rect 32968 8956 32996 9120
rect 32907 8928 32996 8956
rect 33413 8959 33471 8965
rect 32907 8925 32919 8928
rect 32861 8919 32919 8925
rect 33413 8925 33425 8959
rect 33459 8956 33471 8959
rect 33873 8959 33931 8965
rect 33873 8956 33885 8959
rect 33459 8928 33885 8956
rect 33459 8925 33471 8928
rect 33413 8919 33471 8925
rect 33873 8925 33885 8928
rect 33919 8956 33931 8959
rect 34054 8956 34060 8968
rect 33919 8928 34060 8956
rect 33919 8925 33931 8928
rect 33873 8919 33931 8925
rect 33428 8888 33456 8919
rect 34054 8916 34060 8928
rect 34112 8916 34118 8968
rect 32784 8860 33456 8888
rect 25964 8842 26016 8848
rect 33042 8780 33048 8832
rect 33100 8780 33106 8832
rect 33502 8780 33508 8832
rect 33560 8780 33566 8832
rect 1104 8730 35236 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 35236 8730
rect 1104 8656 35236 8678
rect 32582 8576 32588 8628
rect 32640 8616 32646 8628
rect 32640 8588 32812 8616
rect 32640 8576 32646 8588
rect 26234 8508 26240 8560
rect 26292 8548 26298 8560
rect 27157 8551 27215 8557
rect 27157 8548 27169 8551
rect 26292 8520 27169 8548
rect 26292 8508 26298 8520
rect 27157 8517 27169 8520
rect 27203 8517 27215 8551
rect 27157 8511 27215 8517
rect 32401 8551 32459 8557
rect 32401 8517 32413 8551
rect 32447 8548 32459 8551
rect 32674 8548 32680 8560
rect 32447 8520 32680 8548
rect 32447 8517 32459 8520
rect 32401 8511 32459 8517
rect 27798 8440 27804 8492
rect 27856 8440 27862 8492
rect 32416 8480 32444 8511
rect 32674 8508 32680 8520
rect 32732 8508 32738 8560
rect 32784 8557 32812 8588
rect 34054 8576 34060 8628
rect 34112 8576 34118 8628
rect 32769 8551 32827 8557
rect 32769 8517 32781 8551
rect 32815 8517 32827 8551
rect 32769 8511 32827 8517
rect 33502 8508 33508 8560
rect 33560 8508 33566 8560
rect 32493 8483 32551 8489
rect 32493 8480 32505 8483
rect 32416 8452 32505 8480
rect 32493 8449 32505 8452
rect 32539 8449 32551 8483
rect 34072 8480 34100 8576
rect 34517 8483 34575 8489
rect 34517 8480 34529 8483
rect 34072 8452 34529 8480
rect 32493 8443 32551 8449
rect 34517 8449 34529 8452
rect 34563 8480 34575 8483
rect 34793 8483 34851 8489
rect 34793 8480 34805 8483
rect 34563 8452 34805 8480
rect 34563 8449 34575 8452
rect 34517 8443 34575 8449
rect 34793 8449 34805 8452
rect 34839 8449 34851 8483
rect 34793 8443 34851 8449
rect 34238 8304 34244 8356
rect 34296 8304 34302 8356
rect 34422 8236 34428 8288
rect 34480 8236 34486 8288
rect 1104 8186 35248 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 35248 8186
rect 1104 8112 35248 8134
rect 32674 8032 32680 8084
rect 32732 8032 32738 8084
rect 32692 7936 32720 8032
rect 32769 7939 32827 7945
rect 32769 7936 32781 7939
rect 32692 7908 32781 7936
rect 32769 7905 32781 7908
rect 32815 7905 32827 7939
rect 32769 7899 32827 7905
rect 33042 7896 33048 7948
rect 33100 7896 33106 7948
rect 34422 7868 34428 7880
rect 34178 7840 34428 7868
rect 34422 7828 34428 7840
rect 34480 7828 34486 7880
rect 34514 7692 34520 7744
rect 34572 7692 34578 7744
rect 1104 7642 35236 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 35236 7642
rect 1104 7568 35236 7590
rect 34606 7352 34612 7404
rect 34664 7392 34670 7404
rect 34701 7395 34759 7401
rect 34701 7392 34713 7395
rect 34664 7364 34713 7392
rect 34664 7352 34670 7364
rect 34701 7361 34713 7364
rect 34747 7361 34759 7395
rect 34701 7355 34759 7361
rect 34790 7352 34796 7404
rect 34848 7352 34854 7404
rect 34425 7327 34483 7333
rect 34425 7293 34437 7327
rect 34471 7324 34483 7327
rect 34808 7324 34836 7352
rect 34471 7296 34836 7324
rect 34471 7293 34483 7296
rect 34425 7287 34483 7293
rect 1104 7098 35248 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 35248 7098
rect 1104 7024 35248 7046
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 992 6752 1409 6780
rect 992 6740 998 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1486 6604 1492 6656
rect 1544 6644 1550 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 1544 6616 1593 6644
rect 1544 6604 1550 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 1581 6607 1639 6613
rect 1104 6554 35236 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 35236 6554
rect 1104 6480 35236 6502
rect 1104 6010 35248 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 35248 6010
rect 1104 5936 35248 5958
rect 34057 5763 34115 5769
rect 34057 5729 34069 5763
rect 34103 5729 34115 5763
rect 34057 5723 34115 5729
rect 34072 5636 34100 5723
rect 34330 5652 34336 5704
rect 34388 5652 34394 5704
rect 34054 5584 34060 5636
rect 34112 5584 34118 5636
rect 1104 5466 35236 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 35236 5466
rect 1104 5392 35236 5414
rect 1104 4922 35248 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 35248 4922
rect 1104 4848 35248 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 2958 4808 2964 4820
rect 1627 4780 2964 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1104 4378 35236 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 35236 4378
rect 1104 4304 35236 4326
rect 1104 3834 35248 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 35248 3834
rect 1104 3760 35248 3782
rect 34057 3587 34115 3593
rect 34057 3553 34069 3587
rect 34103 3584 34115 3587
rect 34103 3556 34652 3584
rect 34103 3553 34115 3556
rect 34057 3547 34115 3553
rect 34425 3519 34483 3525
rect 34425 3485 34437 3519
rect 34471 3516 34483 3519
rect 34514 3516 34520 3528
rect 34471 3488 34520 3516
rect 34471 3485 34483 3488
rect 34425 3479 34483 3485
rect 34514 3476 34520 3488
rect 34572 3476 34578 3528
rect 34624 3460 34652 3556
rect 34606 3408 34612 3460
rect 34664 3408 34670 3460
rect 1104 3290 35236 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 35236 3290
rect 1104 3216 35236 3238
rect 1104 2746 35248 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 35248 2746
rect 1104 2672 35248 2694
rect 1394 2592 1400 2644
rect 1452 2632 1458 2644
rect 1581 2635 1639 2641
rect 1581 2632 1593 2635
rect 1452 2604 1593 2632
rect 1452 2592 1458 2604
rect 1581 2601 1593 2604
rect 1627 2601 1639 2635
rect 1581 2595 1639 2601
rect 27525 2635 27583 2641
rect 27525 2601 27537 2635
rect 27571 2632 27583 2635
rect 27798 2632 27804 2644
rect 27571 2604 27804 2632
rect 27571 2601 27583 2604
rect 27525 2595 27583 2601
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 9582 2456 9588 2508
rect 9640 2456 9646 2508
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 27338 2388 27344 2440
rect 27396 2388 27402 2440
rect 1104 2202 35236 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 35236 2202
rect 1104 2128 35236 2150
<< via1 >>
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 940 36116 992 36168
rect 33140 36159 33192 36168
rect 33140 36125 33149 36159
rect 33149 36125 33183 36159
rect 33183 36125 33192 36159
rect 33140 36116 33192 36125
rect 34336 36091 34388 36100
rect 34336 36057 34345 36091
rect 34345 36057 34379 36091
rect 34379 36057 34388 36091
rect 34336 36048 34388 36057
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 940 35028 992 35080
rect 1860 34892 1912 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 34520 33983 34572 33992
rect 34520 33949 34529 33983
rect 34529 33949 34563 33983
rect 34563 33949 34572 33983
rect 34520 33940 34572 33949
rect 34612 33872 34664 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 940 32852 992 32904
rect 4068 32716 4120 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 34428 31807 34480 31816
rect 34428 31773 34437 31807
rect 34437 31773 34471 31807
rect 34471 31773 34480 31807
rect 34428 31764 34480 31773
rect 34060 31696 34112 31748
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 2872 30540 2924 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 34612 29520 34664 29572
rect 34796 29452 34848 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 34520 28747 34572 28756
rect 34520 28713 34529 28747
rect 34529 28713 34563 28747
rect 34563 28713 34572 28747
rect 34520 28704 34572 28713
rect 940 28500 992 28552
rect 19984 28500 20036 28552
rect 20352 28568 20404 28620
rect 20168 28432 20220 28484
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 19340 28364 19392 28416
rect 19892 28407 19944 28416
rect 19892 28373 19901 28407
rect 19901 28373 19935 28407
rect 19935 28373 19944 28407
rect 19892 28364 19944 28373
rect 19984 28364 20036 28416
rect 34152 28500 34204 28552
rect 33048 28475 33100 28484
rect 33048 28441 33057 28475
rect 33057 28441 33091 28475
rect 33091 28441 33100 28475
rect 33048 28432 33100 28441
rect 21548 28407 21600 28416
rect 21548 28373 21557 28407
rect 21557 28373 21591 28407
rect 21591 28373 21600 28407
rect 21548 28364 21600 28373
rect 32588 28407 32640 28416
rect 32588 28373 32597 28407
rect 32597 28373 32631 28407
rect 32631 28373 32640 28407
rect 32588 28364 32640 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 19800 28160 19852 28212
rect 19340 28024 19392 28076
rect 21456 28160 21508 28212
rect 21548 28160 21600 28212
rect 20076 28092 20128 28144
rect 21088 28067 21140 28076
rect 21088 28033 21097 28067
rect 21097 28033 21131 28067
rect 21131 28033 21140 28067
rect 21088 28024 21140 28033
rect 19432 27956 19484 28008
rect 19524 27999 19576 28008
rect 19524 27965 19533 27999
rect 19533 27965 19567 27999
rect 19567 27965 19576 27999
rect 19524 27956 19576 27965
rect 20076 27999 20128 28008
rect 20076 27965 20085 27999
rect 20085 27965 20119 27999
rect 20119 27965 20128 27999
rect 20076 27956 20128 27965
rect 20168 27999 20220 28008
rect 20168 27965 20177 27999
rect 20177 27965 20211 27999
rect 20211 27965 20220 27999
rect 20168 27956 20220 27965
rect 34428 28203 34480 28212
rect 34428 28169 34437 28203
rect 34437 28169 34471 28203
rect 34471 28169 34480 28203
rect 34428 28160 34480 28169
rect 22560 28067 22612 28076
rect 22560 28033 22569 28067
rect 22569 28033 22603 28067
rect 22603 28033 22612 28067
rect 22560 28024 22612 28033
rect 33692 28092 33744 28144
rect 32956 27999 33008 28008
rect 32956 27965 32965 27999
rect 32965 27965 32999 27999
rect 32999 27965 33008 27999
rect 32956 27956 33008 27965
rect 19340 27863 19392 27872
rect 19340 27829 19349 27863
rect 19349 27829 19383 27863
rect 19383 27829 19392 27863
rect 19340 27820 19392 27829
rect 20812 27863 20864 27872
rect 20812 27829 20821 27863
rect 20821 27829 20855 27863
rect 20855 27829 20864 27863
rect 20812 27820 20864 27829
rect 22836 27863 22888 27872
rect 22836 27829 22845 27863
rect 22845 27829 22879 27863
rect 22879 27829 22888 27863
rect 22836 27820 22888 27829
rect 30656 27863 30708 27872
rect 30656 27829 30665 27863
rect 30665 27829 30699 27863
rect 30699 27829 30708 27863
rect 30656 27820 30708 27829
rect 30932 27863 30984 27872
rect 30932 27829 30941 27863
rect 30941 27829 30975 27863
rect 30975 27829 30984 27863
rect 30932 27820 30984 27829
rect 31024 27820 31076 27872
rect 31760 27863 31812 27872
rect 31760 27829 31769 27863
rect 31769 27829 31803 27863
rect 31803 27829 31812 27863
rect 32588 27863 32640 27872
rect 31760 27820 31812 27829
rect 32588 27829 32597 27863
rect 32597 27829 32631 27863
rect 32631 27829 32640 27863
rect 32588 27820 32640 27829
rect 34704 27863 34756 27872
rect 34704 27829 34713 27863
rect 34713 27829 34747 27863
rect 34747 27829 34756 27863
rect 34704 27820 34756 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 2872 27616 2924 27668
rect 19432 27616 19484 27668
rect 19524 27548 19576 27600
rect 14924 27480 14976 27532
rect 14832 27455 14884 27464
rect 14832 27421 14841 27455
rect 14841 27421 14875 27455
rect 14875 27421 14884 27455
rect 14832 27412 14884 27421
rect 15108 27455 15160 27464
rect 15108 27421 15117 27455
rect 15117 27421 15151 27455
rect 15151 27421 15160 27455
rect 15108 27412 15160 27421
rect 16764 27480 16816 27532
rect 20076 27616 20128 27668
rect 21456 27616 21508 27668
rect 22836 27616 22888 27668
rect 33692 27659 33744 27668
rect 33692 27625 33701 27659
rect 33701 27625 33735 27659
rect 33735 27625 33744 27659
rect 33692 27616 33744 27625
rect 34152 27659 34204 27668
rect 34152 27625 34161 27659
rect 34161 27625 34195 27659
rect 34195 27625 34204 27659
rect 34152 27616 34204 27625
rect 4160 27344 4212 27396
rect 17316 27412 17368 27464
rect 20168 27455 20220 27464
rect 20168 27421 20177 27455
rect 20177 27421 20211 27455
rect 20211 27421 20220 27455
rect 20168 27412 20220 27421
rect 23388 27455 23440 27464
rect 3608 27276 3660 27328
rect 5540 27319 5592 27328
rect 5540 27285 5549 27319
rect 5549 27285 5583 27319
rect 5583 27285 5592 27319
rect 5540 27276 5592 27285
rect 5816 27319 5868 27328
rect 5816 27285 5825 27319
rect 5825 27285 5859 27319
rect 5859 27285 5868 27319
rect 5816 27276 5868 27285
rect 15660 27319 15712 27328
rect 15660 27285 15669 27319
rect 15669 27285 15703 27319
rect 15703 27285 15712 27319
rect 15660 27276 15712 27285
rect 15936 27276 15988 27328
rect 16856 27276 16908 27328
rect 17500 27319 17552 27328
rect 17500 27285 17509 27319
rect 17509 27285 17543 27319
rect 17543 27285 17552 27319
rect 17500 27276 17552 27285
rect 17960 27276 18012 27328
rect 18512 27319 18564 27328
rect 18512 27285 18521 27319
rect 18521 27285 18555 27319
rect 18555 27285 18564 27319
rect 18512 27276 18564 27285
rect 18696 27276 18748 27328
rect 21456 27276 21508 27328
rect 23388 27421 23397 27455
rect 23397 27421 23431 27455
rect 23431 27421 23440 27455
rect 23388 27412 23440 27421
rect 23480 27455 23532 27464
rect 23480 27421 23489 27455
rect 23489 27421 23523 27455
rect 23523 27421 23532 27455
rect 23480 27412 23532 27421
rect 23664 27523 23716 27532
rect 23664 27489 23673 27523
rect 23673 27489 23707 27523
rect 23707 27489 23716 27523
rect 23664 27480 23716 27489
rect 25964 27344 26016 27396
rect 29736 27455 29788 27464
rect 29736 27421 29745 27455
rect 29745 27421 29779 27455
rect 29779 27421 29788 27455
rect 29736 27412 29788 27421
rect 30656 27455 30708 27464
rect 30656 27421 30665 27455
rect 30665 27421 30699 27455
rect 30699 27421 30708 27455
rect 30656 27412 30708 27421
rect 30840 27523 30892 27532
rect 30840 27489 30849 27523
rect 30849 27489 30883 27523
rect 30883 27489 30892 27523
rect 30840 27480 30892 27489
rect 33140 27591 33192 27600
rect 33140 27557 33149 27591
rect 33149 27557 33183 27591
rect 33183 27557 33192 27591
rect 33140 27548 33192 27557
rect 31024 27455 31076 27464
rect 31024 27421 31033 27455
rect 31033 27421 31067 27455
rect 31067 27421 31076 27455
rect 31024 27412 31076 27421
rect 31208 27344 31260 27396
rect 26700 27276 26752 27328
rect 27068 27319 27120 27328
rect 27068 27285 27077 27319
rect 27077 27285 27111 27319
rect 27111 27285 27120 27319
rect 27068 27276 27120 27285
rect 27252 27319 27304 27328
rect 27252 27285 27261 27319
rect 27261 27285 27295 27319
rect 27295 27285 27304 27319
rect 27252 27276 27304 27285
rect 30012 27276 30064 27328
rect 30840 27319 30892 27328
rect 30840 27285 30849 27319
rect 30849 27285 30883 27319
rect 30883 27285 30892 27319
rect 30840 27276 30892 27285
rect 33416 27455 33468 27464
rect 33416 27421 33425 27455
rect 33425 27421 33459 27455
rect 33459 27421 33468 27455
rect 33416 27412 33468 27421
rect 34152 27412 34204 27464
rect 34704 27480 34756 27532
rect 31760 27344 31812 27396
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4160 27115 4212 27124
rect 4160 27081 4169 27115
rect 4169 27081 4203 27115
rect 4203 27081 4212 27115
rect 4160 27072 4212 27081
rect 15660 27072 15712 27124
rect 15936 27047 15988 27056
rect 15936 27013 15945 27047
rect 15945 27013 15979 27047
rect 15979 27013 15988 27047
rect 15936 27004 15988 27013
rect 3608 26775 3660 26784
rect 3608 26741 3617 26775
rect 3617 26741 3651 26775
rect 3651 26741 3660 26775
rect 3608 26732 3660 26741
rect 14924 26936 14976 26988
rect 4988 26732 5040 26784
rect 16304 26979 16356 26988
rect 16304 26945 16313 26979
rect 16313 26945 16347 26979
rect 16347 26945 16356 26979
rect 16304 26936 16356 26945
rect 20076 27072 20128 27124
rect 19340 27047 19392 27056
rect 17316 26936 17368 26988
rect 17500 26936 17552 26988
rect 19340 27013 19349 27047
rect 19349 27013 19383 27047
rect 19383 27013 19392 27047
rect 19340 27004 19392 27013
rect 22560 27115 22612 27124
rect 22560 27081 22569 27115
rect 22569 27081 22603 27115
rect 22603 27081 22612 27115
rect 22560 27072 22612 27081
rect 23480 27072 23532 27124
rect 23664 27072 23716 27124
rect 25964 27115 26016 27124
rect 25964 27081 25973 27115
rect 25973 27081 26007 27115
rect 26007 27081 26016 27115
rect 25964 27072 26016 27081
rect 26700 27115 26752 27124
rect 26700 27081 26709 27115
rect 26709 27081 26743 27115
rect 26743 27081 26752 27115
rect 26700 27072 26752 27081
rect 27068 27072 27120 27124
rect 27252 27072 27304 27124
rect 29736 27072 29788 27124
rect 30840 27072 30892 27124
rect 32956 27072 33008 27124
rect 18420 26979 18472 26988
rect 18420 26945 18429 26979
rect 18429 26945 18463 26979
rect 18463 26945 18472 26979
rect 18420 26936 18472 26945
rect 18512 26936 18564 26988
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 18696 26936 18748 26945
rect 18788 26979 18840 26988
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 19524 26979 19576 26988
rect 19524 26945 19533 26979
rect 19533 26945 19567 26979
rect 19567 26945 19576 26979
rect 19524 26936 19576 26945
rect 15844 26843 15896 26852
rect 15844 26809 15853 26843
rect 15853 26809 15887 26843
rect 15887 26809 15896 26843
rect 15844 26800 15896 26809
rect 16856 26800 16908 26852
rect 19340 26868 19392 26920
rect 20076 26979 20128 26988
rect 20076 26945 20085 26979
rect 20085 26945 20119 26979
rect 20119 26945 20128 26979
rect 20076 26936 20128 26945
rect 20260 26979 20312 26988
rect 20260 26945 20269 26979
rect 20269 26945 20303 26979
rect 20303 26945 20312 26979
rect 20260 26936 20312 26945
rect 21640 27004 21692 27056
rect 20720 26936 20772 26988
rect 20812 26868 20864 26920
rect 21824 26979 21876 26988
rect 21824 26945 21833 26979
rect 21833 26945 21867 26979
rect 21867 26945 21876 26979
rect 21824 26936 21876 26945
rect 22284 26936 22336 26988
rect 23388 27004 23440 27056
rect 24860 26979 24912 26988
rect 24860 26945 24869 26979
rect 24869 26945 24903 26979
rect 24903 26945 24912 26979
rect 24860 26936 24912 26945
rect 26700 26936 26752 26988
rect 26884 26936 26936 26988
rect 15292 26732 15344 26784
rect 15384 26732 15436 26784
rect 19340 26775 19392 26784
rect 19340 26741 19349 26775
rect 19349 26741 19383 26775
rect 19383 26741 19392 26775
rect 19340 26732 19392 26741
rect 22376 26800 22428 26852
rect 23388 26800 23440 26852
rect 24308 26775 24360 26784
rect 24308 26741 24317 26775
rect 24317 26741 24351 26775
rect 24351 26741 24360 26775
rect 24308 26732 24360 26741
rect 28908 26775 28960 26784
rect 28908 26741 28917 26775
rect 28917 26741 28951 26775
rect 28951 26741 28960 26775
rect 28908 26732 28960 26741
rect 33416 27072 33468 27124
rect 31208 26936 31260 26988
rect 33692 26979 33744 26988
rect 33692 26945 33701 26979
rect 33701 26945 33735 26979
rect 33735 26945 33744 26979
rect 33692 26936 33744 26945
rect 34704 26979 34756 26988
rect 34704 26945 34713 26979
rect 34713 26945 34747 26979
rect 34747 26945 34756 26979
rect 34704 26936 34756 26945
rect 30932 26868 30984 26920
rect 29920 26732 29972 26784
rect 30012 26732 30064 26784
rect 33048 26732 33100 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5816 26571 5868 26580
rect 5816 26537 5825 26571
rect 5825 26537 5859 26571
rect 5859 26537 5868 26571
rect 5816 26528 5868 26537
rect 14832 26528 14884 26580
rect 16764 26528 16816 26580
rect 16856 26571 16908 26580
rect 16856 26537 16865 26571
rect 16865 26537 16899 26571
rect 16899 26537 16908 26571
rect 16856 26528 16908 26537
rect 17500 26528 17552 26580
rect 1676 26435 1728 26444
rect 1676 26401 1685 26435
rect 1685 26401 1719 26435
rect 1719 26401 1728 26435
rect 1676 26392 1728 26401
rect 2136 26256 2188 26308
rect 2044 26188 2096 26240
rect 3608 26392 3660 26444
rect 9312 26392 9364 26444
rect 9772 26392 9824 26444
rect 12992 26435 13044 26444
rect 12992 26401 13001 26435
rect 13001 26401 13035 26435
rect 13035 26401 13044 26435
rect 12992 26392 13044 26401
rect 15844 26392 15896 26444
rect 6828 26367 6880 26376
rect 6828 26333 6837 26367
rect 6837 26333 6871 26367
rect 6871 26333 6880 26367
rect 6828 26324 6880 26333
rect 3976 26256 4028 26308
rect 4068 26299 4120 26308
rect 4068 26265 4077 26299
rect 4077 26265 4111 26299
rect 4111 26265 4120 26299
rect 4068 26256 4120 26265
rect 4712 26256 4764 26308
rect 8300 26256 8352 26308
rect 12900 26367 12952 26376
rect 12900 26333 12909 26367
rect 12909 26333 12943 26367
rect 12943 26333 12952 26367
rect 12900 26324 12952 26333
rect 13636 26367 13688 26376
rect 13636 26333 13645 26367
rect 13645 26333 13679 26367
rect 13679 26333 13688 26367
rect 13636 26324 13688 26333
rect 14924 26324 14976 26376
rect 9312 26256 9364 26308
rect 9680 26256 9732 26308
rect 10692 26256 10744 26308
rect 15384 26299 15436 26308
rect 15384 26265 15393 26299
rect 15393 26265 15427 26299
rect 15427 26265 15436 26299
rect 15384 26256 15436 26265
rect 16304 26324 16356 26376
rect 15936 26256 15988 26308
rect 18420 26528 18472 26580
rect 19340 26528 19392 26580
rect 20076 26528 20128 26580
rect 20352 26571 20404 26580
rect 20352 26537 20361 26571
rect 20361 26537 20395 26571
rect 20395 26537 20404 26571
rect 20352 26528 20404 26537
rect 21456 26571 21508 26580
rect 21456 26537 21465 26571
rect 21465 26537 21499 26571
rect 21499 26537 21508 26571
rect 21456 26528 21508 26537
rect 21824 26528 21876 26580
rect 22100 26528 22152 26580
rect 22284 26571 22336 26580
rect 22284 26537 22293 26571
rect 22293 26537 22327 26571
rect 22327 26537 22336 26571
rect 22284 26528 22336 26537
rect 23388 26528 23440 26580
rect 24860 26528 24912 26580
rect 26884 26571 26936 26580
rect 26884 26537 26893 26571
rect 26893 26537 26927 26571
rect 26927 26537 26936 26571
rect 26884 26528 26936 26537
rect 30012 26528 30064 26580
rect 31024 26528 31076 26580
rect 34796 26528 34848 26580
rect 18052 26367 18104 26376
rect 18052 26333 18061 26367
rect 18061 26333 18095 26367
rect 18095 26333 18104 26367
rect 18052 26324 18104 26333
rect 18236 26367 18288 26376
rect 18236 26333 18245 26367
rect 18245 26333 18279 26367
rect 18279 26333 18288 26367
rect 18236 26324 18288 26333
rect 5540 26231 5592 26240
rect 5540 26197 5549 26231
rect 5549 26197 5583 26231
rect 5583 26197 5592 26231
rect 5540 26188 5592 26197
rect 13268 26231 13320 26240
rect 13268 26197 13277 26231
rect 13277 26197 13311 26231
rect 13311 26197 13320 26231
rect 13268 26188 13320 26197
rect 16396 26188 16448 26240
rect 19524 26392 19576 26444
rect 18788 26324 18840 26376
rect 19984 26324 20036 26376
rect 20444 26324 20496 26376
rect 21640 26392 21692 26444
rect 21548 26367 21600 26376
rect 21548 26333 21557 26367
rect 21557 26333 21591 26367
rect 21591 26333 21600 26367
rect 21548 26324 21600 26333
rect 22376 26324 22428 26376
rect 22652 26367 22704 26376
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 24308 26460 24360 26512
rect 26700 26460 26752 26512
rect 28908 26324 28960 26376
rect 30472 26299 30524 26308
rect 30472 26265 30481 26299
rect 30481 26265 30515 26299
rect 30515 26265 30524 26299
rect 30472 26256 30524 26265
rect 30564 26256 30616 26308
rect 20444 26188 20496 26240
rect 30748 26188 30800 26240
rect 31576 26188 31628 26240
rect 32588 26324 32640 26376
rect 32128 26188 32180 26240
rect 33048 26299 33100 26308
rect 33048 26265 33057 26299
rect 33057 26265 33091 26299
rect 33091 26265 33100 26299
rect 33048 26256 33100 26265
rect 34336 26256 34388 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 2136 25984 2188 26036
rect 4712 26027 4764 26036
rect 4712 25993 4721 26027
rect 4721 25993 4755 26027
rect 4755 25993 4764 26027
rect 4712 25984 4764 25993
rect 6828 25984 6880 26036
rect 9680 25984 9732 26036
rect 13636 25984 13688 26036
rect 1584 25916 1636 25968
rect 940 25848 992 25900
rect 1768 25644 1820 25696
rect 2044 25823 2096 25832
rect 2044 25789 2053 25823
rect 2053 25789 2087 25823
rect 2087 25789 2096 25823
rect 2044 25780 2096 25789
rect 2872 25644 2924 25696
rect 5908 25891 5960 25900
rect 5908 25857 5917 25891
rect 5917 25857 5951 25891
rect 5951 25857 5960 25891
rect 5908 25848 5960 25857
rect 12992 25916 13044 25968
rect 15660 25916 15712 25968
rect 6000 25780 6052 25832
rect 4620 25712 4672 25764
rect 12900 25891 12952 25900
rect 12900 25857 12909 25891
rect 12909 25857 12943 25891
rect 12943 25857 12952 25891
rect 12900 25848 12952 25857
rect 16120 25891 16172 25900
rect 13268 25780 13320 25832
rect 9864 25644 9916 25696
rect 16120 25857 16129 25891
rect 16129 25857 16163 25891
rect 16163 25857 16172 25891
rect 16120 25848 16172 25857
rect 15936 25823 15988 25832
rect 15936 25789 15945 25823
rect 15945 25789 15979 25823
rect 15979 25789 15988 25823
rect 18052 25984 18104 26036
rect 18696 25984 18748 26036
rect 19892 25984 19944 26036
rect 21088 25984 21140 26036
rect 21548 25984 21600 26036
rect 22192 26027 22244 26036
rect 22192 25993 22201 26027
rect 22201 25993 22235 26027
rect 22235 25993 22244 26027
rect 22192 25984 22244 25993
rect 22652 25984 22704 26036
rect 30564 25984 30616 26036
rect 33048 25984 33100 26036
rect 33692 25984 33744 26036
rect 34336 26027 34388 26036
rect 34336 25993 34345 26027
rect 34345 25993 34379 26027
rect 34379 25993 34388 26027
rect 34336 25984 34388 25993
rect 16764 25891 16816 25900
rect 16764 25857 16773 25891
rect 16773 25857 16807 25891
rect 16807 25857 16816 25891
rect 16764 25848 16816 25857
rect 15936 25780 15988 25789
rect 16580 25780 16632 25832
rect 18236 25916 18288 25968
rect 18880 25916 18932 25968
rect 17868 25823 17920 25832
rect 17868 25789 17877 25823
rect 17877 25789 17911 25823
rect 17911 25789 17920 25823
rect 17868 25780 17920 25789
rect 17960 25823 18012 25832
rect 17960 25789 17969 25823
rect 17969 25789 18003 25823
rect 18003 25789 18012 25823
rect 17960 25780 18012 25789
rect 19432 25848 19484 25900
rect 20076 25848 20128 25900
rect 20352 25891 20404 25900
rect 20352 25857 20361 25891
rect 20361 25857 20395 25891
rect 20395 25857 20404 25891
rect 20352 25848 20404 25857
rect 20536 25891 20588 25900
rect 20536 25857 20545 25891
rect 20545 25857 20579 25891
rect 20579 25857 20588 25891
rect 20536 25848 20588 25857
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 26700 25916 26752 25968
rect 22100 25848 22152 25857
rect 20444 25780 20496 25832
rect 21272 25823 21324 25832
rect 21272 25789 21281 25823
rect 21281 25789 21315 25823
rect 21315 25789 21324 25823
rect 21272 25780 21324 25789
rect 21916 25780 21968 25832
rect 23388 25848 23440 25900
rect 29920 25891 29972 25900
rect 29920 25857 29929 25891
rect 29929 25857 29963 25891
rect 29963 25857 29972 25891
rect 30656 25916 30708 25968
rect 29920 25848 29972 25857
rect 22376 25712 22428 25764
rect 34152 25891 34204 25900
rect 34152 25857 34161 25891
rect 34161 25857 34195 25891
rect 34195 25857 34204 25891
rect 34152 25848 34204 25857
rect 32128 25823 32180 25832
rect 32128 25789 32137 25823
rect 32137 25789 32171 25823
rect 32171 25789 32180 25823
rect 32128 25780 32180 25789
rect 32404 25823 32456 25832
rect 32404 25789 32413 25823
rect 32413 25789 32447 25823
rect 32447 25789 32456 25823
rect 32404 25780 32456 25789
rect 14648 25687 14700 25696
rect 14648 25653 14657 25687
rect 14657 25653 14691 25687
rect 14691 25653 14700 25687
rect 14648 25644 14700 25653
rect 15108 25687 15160 25696
rect 15108 25653 15117 25687
rect 15117 25653 15151 25687
rect 15151 25653 15160 25687
rect 15108 25644 15160 25653
rect 16304 25687 16356 25696
rect 16304 25653 16313 25687
rect 16313 25653 16347 25687
rect 16347 25653 16356 25687
rect 16304 25644 16356 25653
rect 17132 25687 17184 25696
rect 17132 25653 17141 25687
rect 17141 25653 17175 25687
rect 17175 25653 17184 25687
rect 17132 25644 17184 25653
rect 18972 25644 19024 25696
rect 20720 25687 20772 25696
rect 20720 25653 20729 25687
rect 20729 25653 20763 25687
rect 20763 25653 20772 25687
rect 20720 25644 20772 25653
rect 26884 25644 26936 25696
rect 27712 25687 27764 25696
rect 27712 25653 27721 25687
rect 27721 25653 27755 25687
rect 27755 25653 27764 25687
rect 27712 25644 27764 25653
rect 30104 25644 30156 25696
rect 31576 25644 31628 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 5908 25440 5960 25492
rect 8300 25440 8352 25492
rect 10692 25483 10744 25492
rect 10692 25449 10701 25483
rect 10701 25449 10735 25483
rect 10735 25449 10744 25483
rect 10692 25440 10744 25449
rect 16120 25440 16172 25492
rect 16764 25440 16816 25492
rect 18236 25440 18288 25492
rect 18972 25483 19024 25492
rect 18972 25449 18981 25483
rect 18981 25449 19015 25483
rect 19015 25449 19024 25483
rect 18972 25440 19024 25449
rect 20260 25440 20312 25492
rect 21272 25440 21324 25492
rect 22376 25483 22428 25492
rect 22376 25449 22385 25483
rect 22385 25449 22419 25483
rect 22419 25449 22428 25483
rect 22376 25440 22428 25449
rect 23388 25440 23440 25492
rect 5540 25372 5592 25424
rect 15660 25372 15712 25424
rect 2872 25100 2924 25152
rect 3608 25100 3660 25152
rect 4160 25100 4212 25152
rect 5080 25100 5132 25152
rect 11244 25304 11296 25356
rect 12900 25304 12952 25356
rect 12992 25347 13044 25356
rect 12992 25313 13001 25347
rect 13001 25313 13035 25347
rect 13035 25313 13044 25347
rect 12992 25304 13044 25313
rect 16580 25347 16632 25356
rect 16580 25313 16589 25347
rect 16589 25313 16623 25347
rect 16623 25313 16632 25347
rect 22192 25372 22244 25424
rect 16580 25304 16632 25313
rect 20076 25304 20128 25356
rect 11152 25236 11204 25288
rect 11060 25168 11112 25220
rect 12440 25236 12492 25288
rect 14556 25236 14608 25288
rect 16028 25236 16080 25288
rect 16304 25279 16356 25288
rect 16304 25245 16313 25279
rect 16313 25245 16347 25279
rect 16347 25245 16356 25279
rect 16304 25236 16356 25245
rect 18880 25236 18932 25288
rect 19340 25236 19392 25288
rect 12532 25168 12584 25220
rect 15200 25168 15252 25220
rect 20260 25236 20312 25288
rect 20720 25236 20772 25288
rect 21916 25279 21968 25288
rect 21916 25245 21925 25279
rect 21925 25245 21959 25279
rect 21959 25245 21968 25279
rect 23388 25304 23440 25356
rect 21916 25236 21968 25245
rect 23204 25236 23256 25288
rect 23940 25236 23992 25288
rect 24584 25279 24636 25288
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 25412 25279 25464 25288
rect 25412 25245 25421 25279
rect 25421 25245 25455 25279
rect 25455 25245 25464 25279
rect 25412 25236 25464 25245
rect 26884 25440 26936 25492
rect 32404 25440 32456 25492
rect 30932 25347 30984 25356
rect 30932 25313 30941 25347
rect 30941 25313 30975 25347
rect 30975 25313 30984 25347
rect 30932 25304 30984 25313
rect 30840 25279 30892 25288
rect 30840 25245 30849 25279
rect 30849 25245 30883 25279
rect 30883 25245 30892 25279
rect 30840 25236 30892 25245
rect 34336 25279 34388 25288
rect 34336 25245 34345 25279
rect 34345 25245 34379 25279
rect 34379 25245 34388 25279
rect 34336 25236 34388 25245
rect 5632 25100 5684 25152
rect 14372 25143 14424 25152
rect 14372 25109 14381 25143
rect 14381 25109 14415 25143
rect 14415 25109 14424 25143
rect 14372 25100 14424 25109
rect 16120 25100 16172 25152
rect 16764 25100 16816 25152
rect 17684 25100 17736 25152
rect 17960 25100 18012 25152
rect 27804 25168 27856 25220
rect 34060 25168 34112 25220
rect 32128 25100 32180 25152
rect 32404 25100 32456 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 11152 24939 11204 24948
rect 11152 24905 11161 24939
rect 11161 24905 11195 24939
rect 11195 24905 11204 24939
rect 11152 24896 11204 24905
rect 11244 24896 11296 24948
rect 12440 24896 12492 24948
rect 12532 24939 12584 24948
rect 12532 24905 12541 24939
rect 12541 24905 12575 24939
rect 12575 24905 12584 24939
rect 12532 24896 12584 24905
rect 14556 24939 14608 24948
rect 14556 24905 14565 24939
rect 14565 24905 14599 24939
rect 14599 24905 14608 24939
rect 14556 24896 14608 24905
rect 14924 24939 14976 24948
rect 14924 24905 14933 24939
rect 14933 24905 14967 24939
rect 14967 24905 14976 24939
rect 14924 24896 14976 24905
rect 15384 24939 15436 24948
rect 15384 24905 15393 24939
rect 15393 24905 15427 24939
rect 15427 24905 15436 24939
rect 15384 24896 15436 24905
rect 16580 24896 16632 24948
rect 17132 24896 17184 24948
rect 3976 24828 4028 24880
rect 940 24760 992 24812
rect 4068 24803 4120 24812
rect 4068 24769 4077 24803
rect 4077 24769 4111 24803
rect 4111 24769 4120 24803
rect 4068 24760 4120 24769
rect 4252 24803 4304 24812
rect 4252 24769 4261 24803
rect 4261 24769 4295 24803
rect 4295 24769 4304 24803
rect 4252 24760 4304 24769
rect 4620 24760 4672 24812
rect 5356 24760 5408 24812
rect 6000 24828 6052 24880
rect 9404 24828 9456 24880
rect 10692 24828 10744 24880
rect 5540 24760 5592 24812
rect 5908 24760 5960 24812
rect 7932 24760 7984 24812
rect 8300 24760 8352 24812
rect 5724 24735 5776 24744
rect 5724 24701 5733 24735
rect 5733 24701 5767 24735
rect 5767 24701 5776 24735
rect 5724 24692 5776 24701
rect 1584 24599 1636 24608
rect 1584 24565 1593 24599
rect 1593 24565 1627 24599
rect 1627 24565 1636 24599
rect 1584 24556 1636 24565
rect 3608 24556 3660 24608
rect 4712 24556 4764 24608
rect 11152 24760 11204 24812
rect 11428 24760 11480 24812
rect 11704 24803 11756 24812
rect 11704 24769 11713 24803
rect 11713 24769 11747 24803
rect 11747 24769 11756 24803
rect 11704 24760 11756 24769
rect 12164 24803 12216 24812
rect 12164 24769 12173 24803
rect 12173 24769 12207 24803
rect 12207 24769 12216 24803
rect 12164 24760 12216 24769
rect 12348 24803 12400 24812
rect 12348 24769 12357 24803
rect 12357 24769 12391 24803
rect 12391 24769 12400 24803
rect 12348 24760 12400 24769
rect 12440 24803 12492 24812
rect 12440 24769 12449 24803
rect 12449 24769 12483 24803
rect 12483 24769 12492 24803
rect 15016 24828 15068 24880
rect 12440 24760 12492 24769
rect 14188 24760 14240 24812
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 15568 24871 15620 24880
rect 15568 24837 15595 24871
rect 15595 24837 15620 24871
rect 15568 24828 15620 24837
rect 15660 24828 15712 24880
rect 16396 24760 16448 24812
rect 17224 24828 17276 24880
rect 14464 24624 14516 24676
rect 15200 24624 15252 24676
rect 10140 24599 10192 24608
rect 10140 24565 10149 24599
rect 10149 24565 10183 24599
rect 10183 24565 10192 24599
rect 10140 24556 10192 24565
rect 11980 24599 12032 24608
rect 11980 24565 11989 24599
rect 11989 24565 12023 24599
rect 12023 24565 12032 24599
rect 11980 24556 12032 24565
rect 13544 24556 13596 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 14648 24556 14700 24608
rect 16764 24692 16816 24744
rect 17040 24803 17092 24812
rect 17040 24769 17049 24803
rect 17049 24769 17083 24803
rect 17083 24769 17092 24803
rect 17040 24760 17092 24769
rect 18236 24760 18288 24812
rect 18788 24803 18840 24812
rect 18788 24769 18797 24803
rect 18797 24769 18831 24803
rect 18831 24769 18840 24803
rect 18788 24760 18840 24769
rect 23204 24939 23256 24948
rect 23204 24905 23213 24939
rect 23213 24905 23247 24939
rect 23247 24905 23256 24939
rect 23204 24896 23256 24905
rect 23940 24939 23992 24948
rect 23940 24905 23949 24939
rect 23949 24905 23983 24939
rect 23983 24905 23992 24939
rect 23940 24896 23992 24905
rect 24584 24939 24636 24948
rect 24584 24905 24593 24939
rect 24593 24905 24627 24939
rect 24627 24905 24636 24939
rect 24584 24896 24636 24905
rect 25412 24896 25464 24948
rect 30472 24939 30524 24948
rect 30472 24905 30481 24939
rect 30481 24905 30515 24939
rect 30515 24905 30524 24939
rect 30472 24896 30524 24905
rect 30932 24896 30984 24948
rect 34336 24896 34388 24948
rect 23388 24803 23440 24812
rect 16120 24667 16172 24676
rect 16120 24633 16129 24667
rect 16129 24633 16163 24667
rect 16163 24633 16172 24667
rect 16120 24624 16172 24633
rect 15476 24556 15528 24608
rect 23388 24769 23397 24803
rect 23397 24769 23431 24803
rect 23431 24769 23440 24803
rect 23388 24760 23440 24769
rect 23940 24760 23992 24812
rect 18880 24624 18932 24676
rect 19248 24624 19300 24676
rect 21548 24624 21600 24676
rect 24032 24692 24084 24744
rect 24492 24803 24544 24812
rect 24492 24769 24501 24803
rect 24501 24769 24535 24803
rect 24535 24769 24544 24803
rect 24492 24760 24544 24769
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 18328 24556 18380 24608
rect 19616 24556 19668 24608
rect 23112 24556 23164 24608
rect 23204 24556 23256 24608
rect 23940 24556 23992 24608
rect 24860 24692 24912 24744
rect 25228 24760 25280 24812
rect 26608 24760 26660 24812
rect 27344 24556 27396 24608
rect 30656 24556 30708 24608
rect 33784 24760 33836 24812
rect 31576 24692 31628 24744
rect 32680 24735 32732 24744
rect 32680 24701 32689 24735
rect 32689 24701 32723 24735
rect 32723 24701 32732 24735
rect 32680 24692 32732 24701
rect 30840 24599 30892 24608
rect 30840 24565 30849 24599
rect 30849 24565 30883 24599
rect 30883 24565 30892 24599
rect 30840 24556 30892 24565
rect 31576 24599 31628 24608
rect 31576 24565 31585 24599
rect 31585 24565 31619 24599
rect 31619 24565 31628 24599
rect 31576 24556 31628 24565
rect 31668 24556 31720 24608
rect 32404 24556 32456 24608
rect 33324 24556 33376 24608
rect 34152 24556 34204 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1400 24216 1452 24268
rect 2044 24352 2096 24404
rect 3608 24352 3660 24404
rect 4620 24352 4672 24404
rect 5356 24352 5408 24404
rect 5724 24395 5776 24404
rect 5724 24361 5733 24395
rect 5733 24361 5767 24395
rect 5767 24361 5776 24395
rect 5724 24352 5776 24361
rect 7932 24352 7984 24404
rect 9404 24352 9456 24404
rect 9588 24352 9640 24404
rect 10140 24352 10192 24404
rect 14832 24352 14884 24404
rect 15016 24352 15068 24404
rect 1860 24259 1912 24268
rect 1860 24225 1869 24259
rect 1869 24225 1903 24259
rect 1903 24225 1912 24259
rect 1860 24216 1912 24225
rect 4160 24148 4212 24200
rect 4896 24148 4948 24200
rect 5080 24148 5132 24200
rect 5632 24148 5684 24200
rect 4068 24012 4120 24064
rect 4620 24012 4672 24064
rect 5080 24012 5132 24064
rect 12164 24148 12216 24200
rect 14648 24284 14700 24336
rect 15568 24352 15620 24404
rect 16028 24352 16080 24404
rect 18236 24352 18288 24404
rect 18604 24352 18656 24404
rect 19340 24395 19392 24404
rect 19340 24361 19349 24395
rect 19349 24361 19383 24395
rect 19383 24361 19392 24395
rect 19340 24352 19392 24361
rect 19616 24352 19668 24404
rect 13912 24191 13964 24200
rect 13912 24157 13921 24191
rect 13921 24157 13955 24191
rect 13955 24157 13964 24191
rect 13912 24148 13964 24157
rect 14096 24191 14148 24200
rect 14096 24157 14106 24191
rect 14106 24157 14140 24191
rect 14140 24157 14148 24191
rect 14096 24148 14148 24157
rect 14188 24191 14240 24200
rect 14188 24157 14197 24191
rect 14197 24157 14231 24191
rect 14231 24157 14240 24191
rect 14188 24148 14240 24157
rect 14280 24148 14332 24200
rect 15660 24284 15712 24336
rect 17316 24284 17368 24336
rect 17408 24284 17460 24336
rect 27344 24352 27396 24404
rect 27804 24352 27856 24404
rect 32680 24352 32732 24404
rect 33784 24352 33836 24404
rect 20996 24327 21048 24336
rect 20996 24293 21005 24327
rect 21005 24293 21039 24327
rect 21039 24293 21048 24327
rect 20996 24284 21048 24293
rect 33140 24284 33192 24336
rect 33324 24327 33376 24336
rect 33324 24293 33333 24327
rect 33333 24293 33367 24327
rect 33367 24293 33376 24327
rect 33324 24284 33376 24293
rect 15108 24191 15160 24200
rect 15108 24157 15119 24191
rect 15119 24157 15160 24191
rect 12992 24080 13044 24132
rect 13544 24123 13596 24132
rect 13544 24089 13553 24123
rect 13553 24089 13587 24123
rect 13587 24089 13596 24123
rect 13544 24080 13596 24089
rect 15108 24148 15160 24157
rect 15568 24191 15620 24200
rect 15568 24157 15577 24191
rect 15577 24157 15611 24191
rect 15611 24157 15620 24191
rect 16028 24191 16080 24200
rect 15568 24148 15620 24157
rect 16028 24157 16037 24191
rect 16037 24157 16071 24191
rect 16071 24157 16080 24191
rect 16028 24148 16080 24157
rect 9864 24012 9916 24064
rect 11428 24012 11480 24064
rect 12532 24012 12584 24064
rect 13912 24012 13964 24064
rect 14372 24055 14424 24064
rect 14372 24021 14381 24055
rect 14381 24021 14415 24055
rect 14415 24021 14424 24055
rect 14372 24012 14424 24021
rect 14556 24055 14608 24064
rect 14556 24021 14565 24055
rect 14565 24021 14599 24055
rect 14599 24021 14608 24055
rect 14556 24012 14608 24021
rect 15108 24012 15160 24064
rect 15476 24012 15528 24064
rect 17040 24148 17092 24200
rect 17316 24148 17368 24200
rect 17868 24148 17920 24200
rect 16212 24055 16264 24064
rect 16212 24021 16221 24055
rect 16221 24021 16255 24055
rect 16255 24021 16264 24055
rect 17684 24123 17736 24132
rect 17684 24089 17693 24123
rect 17693 24089 17727 24123
rect 17727 24089 17736 24123
rect 17684 24080 17736 24089
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 19248 24191 19300 24200
rect 16212 24012 16264 24021
rect 17132 24012 17184 24064
rect 17224 24012 17276 24064
rect 19248 24157 19257 24191
rect 19257 24157 19291 24191
rect 19291 24157 19300 24191
rect 19248 24148 19300 24157
rect 19984 24148 20036 24200
rect 21088 24216 21140 24268
rect 23112 24216 23164 24268
rect 25044 24216 25096 24268
rect 27068 24216 27120 24268
rect 30104 24216 30156 24268
rect 20812 24123 20864 24132
rect 20812 24089 20821 24123
rect 20821 24089 20855 24123
rect 20855 24089 20864 24123
rect 20812 24080 20864 24089
rect 20904 24080 20956 24132
rect 30656 24148 30708 24200
rect 31668 24080 31720 24132
rect 21180 24012 21232 24064
rect 29552 24012 29604 24064
rect 31576 24012 31628 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23808 1636 23860
rect 3792 23808 3844 23860
rect 4068 23851 4120 23860
rect 4068 23817 4077 23851
rect 4077 23817 4111 23851
rect 4111 23817 4120 23851
rect 4068 23808 4120 23817
rect 4988 23808 5040 23860
rect 2780 23672 2832 23724
rect 6368 23715 6420 23724
rect 6368 23681 6377 23715
rect 6377 23681 6411 23715
rect 6411 23681 6420 23715
rect 6368 23672 6420 23681
rect 1400 23647 1452 23656
rect 1400 23613 1409 23647
rect 1409 23613 1443 23647
rect 1443 23613 1452 23647
rect 1400 23604 1452 23613
rect 11428 23808 11480 23860
rect 12716 23808 12768 23860
rect 8300 23740 8352 23792
rect 8852 23740 8904 23792
rect 12440 23740 12492 23792
rect 9036 23715 9088 23724
rect 9036 23681 9045 23715
rect 9045 23681 9079 23715
rect 9079 23681 9088 23715
rect 9036 23672 9088 23681
rect 9772 23672 9824 23724
rect 12348 23672 12400 23724
rect 12716 23715 12768 23724
rect 12716 23681 12725 23715
rect 12725 23681 12759 23715
rect 12759 23681 12768 23715
rect 12716 23672 12768 23681
rect 12900 23672 12952 23724
rect 14372 23808 14424 23860
rect 14556 23808 14608 23860
rect 15108 23808 15160 23860
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 14280 23672 14332 23724
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 14556 23672 14608 23681
rect 16396 23851 16448 23860
rect 16396 23817 16405 23851
rect 16405 23817 16439 23851
rect 16439 23817 16448 23851
rect 16396 23808 16448 23817
rect 20996 23808 21048 23860
rect 21640 23808 21692 23860
rect 4068 23536 4120 23588
rect 11704 23536 11756 23588
rect 12624 23536 12676 23588
rect 15108 23647 15160 23656
rect 15108 23613 15117 23647
rect 15117 23613 15151 23647
rect 15151 23613 15160 23647
rect 15108 23604 15160 23613
rect 15200 23647 15252 23656
rect 15200 23613 15209 23647
rect 15209 23613 15243 23647
rect 15243 23613 15252 23647
rect 15200 23604 15252 23613
rect 17132 23740 17184 23792
rect 18328 23740 18380 23792
rect 20260 23740 20312 23792
rect 18420 23715 18472 23724
rect 18420 23681 18429 23715
rect 18429 23681 18463 23715
rect 18463 23681 18472 23715
rect 18420 23672 18472 23681
rect 18604 23715 18656 23724
rect 18604 23681 18613 23715
rect 18613 23681 18647 23715
rect 18647 23681 18656 23715
rect 18604 23672 18656 23681
rect 20444 23672 20496 23724
rect 21180 23740 21232 23792
rect 15752 23604 15804 23656
rect 16764 23604 16816 23656
rect 17316 23647 17368 23656
rect 17316 23613 17325 23647
rect 17325 23613 17359 23647
rect 17359 23613 17368 23647
rect 17316 23604 17368 23613
rect 19984 23604 20036 23656
rect 20628 23604 20680 23656
rect 20812 23647 20864 23656
rect 20812 23613 20821 23647
rect 20821 23613 20855 23647
rect 20855 23613 20864 23647
rect 20812 23604 20864 23613
rect 21272 23672 21324 23724
rect 21456 23715 21508 23724
rect 21456 23681 21487 23715
rect 21487 23681 21508 23715
rect 21456 23672 21508 23681
rect 22652 23740 22704 23792
rect 21916 23672 21968 23724
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 22836 23715 22888 23724
rect 22836 23681 22845 23715
rect 22845 23681 22879 23715
rect 22879 23681 22888 23715
rect 22836 23672 22888 23681
rect 3608 23468 3660 23520
rect 5080 23468 5132 23520
rect 7012 23468 7064 23520
rect 8760 23468 8812 23520
rect 9864 23511 9916 23520
rect 9864 23477 9873 23511
rect 9873 23477 9907 23511
rect 9907 23477 9916 23511
rect 9864 23468 9916 23477
rect 10600 23468 10652 23520
rect 11244 23511 11296 23520
rect 11244 23477 11253 23511
rect 11253 23477 11287 23511
rect 11287 23477 11296 23511
rect 11244 23468 11296 23477
rect 11980 23468 12032 23520
rect 14556 23536 14608 23588
rect 15016 23536 15068 23588
rect 16856 23468 16908 23520
rect 17684 23468 17736 23520
rect 23204 23715 23256 23724
rect 23204 23681 23213 23715
rect 23213 23681 23247 23715
rect 23247 23681 23256 23715
rect 23204 23672 23256 23681
rect 23940 23808 23992 23860
rect 26884 23808 26936 23860
rect 29552 23851 29604 23860
rect 29552 23817 29561 23851
rect 29561 23817 29595 23851
rect 29595 23817 29604 23851
rect 29552 23808 29604 23817
rect 24492 23672 24544 23724
rect 26240 23672 26292 23724
rect 27712 23672 27764 23724
rect 23020 23604 23072 23656
rect 23572 23647 23624 23656
rect 23572 23613 23581 23647
rect 23581 23613 23615 23647
rect 23615 23613 23624 23647
rect 23572 23604 23624 23613
rect 26148 23604 26200 23656
rect 26700 23647 26752 23656
rect 26700 23613 26709 23647
rect 26709 23613 26743 23647
rect 26743 23613 26752 23647
rect 26700 23604 26752 23613
rect 24768 23536 24820 23588
rect 22928 23468 22980 23520
rect 23112 23468 23164 23520
rect 30104 23511 30156 23520
rect 30104 23477 30113 23511
rect 30113 23477 30147 23511
rect 30147 23477 30156 23511
rect 30104 23468 30156 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 2780 23264 2832 23316
rect 4896 23307 4948 23316
rect 4896 23273 4905 23307
rect 4905 23273 4939 23307
rect 4939 23273 4948 23307
rect 4896 23264 4948 23273
rect 6368 23264 6420 23316
rect 4344 23128 4396 23180
rect 5724 23171 5776 23180
rect 5724 23137 5733 23171
rect 5733 23137 5767 23171
rect 5767 23137 5776 23171
rect 5724 23128 5776 23137
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 9036 23264 9088 23316
rect 11980 23264 12032 23316
rect 13820 23264 13872 23316
rect 14096 23264 14148 23316
rect 15108 23264 15160 23316
rect 15660 23307 15712 23316
rect 15660 23273 15669 23307
rect 15669 23273 15703 23307
rect 15703 23273 15712 23307
rect 15660 23264 15712 23273
rect 16028 23264 16080 23316
rect 18420 23264 18472 23316
rect 20812 23264 20864 23316
rect 21088 23264 21140 23316
rect 21456 23264 21508 23316
rect 23020 23264 23072 23316
rect 23572 23264 23624 23316
rect 26240 23264 26292 23316
rect 26700 23264 26752 23316
rect 27712 23307 27764 23316
rect 27712 23273 27721 23307
rect 27721 23273 27755 23307
rect 27755 23273 27764 23307
rect 27712 23264 27764 23273
rect 28356 23264 28408 23316
rect 15476 23196 15528 23248
rect 21180 23196 21232 23248
rect 2872 23060 2924 23112
rect 4160 23103 4212 23112
rect 4160 23069 4169 23103
rect 4169 23069 4203 23103
rect 4203 23069 4212 23103
rect 4160 23060 4212 23069
rect 5632 23060 5684 23112
rect 5816 23103 5868 23112
rect 5816 23069 5825 23103
rect 5825 23069 5859 23103
rect 5859 23069 5868 23103
rect 5816 23060 5868 23069
rect 5080 22992 5132 23044
rect 5172 22992 5224 23044
rect 6368 23060 6420 23112
rect 8760 23103 8812 23112
rect 8760 23069 8769 23103
rect 8769 23069 8803 23103
rect 8803 23069 8812 23103
rect 8760 23060 8812 23069
rect 8852 23060 8904 23112
rect 15016 23128 15068 23180
rect 15568 23128 15620 23180
rect 18236 23128 18288 23180
rect 11244 23060 11296 23112
rect 12992 23060 13044 23112
rect 3424 22924 3476 22976
rect 3608 22967 3660 22976
rect 3608 22933 3617 22967
rect 3617 22933 3651 22967
rect 3651 22933 3660 22967
rect 3608 22924 3660 22933
rect 4068 22924 4120 22976
rect 5264 22924 5316 22976
rect 8392 22924 8444 22976
rect 9956 22992 10008 23044
rect 11888 22992 11940 23044
rect 12348 22992 12400 23044
rect 14372 23060 14424 23112
rect 12716 22924 12768 22976
rect 18236 23035 18288 23044
rect 18236 23001 18245 23035
rect 18245 23001 18279 23035
rect 18279 23001 18288 23035
rect 18788 23060 18840 23112
rect 20444 23103 20496 23112
rect 20444 23069 20453 23103
rect 20453 23069 20487 23103
rect 20487 23069 20496 23103
rect 20444 23060 20496 23069
rect 20628 23103 20680 23112
rect 20628 23069 20637 23103
rect 20637 23069 20671 23103
rect 20671 23069 20680 23103
rect 20628 23060 20680 23069
rect 18236 22992 18288 23001
rect 18512 22924 18564 22976
rect 19984 22967 20036 22976
rect 19984 22933 19993 22967
rect 19993 22933 20027 22967
rect 20027 22933 20036 22967
rect 20904 23060 20956 23112
rect 19984 22924 20036 22933
rect 22928 23128 22980 23180
rect 23388 23171 23440 23180
rect 23388 23137 23397 23171
rect 23397 23137 23431 23171
rect 23431 23137 23440 23171
rect 23388 23128 23440 23137
rect 22008 22992 22060 23044
rect 21364 22924 21416 22976
rect 24768 23196 24820 23248
rect 25228 23196 25280 23248
rect 23296 22992 23348 23044
rect 22652 22967 22704 22976
rect 22652 22933 22661 22967
rect 22661 22933 22695 22967
rect 22695 22933 22704 22967
rect 22652 22924 22704 22933
rect 24492 23103 24544 23112
rect 24492 23069 24501 23103
rect 24501 23069 24535 23103
rect 24535 23069 24544 23103
rect 24492 23060 24544 23069
rect 25136 23103 25188 23112
rect 25136 23069 25145 23103
rect 25145 23069 25179 23103
rect 25179 23069 25188 23103
rect 25136 23060 25188 23069
rect 24400 22992 24452 23044
rect 24584 23035 24636 23044
rect 24584 23001 24593 23035
rect 24593 23001 24627 23035
rect 24627 23001 24636 23035
rect 24584 22992 24636 23001
rect 25320 22924 25372 22976
rect 26056 23103 26108 23112
rect 26056 23069 26065 23103
rect 26065 23069 26099 23103
rect 26099 23069 26108 23103
rect 26056 23060 26108 23069
rect 26148 23060 26200 23112
rect 26884 23060 26936 23112
rect 34336 23103 34388 23112
rect 34336 23069 34345 23103
rect 34345 23069 34379 23103
rect 34379 23069 34388 23103
rect 34336 23060 34388 23069
rect 34612 22992 34664 23044
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4344 22763 4396 22772
rect 4344 22729 4353 22763
rect 4353 22729 4387 22763
rect 4387 22729 4396 22763
rect 4344 22720 4396 22729
rect 5172 22720 5224 22772
rect 5632 22720 5684 22772
rect 5724 22720 5776 22772
rect 1768 22652 1820 22704
rect 2872 22652 2924 22704
rect 4620 22584 4672 22636
rect 5264 22627 5316 22636
rect 5264 22593 5273 22627
rect 5273 22593 5307 22627
rect 5307 22593 5316 22627
rect 5264 22584 5316 22593
rect 9956 22763 10008 22772
rect 9956 22729 9965 22763
rect 9965 22729 9999 22763
rect 9999 22729 10008 22763
rect 9956 22720 10008 22729
rect 20720 22720 20772 22772
rect 21916 22720 21968 22772
rect 23296 22720 23348 22772
rect 23388 22720 23440 22772
rect 24308 22720 24360 22772
rect 8392 22627 8444 22636
rect 8392 22593 8401 22627
rect 8401 22593 8435 22627
rect 8435 22593 8444 22627
rect 8392 22584 8444 22593
rect 3976 22516 4028 22568
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 6368 22559 6420 22568
rect 6368 22525 6377 22559
rect 6377 22525 6411 22559
rect 6411 22525 6420 22559
rect 6368 22516 6420 22525
rect 11152 22584 11204 22636
rect 12532 22584 12584 22636
rect 15384 22627 15436 22636
rect 15384 22593 15393 22627
rect 15393 22593 15427 22627
rect 15427 22593 15436 22627
rect 15384 22584 15436 22593
rect 15660 22584 15712 22636
rect 16948 22627 17000 22636
rect 16948 22593 16957 22627
rect 16957 22593 16991 22627
rect 16991 22593 17000 22627
rect 16948 22584 17000 22593
rect 20444 22652 20496 22704
rect 22008 22652 22060 22704
rect 17684 22627 17736 22636
rect 17684 22593 17693 22627
rect 17693 22593 17727 22627
rect 17727 22593 17736 22627
rect 17684 22584 17736 22593
rect 17868 22584 17920 22636
rect 18052 22627 18104 22636
rect 18052 22593 18061 22627
rect 18061 22593 18095 22627
rect 18095 22593 18104 22627
rect 18052 22584 18104 22593
rect 18236 22627 18288 22636
rect 18236 22593 18245 22627
rect 18245 22593 18279 22627
rect 18279 22593 18288 22627
rect 18236 22584 18288 22593
rect 21272 22584 21324 22636
rect 24400 22652 24452 22704
rect 24952 22627 25004 22636
rect 9772 22516 9824 22568
rect 13268 22516 13320 22568
rect 4712 22448 4764 22500
rect 2320 22380 2372 22432
rect 5356 22448 5408 22500
rect 8852 22448 8904 22500
rect 13820 22448 13872 22500
rect 14464 22448 14516 22500
rect 16856 22448 16908 22500
rect 22652 22516 22704 22568
rect 23848 22559 23900 22568
rect 23848 22525 23857 22559
rect 23857 22525 23891 22559
rect 23891 22525 23900 22559
rect 23848 22516 23900 22525
rect 24952 22593 24961 22627
rect 24961 22593 24995 22627
rect 24995 22593 25004 22627
rect 24952 22584 25004 22593
rect 25320 22627 25372 22636
rect 25320 22593 25329 22627
rect 25329 22593 25363 22627
rect 25363 22593 25372 22627
rect 25320 22584 25372 22593
rect 18512 22491 18564 22500
rect 18512 22457 18521 22491
rect 18521 22457 18555 22491
rect 18555 22457 18564 22491
rect 18512 22448 18564 22457
rect 23388 22448 23440 22500
rect 25872 22516 25924 22568
rect 24308 22448 24360 22500
rect 26056 22448 26108 22500
rect 5080 22380 5132 22432
rect 5172 22380 5224 22432
rect 14924 22423 14976 22432
rect 14924 22389 14933 22423
rect 14933 22389 14967 22423
rect 14967 22389 14976 22423
rect 14924 22380 14976 22389
rect 15568 22380 15620 22432
rect 17040 22423 17092 22432
rect 17040 22389 17049 22423
rect 17049 22389 17083 22423
rect 17083 22389 17092 22423
rect 17040 22380 17092 22389
rect 22744 22423 22796 22432
rect 22744 22389 22753 22423
rect 22753 22389 22787 22423
rect 22787 22389 22796 22423
rect 22744 22380 22796 22389
rect 23940 22423 23992 22432
rect 23940 22389 23949 22423
rect 23949 22389 23983 22423
rect 23983 22389 23992 22423
rect 23940 22380 23992 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 2872 22176 2924 22228
rect 3976 22176 4028 22228
rect 4528 22176 4580 22228
rect 4712 22219 4764 22228
rect 4712 22185 4721 22219
rect 4721 22185 4755 22219
rect 4755 22185 4764 22219
rect 4712 22176 4764 22185
rect 5264 22176 5316 22228
rect 5356 22108 5408 22160
rect 940 21972 992 22024
rect 3148 22040 3200 22092
rect 3792 22040 3844 22092
rect 8852 22176 8904 22228
rect 15384 22219 15436 22228
rect 15384 22185 15393 22219
rect 15393 22185 15427 22219
rect 15427 22185 15436 22219
rect 15384 22176 15436 22185
rect 15660 22219 15712 22228
rect 15660 22185 15669 22219
rect 15669 22185 15703 22219
rect 15703 22185 15712 22219
rect 15660 22176 15712 22185
rect 16948 22176 17000 22228
rect 20720 22219 20772 22228
rect 20720 22185 20729 22219
rect 20729 22185 20763 22219
rect 20763 22185 20772 22219
rect 20720 22176 20772 22185
rect 17776 22108 17828 22160
rect 14004 21972 14056 22024
rect 14556 21972 14608 22024
rect 14924 21972 14976 22024
rect 15476 22015 15528 22024
rect 15476 21981 15485 22015
rect 15485 21981 15519 22015
rect 15519 21981 15528 22015
rect 15476 21972 15528 21981
rect 15568 22015 15620 22024
rect 15568 21981 15577 22015
rect 15577 21981 15611 22015
rect 15611 21981 15620 22015
rect 15568 21972 15620 21981
rect 15752 22015 15804 22024
rect 15752 21981 15761 22015
rect 15761 21981 15795 22015
rect 15795 21981 15804 22015
rect 15752 21972 15804 21981
rect 16212 22015 16264 22024
rect 16212 21981 16221 22015
rect 16221 21981 16255 22015
rect 16255 21981 16264 22015
rect 16212 21972 16264 21981
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 16488 22015 16540 22024
rect 16488 21981 16497 22015
rect 16497 21981 16531 22015
rect 16531 21981 16540 22015
rect 16488 21972 16540 21981
rect 17040 22040 17092 22092
rect 16856 21972 16908 22024
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 3976 21836 4028 21888
rect 4804 21836 4856 21888
rect 4988 21836 5040 21888
rect 6368 21836 6420 21888
rect 8300 21904 8352 21956
rect 17592 21947 17644 21956
rect 17592 21913 17601 21947
rect 17601 21913 17635 21947
rect 17635 21913 17644 21947
rect 17592 21904 17644 21913
rect 17868 21972 17920 22024
rect 18696 21972 18748 22024
rect 21180 22108 21232 22160
rect 21364 22176 21416 22228
rect 22560 22219 22612 22228
rect 22560 22185 22569 22219
rect 22569 22185 22603 22219
rect 22603 22185 22612 22219
rect 22560 22176 22612 22185
rect 23664 22219 23716 22228
rect 23664 22185 23673 22219
rect 23673 22185 23707 22219
rect 23707 22185 23716 22219
rect 23664 22176 23716 22185
rect 23940 22176 23992 22228
rect 21272 22040 21324 22092
rect 26148 22108 26200 22160
rect 34336 22176 34388 22228
rect 21180 21972 21232 22024
rect 21916 22015 21968 22024
rect 21916 21981 21925 22015
rect 21925 21981 21959 22015
rect 21959 21981 21968 22015
rect 21916 21972 21968 21981
rect 22192 21947 22244 21956
rect 22192 21913 22197 21947
rect 22197 21913 22231 21947
rect 22231 21913 22244 21947
rect 8392 21836 8444 21888
rect 9404 21836 9456 21888
rect 11612 21836 11664 21888
rect 13268 21836 13320 21888
rect 13636 21836 13688 21888
rect 13912 21836 13964 21888
rect 16304 21836 16356 21888
rect 16856 21836 16908 21888
rect 17224 21836 17276 21888
rect 20352 21879 20404 21888
rect 20352 21845 20361 21879
rect 20361 21845 20395 21879
rect 20395 21845 20404 21879
rect 20352 21836 20404 21845
rect 20904 21879 20956 21888
rect 20904 21845 20913 21879
rect 20913 21845 20947 21879
rect 20947 21845 20956 21879
rect 22192 21904 22244 21913
rect 20904 21836 20956 21845
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 23020 22015 23072 22024
rect 23020 21981 23029 22015
rect 23029 21981 23063 22015
rect 23063 21981 23072 22015
rect 23020 21972 23072 21981
rect 23388 22015 23440 22024
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23388 21972 23440 21981
rect 23756 21972 23808 22024
rect 31116 22083 31168 22092
rect 31116 22049 31125 22083
rect 31125 22049 31159 22083
rect 31159 22049 31168 22083
rect 31116 22040 31168 22049
rect 31668 22083 31720 22092
rect 31668 22049 31677 22083
rect 31677 22049 31711 22083
rect 31711 22049 31720 22083
rect 31668 22040 31720 22049
rect 32312 22083 32364 22092
rect 32312 22049 32321 22083
rect 32321 22049 32355 22083
rect 32355 22049 32364 22083
rect 32312 22040 32364 22049
rect 23204 21836 23256 21888
rect 32036 21947 32088 21956
rect 32036 21913 32045 21947
rect 32045 21913 32079 21947
rect 32079 21913 32088 21947
rect 32036 21904 32088 21913
rect 33324 21904 33376 21956
rect 23572 21836 23624 21888
rect 30288 21836 30340 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1584 21632 1636 21684
rect 4804 21632 4856 21684
rect 3332 21564 3384 21616
rect 2320 21539 2372 21548
rect 2320 21505 2329 21539
rect 2329 21505 2363 21539
rect 2363 21505 2372 21539
rect 2320 21496 2372 21505
rect 4436 21539 4488 21548
rect 4436 21505 4445 21539
rect 4445 21505 4479 21539
rect 4479 21505 4488 21539
rect 4436 21496 4488 21505
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 7380 21564 7432 21616
rect 5356 21539 5408 21548
rect 5356 21505 5365 21539
rect 5365 21505 5399 21539
rect 5399 21505 5408 21539
rect 5356 21496 5408 21505
rect 3976 21428 4028 21480
rect 4988 21428 5040 21480
rect 6368 21471 6420 21480
rect 6368 21437 6377 21471
rect 6377 21437 6411 21471
rect 6411 21437 6420 21471
rect 6368 21428 6420 21437
rect 9680 21496 9732 21548
rect 11152 21632 11204 21684
rect 11612 21675 11664 21684
rect 11244 21564 11296 21616
rect 11612 21641 11621 21675
rect 11621 21641 11655 21675
rect 11655 21641 11664 21675
rect 11612 21632 11664 21641
rect 11980 21675 12032 21684
rect 11980 21641 11989 21675
rect 11989 21641 12023 21675
rect 12023 21641 12032 21675
rect 11980 21632 12032 21641
rect 13268 21675 13320 21684
rect 13268 21641 13277 21675
rect 13277 21641 13311 21675
rect 13311 21641 13320 21675
rect 13268 21632 13320 21641
rect 13452 21632 13504 21684
rect 11520 21539 11572 21548
rect 11520 21505 11529 21539
rect 11529 21505 11563 21539
rect 11563 21505 11572 21539
rect 11520 21496 11572 21505
rect 10784 21428 10836 21480
rect 10968 21428 11020 21480
rect 13268 21496 13320 21548
rect 12348 21428 12400 21480
rect 13544 21496 13596 21548
rect 13912 21496 13964 21548
rect 14004 21539 14056 21548
rect 14004 21505 14013 21539
rect 14013 21505 14047 21539
rect 14047 21505 14056 21539
rect 14004 21496 14056 21505
rect 16212 21632 16264 21684
rect 16488 21632 16540 21684
rect 17224 21632 17276 21684
rect 17684 21632 17736 21684
rect 17960 21632 18012 21684
rect 18052 21632 18104 21684
rect 21180 21632 21232 21684
rect 23204 21632 23256 21684
rect 23664 21632 23716 21684
rect 4436 21292 4488 21344
rect 4896 21292 4948 21344
rect 5172 21292 5224 21344
rect 9404 21292 9456 21344
rect 10416 21335 10468 21344
rect 10416 21301 10425 21335
rect 10425 21301 10459 21335
rect 10459 21301 10468 21335
rect 10416 21292 10468 21301
rect 10508 21335 10560 21344
rect 10508 21301 10517 21335
rect 10517 21301 10551 21335
rect 10551 21301 10560 21335
rect 10508 21292 10560 21301
rect 11796 21292 11848 21344
rect 13912 21335 13964 21344
rect 13912 21301 13921 21335
rect 13921 21301 13955 21335
rect 13955 21301 13964 21335
rect 13912 21292 13964 21301
rect 14372 21292 14424 21344
rect 15016 21292 15068 21344
rect 15476 21292 15528 21344
rect 15660 21292 15712 21344
rect 17500 21539 17552 21548
rect 17500 21505 17509 21539
rect 17509 21505 17543 21539
rect 17543 21505 17552 21539
rect 17500 21496 17552 21505
rect 17776 21539 17828 21548
rect 17776 21505 17785 21539
rect 17785 21505 17819 21539
rect 17819 21505 17828 21539
rect 17776 21496 17828 21505
rect 17868 21496 17920 21548
rect 18052 21496 18104 21548
rect 22192 21564 22244 21616
rect 20444 21539 20496 21548
rect 20444 21505 20453 21539
rect 20453 21505 20487 21539
rect 20487 21505 20496 21539
rect 20444 21496 20496 21505
rect 20536 21539 20588 21548
rect 20536 21505 20545 21539
rect 20545 21505 20579 21539
rect 20579 21505 20588 21539
rect 20536 21496 20588 21505
rect 20720 21539 20772 21548
rect 20720 21505 20729 21539
rect 20729 21505 20763 21539
rect 20763 21505 20772 21539
rect 20720 21496 20772 21505
rect 20904 21496 20956 21548
rect 20996 21496 21048 21548
rect 21916 21496 21968 21548
rect 28356 21607 28408 21616
rect 28356 21573 28365 21607
rect 28365 21573 28399 21607
rect 28399 21573 28408 21607
rect 28356 21564 28408 21573
rect 30288 21675 30340 21684
rect 30288 21641 30297 21675
rect 30297 21641 30331 21675
rect 30331 21641 30340 21675
rect 30288 21632 30340 21641
rect 31116 21675 31168 21684
rect 31116 21641 31125 21675
rect 31125 21641 31159 21675
rect 31159 21641 31168 21675
rect 31116 21632 31168 21641
rect 31576 21675 31628 21684
rect 31576 21641 31585 21675
rect 31585 21641 31619 21675
rect 31619 21641 31628 21675
rect 31576 21632 31628 21641
rect 33324 21675 33376 21684
rect 33324 21641 33333 21675
rect 33333 21641 33367 21675
rect 33367 21641 33376 21675
rect 33324 21632 33376 21641
rect 23572 21539 23624 21548
rect 23572 21505 23581 21539
rect 23581 21505 23615 21539
rect 23615 21505 23624 21539
rect 23572 21496 23624 21505
rect 24952 21496 25004 21548
rect 26424 21539 26476 21548
rect 26424 21505 26433 21539
rect 26433 21505 26467 21539
rect 26467 21505 26476 21539
rect 26424 21496 26476 21505
rect 30104 21496 30156 21548
rect 31024 21496 31076 21548
rect 32036 21496 32088 21548
rect 21272 21428 21324 21480
rect 24860 21428 24912 21480
rect 17868 21360 17920 21412
rect 23756 21360 23808 21412
rect 18696 21335 18748 21344
rect 18696 21301 18705 21335
rect 18705 21301 18739 21335
rect 18739 21301 18748 21335
rect 18696 21292 18748 21301
rect 32404 21335 32456 21344
rect 32404 21301 32413 21335
rect 32413 21301 32447 21335
rect 32447 21301 32456 21335
rect 32404 21292 32456 21301
rect 32680 21292 32732 21344
rect 33140 21335 33192 21344
rect 33140 21301 33149 21335
rect 33149 21301 33183 21335
rect 33183 21301 33192 21335
rect 33140 21292 33192 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3148 21131 3200 21140
rect 3148 21097 3157 21131
rect 3157 21097 3191 21131
rect 3191 21097 3200 21131
rect 3148 21088 3200 21097
rect 3332 21131 3384 21140
rect 3332 21097 3341 21131
rect 3341 21097 3375 21131
rect 3375 21097 3384 21131
rect 3332 21088 3384 21097
rect 3240 20927 3292 20936
rect 3240 20893 3249 20927
rect 3249 20893 3283 20927
rect 3283 20893 3292 20927
rect 3240 20884 3292 20893
rect 5080 21088 5132 21140
rect 5172 21088 5224 21140
rect 5816 21088 5868 21140
rect 7380 21131 7432 21140
rect 7380 21097 7389 21131
rect 7389 21097 7423 21131
rect 7423 21097 7432 21131
rect 7380 21088 7432 21097
rect 10416 21088 10468 21140
rect 10508 21088 10560 21140
rect 15752 21088 15804 21140
rect 17224 21088 17276 21140
rect 17500 21088 17552 21140
rect 17868 21131 17920 21140
rect 17868 21097 17877 21131
rect 17877 21097 17911 21131
rect 17911 21097 17920 21131
rect 17868 21088 17920 21097
rect 23020 21131 23072 21140
rect 23020 21097 23029 21131
rect 23029 21097 23063 21131
rect 23063 21097 23072 21131
rect 23020 21088 23072 21097
rect 26424 21131 26476 21140
rect 26424 21097 26433 21131
rect 26433 21097 26467 21131
rect 26467 21097 26476 21131
rect 26424 21088 26476 21097
rect 9680 21020 9732 21072
rect 6000 20952 6052 21004
rect 10876 21020 10928 21072
rect 4988 20927 5040 20936
rect 4988 20893 4997 20927
rect 4997 20893 5031 20927
rect 5031 20893 5040 20927
rect 4988 20884 5040 20893
rect 6092 20859 6144 20868
rect 6092 20825 6101 20859
rect 6101 20825 6135 20859
rect 6135 20825 6144 20859
rect 6092 20816 6144 20825
rect 8392 20884 8444 20936
rect 10692 20927 10744 20936
rect 10692 20893 10701 20927
rect 10701 20893 10735 20927
rect 10735 20893 10744 20927
rect 10692 20884 10744 20893
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 10968 20884 11020 20936
rect 11152 20927 11204 20936
rect 11152 20893 11161 20927
rect 11161 20893 11195 20927
rect 11195 20893 11204 20927
rect 11152 20884 11204 20893
rect 11244 20927 11296 20936
rect 11244 20893 11253 20927
rect 11253 20893 11287 20927
rect 11287 20893 11296 20927
rect 11244 20884 11296 20893
rect 13912 20952 13964 21004
rect 11796 20884 11848 20936
rect 9404 20816 9456 20868
rect 4804 20748 4856 20800
rect 7564 20748 7616 20800
rect 9588 20748 9640 20800
rect 11428 20816 11480 20868
rect 14280 20884 14332 20936
rect 14372 20927 14424 20936
rect 14372 20893 14381 20927
rect 14381 20893 14415 20927
rect 14415 20893 14424 20927
rect 14372 20884 14424 20893
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 10876 20748 10928 20800
rect 10968 20791 11020 20800
rect 10968 20757 10977 20791
rect 10977 20757 11011 20791
rect 11011 20757 11020 20791
rect 10968 20748 11020 20757
rect 11704 20748 11756 20800
rect 15200 20927 15252 20936
rect 15200 20893 15209 20927
rect 15209 20893 15243 20927
rect 15243 20893 15252 20927
rect 15200 20884 15252 20893
rect 15476 20927 15528 20936
rect 15476 20893 15485 20927
rect 15485 20893 15519 20927
rect 15519 20893 15528 20927
rect 15476 20884 15528 20893
rect 15660 20927 15712 20936
rect 15660 20893 15669 20927
rect 15669 20893 15703 20927
rect 15703 20893 15712 20927
rect 15660 20884 15712 20893
rect 17316 20884 17368 20936
rect 20352 20995 20404 21004
rect 20352 20961 20361 20995
rect 20361 20961 20395 20995
rect 20395 20961 20404 20995
rect 20352 20952 20404 20961
rect 25136 20995 25188 21004
rect 25136 20961 25145 20995
rect 25145 20961 25179 20995
rect 25179 20961 25188 20995
rect 25136 20952 25188 20961
rect 17960 20884 18012 20936
rect 20720 20884 20772 20936
rect 21732 20927 21784 20936
rect 21732 20893 21741 20927
rect 21741 20893 21775 20927
rect 21775 20893 21784 20927
rect 21732 20884 21784 20893
rect 24860 20884 24912 20936
rect 25044 20884 25096 20936
rect 25504 20927 25556 20936
rect 25504 20893 25513 20927
rect 25513 20893 25547 20927
rect 25547 20893 25556 20927
rect 25504 20884 25556 20893
rect 15568 20816 15620 20868
rect 16304 20816 16356 20868
rect 25780 20927 25832 20936
rect 25780 20893 25789 20927
rect 25789 20893 25823 20927
rect 25823 20893 25832 20927
rect 25780 20884 25832 20893
rect 25872 20884 25924 20936
rect 33324 20927 33376 20936
rect 33324 20893 33333 20927
rect 33333 20893 33367 20927
rect 33367 20893 33376 20927
rect 33324 20884 33376 20893
rect 26332 20816 26384 20868
rect 34336 20859 34388 20868
rect 34336 20825 34345 20859
rect 34345 20825 34379 20859
rect 34379 20825 34388 20859
rect 34336 20816 34388 20825
rect 12900 20791 12952 20800
rect 12900 20757 12909 20791
rect 12909 20757 12943 20791
rect 12943 20757 12952 20791
rect 12900 20748 12952 20757
rect 14372 20748 14424 20800
rect 15384 20791 15436 20800
rect 15384 20757 15393 20791
rect 15393 20757 15427 20791
rect 15427 20757 15436 20791
rect 15384 20748 15436 20757
rect 15476 20748 15528 20800
rect 15752 20748 15804 20800
rect 16120 20748 16172 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 9680 20587 9732 20596
rect 9680 20553 9689 20587
rect 9689 20553 9723 20587
rect 9723 20553 9732 20587
rect 9680 20544 9732 20553
rect 10876 20544 10928 20596
rect 11060 20587 11112 20596
rect 11060 20553 11069 20587
rect 11069 20553 11103 20587
rect 11103 20553 11112 20587
rect 11060 20544 11112 20553
rect 11152 20544 11204 20596
rect 12900 20544 12952 20596
rect 13268 20544 13320 20596
rect 6000 20476 6052 20528
rect 7380 20476 7432 20528
rect 12532 20476 12584 20528
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 10416 20408 10468 20460
rect 11612 20408 11664 20460
rect 11704 20451 11756 20460
rect 11704 20417 11713 20451
rect 11713 20417 11747 20451
rect 11747 20417 11756 20451
rect 11704 20408 11756 20417
rect 10048 20383 10100 20392
rect 10048 20349 10057 20383
rect 10057 20349 10091 20383
rect 10091 20349 10100 20383
rect 10048 20340 10100 20349
rect 10692 20340 10744 20392
rect 9588 20272 9640 20324
rect 12532 20272 12584 20324
rect 12900 20408 12952 20460
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 13268 20451 13320 20460
rect 13268 20417 13277 20451
rect 13277 20417 13311 20451
rect 13311 20417 13320 20451
rect 13268 20408 13320 20417
rect 13360 20451 13412 20460
rect 13360 20417 13405 20451
rect 13405 20417 13412 20451
rect 13360 20408 13412 20417
rect 13544 20451 13596 20460
rect 13544 20417 13553 20451
rect 13553 20417 13587 20451
rect 13587 20417 13596 20451
rect 13544 20408 13596 20417
rect 13728 20408 13780 20460
rect 14280 20587 14332 20596
rect 14280 20553 14289 20587
rect 14289 20553 14323 20587
rect 14323 20553 14332 20587
rect 14280 20544 14332 20553
rect 15200 20544 15252 20596
rect 15568 20587 15620 20596
rect 15568 20553 15577 20587
rect 15577 20553 15611 20587
rect 15611 20553 15620 20587
rect 15568 20544 15620 20553
rect 14096 20451 14148 20460
rect 14096 20417 14105 20451
rect 14105 20417 14139 20451
rect 14139 20417 14148 20451
rect 14096 20408 14148 20417
rect 14280 20408 14332 20460
rect 14556 20408 14608 20460
rect 17684 20544 17736 20596
rect 20444 20544 20496 20596
rect 20904 20587 20956 20596
rect 20904 20553 20913 20587
rect 20913 20553 20947 20587
rect 20947 20553 20956 20587
rect 20904 20544 20956 20553
rect 17040 20476 17092 20528
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 13636 20272 13688 20324
rect 15476 20383 15528 20392
rect 15476 20349 15485 20383
rect 15485 20349 15519 20383
rect 15519 20349 15528 20383
rect 15476 20340 15528 20349
rect 13820 20272 13872 20324
rect 16304 20340 16356 20392
rect 15844 20204 15896 20256
rect 17040 20247 17092 20256
rect 17040 20213 17049 20247
rect 17049 20213 17083 20247
rect 17083 20213 17092 20247
rect 17040 20204 17092 20213
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17960 20383 18012 20392
rect 17960 20349 17969 20383
rect 17969 20349 18003 20383
rect 18003 20349 18012 20383
rect 17960 20340 18012 20349
rect 17316 20272 17368 20324
rect 20352 20408 20404 20460
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 21732 20476 21784 20528
rect 20352 20272 20404 20324
rect 20812 20340 20864 20392
rect 20628 20272 20680 20324
rect 21272 20408 21324 20460
rect 22652 20544 22704 20596
rect 24584 20587 24636 20596
rect 24584 20553 24593 20587
rect 24593 20553 24627 20587
rect 24627 20553 24636 20587
rect 24584 20544 24636 20553
rect 24952 20544 25004 20596
rect 33324 20544 33376 20596
rect 17776 20204 17828 20256
rect 19524 20204 19576 20256
rect 24676 20408 24728 20460
rect 25136 20451 25188 20460
rect 25136 20417 25145 20451
rect 25145 20417 25179 20451
rect 25179 20417 25188 20451
rect 25136 20408 25188 20417
rect 33232 20476 33284 20528
rect 25780 20408 25832 20460
rect 26332 20408 26384 20460
rect 24860 20272 24912 20324
rect 22468 20204 22520 20256
rect 22560 20247 22612 20256
rect 22560 20213 22569 20247
rect 22569 20213 22603 20247
rect 22603 20213 22612 20247
rect 22560 20204 22612 20213
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 23756 20204 23808 20256
rect 25596 20272 25648 20324
rect 26516 20247 26568 20256
rect 26516 20213 26525 20247
rect 26525 20213 26559 20247
rect 26559 20213 26568 20247
rect 26516 20204 26568 20213
rect 32496 20383 32548 20392
rect 32496 20349 32505 20383
rect 32505 20349 32539 20383
rect 32539 20349 32548 20383
rect 32496 20340 32548 20349
rect 32680 20204 32732 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 7380 20043 7432 20052
rect 7380 20009 7389 20043
rect 7389 20009 7423 20043
rect 7423 20009 7432 20043
rect 7380 20000 7432 20009
rect 8300 20043 8352 20052
rect 8300 20009 8309 20043
rect 8309 20009 8343 20043
rect 8343 20009 8352 20043
rect 8300 20000 8352 20009
rect 11060 20043 11112 20052
rect 11060 20009 11069 20043
rect 11069 20009 11103 20043
rect 11103 20009 11112 20043
rect 11060 20000 11112 20009
rect 13728 20000 13780 20052
rect 14096 20000 14148 20052
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 14372 20000 14424 20052
rect 15476 20000 15528 20052
rect 16304 20043 16356 20052
rect 16304 20009 16313 20043
rect 16313 20009 16347 20043
rect 16347 20009 16356 20043
rect 16304 20000 16356 20009
rect 10784 19932 10836 19984
rect 12072 19932 12124 19984
rect 13268 19932 13320 19984
rect 11060 19864 11112 19916
rect 17592 20000 17644 20052
rect 20444 20000 20496 20052
rect 21548 20000 21600 20052
rect 18512 19932 18564 19984
rect 940 19796 992 19848
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 11796 19796 11848 19805
rect 11980 19796 12032 19848
rect 17776 19864 17828 19916
rect 19524 19864 19576 19916
rect 20628 19932 20680 19984
rect 23020 20000 23072 20052
rect 25136 20000 25188 20052
rect 25872 20043 25924 20052
rect 25872 20009 25881 20043
rect 25881 20009 25915 20043
rect 25915 20009 25924 20043
rect 25872 20000 25924 20009
rect 22560 19932 22612 19984
rect 26516 20000 26568 20052
rect 22192 19864 22244 19916
rect 13452 19839 13504 19848
rect 13452 19805 13461 19839
rect 13461 19805 13495 19839
rect 13495 19805 13504 19839
rect 13452 19796 13504 19805
rect 11612 19728 11664 19780
rect 1584 19703 1636 19712
rect 1584 19669 1593 19703
rect 1593 19669 1627 19703
rect 1627 19669 1636 19703
rect 1584 19660 1636 19669
rect 7564 19660 7616 19712
rect 12624 19660 12676 19712
rect 13636 19728 13688 19780
rect 13820 19839 13872 19848
rect 13820 19805 13829 19839
rect 13829 19805 13863 19839
rect 13863 19805 13872 19839
rect 13820 19796 13872 19805
rect 15844 19796 15896 19848
rect 14372 19660 14424 19712
rect 15568 19660 15620 19712
rect 16580 19660 16632 19712
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 22376 19839 22428 19848
rect 22376 19805 22385 19839
rect 22385 19805 22419 19839
rect 22419 19805 22428 19839
rect 22376 19796 22428 19805
rect 22652 19839 22704 19848
rect 22652 19805 22661 19839
rect 22661 19805 22695 19839
rect 22695 19805 22704 19839
rect 22652 19796 22704 19805
rect 27160 19932 27212 19984
rect 24860 19864 24912 19916
rect 25780 19864 25832 19916
rect 30104 20043 30156 20052
rect 30104 20009 30113 20043
rect 30113 20009 30147 20043
rect 30147 20009 30156 20043
rect 30104 20000 30156 20009
rect 20444 19771 20496 19780
rect 20444 19737 20453 19771
rect 20453 19737 20487 19771
rect 20487 19737 20496 19771
rect 20444 19728 20496 19737
rect 17500 19660 17552 19712
rect 20352 19660 20404 19712
rect 23756 19728 23808 19780
rect 25596 19839 25648 19848
rect 25596 19805 25605 19839
rect 25605 19805 25639 19839
rect 25639 19805 25648 19839
rect 25596 19796 25648 19805
rect 25320 19771 25372 19780
rect 25320 19737 25329 19771
rect 25329 19737 25363 19771
rect 25363 19737 25372 19771
rect 25320 19728 25372 19737
rect 27160 19796 27212 19848
rect 31116 19907 31168 19916
rect 31116 19873 31125 19907
rect 31125 19873 31159 19907
rect 31159 19873 31168 19907
rect 31116 19864 31168 19873
rect 32036 20043 32088 20052
rect 32036 20009 32045 20043
rect 32045 20009 32079 20043
rect 32079 20009 32088 20043
rect 32036 20000 32088 20009
rect 32496 20000 32548 20052
rect 33232 20000 33284 20052
rect 31392 19864 31444 19916
rect 33140 19796 33192 19848
rect 25228 19660 25280 19712
rect 25596 19660 25648 19712
rect 26792 19660 26844 19712
rect 27712 19703 27764 19712
rect 27712 19669 27721 19703
rect 27721 19669 27755 19703
rect 27755 19669 27764 19703
rect 27712 19660 27764 19669
rect 29736 19660 29788 19712
rect 30196 19660 30248 19712
rect 31484 19660 31536 19712
rect 33600 19660 33652 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 9772 19456 9824 19508
rect 10048 19456 10100 19508
rect 11980 19499 12032 19508
rect 11980 19465 11989 19499
rect 11989 19465 12023 19499
rect 12023 19465 12032 19499
rect 11980 19456 12032 19465
rect 12072 19499 12124 19508
rect 12072 19465 12081 19499
rect 12081 19465 12115 19499
rect 12115 19465 12124 19499
rect 12072 19456 12124 19465
rect 12164 19456 12216 19508
rect 13360 19456 13412 19508
rect 13820 19499 13872 19508
rect 13820 19465 13829 19499
rect 13829 19465 13863 19499
rect 13863 19465 13872 19499
rect 13820 19456 13872 19465
rect 15568 19456 15620 19508
rect 16120 19456 16172 19508
rect 16580 19456 16632 19508
rect 16672 19456 16724 19508
rect 17500 19499 17552 19508
rect 17500 19465 17509 19499
rect 17509 19465 17543 19499
rect 17543 19465 17552 19499
rect 17500 19456 17552 19465
rect 17960 19499 18012 19508
rect 17960 19465 17969 19499
rect 17969 19465 18003 19499
rect 18003 19465 18012 19499
rect 17960 19456 18012 19465
rect 9864 19320 9916 19372
rect 10968 19252 11020 19304
rect 11520 19295 11572 19304
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 11612 19252 11664 19304
rect 9680 19227 9732 19236
rect 9680 19193 9689 19227
rect 9689 19193 9723 19227
rect 9723 19193 9732 19227
rect 11796 19295 11848 19304
rect 11796 19261 11805 19295
rect 11805 19261 11839 19295
rect 11839 19261 11848 19295
rect 11796 19252 11848 19261
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 12624 19363 12676 19372
rect 12624 19329 12633 19363
rect 12633 19329 12667 19363
rect 12667 19329 12676 19363
rect 12624 19320 12676 19329
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 15200 19388 15252 19440
rect 12164 19295 12216 19304
rect 12164 19261 12173 19295
rect 12173 19261 12207 19295
rect 12207 19261 12216 19295
rect 12164 19252 12216 19261
rect 12348 19252 12400 19304
rect 9680 19184 9732 19193
rect 9220 19159 9272 19168
rect 9220 19125 9229 19159
rect 9229 19125 9263 19159
rect 9263 19125 9272 19159
rect 9220 19116 9272 19125
rect 11152 19116 11204 19168
rect 12532 19227 12584 19236
rect 12532 19193 12541 19227
rect 12541 19193 12575 19227
rect 12575 19193 12584 19227
rect 12532 19184 12584 19193
rect 12624 19116 12676 19168
rect 13268 19159 13320 19168
rect 13268 19125 13277 19159
rect 13277 19125 13311 19159
rect 13311 19125 13320 19159
rect 13268 19116 13320 19125
rect 15292 19320 15344 19372
rect 15384 19252 15436 19304
rect 20352 19456 20404 19508
rect 15752 19363 15804 19372
rect 15752 19329 15761 19363
rect 15761 19329 15795 19363
rect 15795 19329 15804 19363
rect 15752 19320 15804 19329
rect 16672 19320 16724 19372
rect 15660 19295 15712 19304
rect 15660 19261 15669 19295
rect 15669 19261 15703 19295
rect 15703 19261 15712 19295
rect 15660 19252 15712 19261
rect 16580 19252 16632 19304
rect 14740 19116 14792 19168
rect 15200 19116 15252 19168
rect 15936 19116 15988 19168
rect 17960 19320 18012 19372
rect 18052 19363 18104 19372
rect 18052 19329 18061 19363
rect 18061 19329 18095 19363
rect 18095 19329 18104 19363
rect 18052 19320 18104 19329
rect 17684 19295 17736 19304
rect 17684 19261 17693 19295
rect 17693 19261 17727 19295
rect 17727 19261 17736 19295
rect 17684 19252 17736 19261
rect 17776 19295 17828 19304
rect 17776 19261 17785 19295
rect 17785 19261 17819 19295
rect 17819 19261 17828 19295
rect 17776 19252 17828 19261
rect 18144 19295 18196 19304
rect 18144 19261 18153 19295
rect 18153 19261 18187 19295
rect 18187 19261 18196 19295
rect 18144 19252 18196 19261
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 21272 19388 21324 19440
rect 18972 19252 19024 19304
rect 17316 19159 17368 19168
rect 17316 19125 17325 19159
rect 17325 19125 17359 19159
rect 17359 19125 17368 19159
rect 17316 19116 17368 19125
rect 18328 19116 18380 19168
rect 18420 19116 18472 19168
rect 20076 19320 20128 19372
rect 20444 19320 20496 19372
rect 22192 19456 22244 19508
rect 23572 19456 23624 19508
rect 25320 19456 25372 19508
rect 25504 19499 25556 19508
rect 25504 19465 25506 19499
rect 25506 19465 25540 19499
rect 25540 19465 25556 19499
rect 25504 19456 25556 19465
rect 28356 19499 28408 19508
rect 28356 19465 28365 19499
rect 28365 19465 28399 19499
rect 28399 19465 28408 19499
rect 28356 19456 28408 19465
rect 30196 19499 30248 19508
rect 30196 19465 30205 19499
rect 30205 19465 30239 19499
rect 30239 19465 30248 19499
rect 30196 19456 30248 19465
rect 31116 19499 31168 19508
rect 31116 19465 31125 19499
rect 31125 19465 31159 19499
rect 31159 19465 31168 19499
rect 31116 19456 31168 19465
rect 27712 19388 27764 19440
rect 29736 19388 29788 19440
rect 31392 19388 31444 19440
rect 25320 19363 25372 19372
rect 25320 19329 25329 19363
rect 25329 19329 25363 19363
rect 25363 19329 25372 19363
rect 25320 19320 25372 19329
rect 25596 19363 25648 19372
rect 24676 19252 24728 19304
rect 25596 19329 25605 19363
rect 25605 19329 25639 19363
rect 25639 19329 25648 19363
rect 25596 19320 25648 19329
rect 28356 19320 28408 19372
rect 31024 19295 31076 19304
rect 31024 19261 31033 19295
rect 31033 19261 31067 19295
rect 31067 19261 31076 19295
rect 31024 19252 31076 19261
rect 32220 19184 32272 19236
rect 19248 19159 19300 19168
rect 19248 19125 19257 19159
rect 19257 19125 19291 19159
rect 19291 19125 19300 19159
rect 19248 19116 19300 19125
rect 20628 19116 20680 19168
rect 22652 19116 22704 19168
rect 23204 19159 23256 19168
rect 23204 19125 23213 19159
rect 23213 19125 23247 19159
rect 23247 19125 23256 19159
rect 23204 19116 23256 19125
rect 31484 19116 31536 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 12072 18912 12124 18964
rect 12716 18912 12768 18964
rect 13268 18912 13320 18964
rect 13544 18912 13596 18964
rect 14464 18912 14516 18964
rect 15568 18912 15620 18964
rect 15660 18955 15712 18964
rect 15660 18921 15669 18955
rect 15669 18921 15703 18955
rect 15703 18921 15712 18955
rect 15660 18912 15712 18921
rect 15752 18912 15804 18964
rect 17684 18912 17736 18964
rect 18052 18912 18104 18964
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 19248 18912 19300 18964
rect 9680 18708 9732 18760
rect 11520 18776 11572 18828
rect 10324 18751 10376 18760
rect 10324 18717 10333 18751
rect 10333 18717 10367 18751
rect 10367 18717 10376 18751
rect 10324 18708 10376 18717
rect 10968 18640 11020 18692
rect 12348 18819 12400 18828
rect 12348 18785 12357 18819
rect 12357 18785 12391 18819
rect 12391 18785 12400 18819
rect 12348 18776 12400 18785
rect 16580 18844 16632 18896
rect 15292 18776 15344 18828
rect 15200 18708 15252 18760
rect 12256 18640 12308 18692
rect 14372 18640 14424 18692
rect 15108 18640 15160 18692
rect 15936 18751 15988 18760
rect 15936 18717 15945 18751
rect 15945 18717 15979 18751
rect 15979 18717 15988 18751
rect 15936 18708 15988 18717
rect 18972 18844 19024 18896
rect 17960 18776 18012 18828
rect 9864 18572 9916 18624
rect 11704 18572 11756 18624
rect 12348 18572 12400 18624
rect 13084 18572 13136 18624
rect 13452 18615 13504 18624
rect 13452 18581 13461 18615
rect 13461 18581 13495 18615
rect 13495 18581 13504 18615
rect 13452 18572 13504 18581
rect 13912 18615 13964 18624
rect 13912 18581 13921 18615
rect 13921 18581 13955 18615
rect 13955 18581 13964 18615
rect 13912 18572 13964 18581
rect 14740 18572 14792 18624
rect 15752 18572 15804 18624
rect 17040 18751 17092 18760
rect 17040 18717 17049 18751
rect 17049 18717 17083 18751
rect 17083 18717 17092 18751
rect 17040 18708 17092 18717
rect 17224 18751 17276 18760
rect 17224 18717 17233 18751
rect 17233 18717 17267 18751
rect 17267 18717 17276 18751
rect 17224 18708 17276 18717
rect 18328 18708 18380 18760
rect 19340 18776 19392 18828
rect 16580 18640 16632 18692
rect 19432 18708 19484 18760
rect 20352 18887 20404 18896
rect 20352 18853 20361 18887
rect 20361 18853 20395 18887
rect 20395 18853 20404 18887
rect 20352 18844 20404 18853
rect 25320 18912 25372 18964
rect 26792 18955 26844 18964
rect 26792 18921 26801 18955
rect 26801 18921 26835 18955
rect 26835 18921 26844 18955
rect 26792 18912 26844 18921
rect 31392 18912 31444 18964
rect 27160 18844 27212 18896
rect 17960 18572 18012 18624
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 18972 18640 19024 18692
rect 19064 18640 19116 18692
rect 20720 18708 20772 18760
rect 19432 18615 19484 18624
rect 19432 18581 19441 18615
rect 19441 18581 19475 18615
rect 19475 18581 19484 18615
rect 19432 18572 19484 18581
rect 20444 18572 20496 18624
rect 22560 18751 22612 18760
rect 22560 18717 22569 18751
rect 22569 18717 22603 18751
rect 22603 18717 22612 18751
rect 22560 18708 22612 18717
rect 22836 18708 22888 18760
rect 23664 18640 23716 18692
rect 22744 18572 22796 18624
rect 25872 18572 25924 18624
rect 27160 18640 27212 18692
rect 28724 18708 28776 18760
rect 29368 18751 29420 18760
rect 29368 18717 29377 18751
rect 29377 18717 29411 18751
rect 29411 18717 29420 18751
rect 29368 18708 29420 18717
rect 27528 18640 27580 18692
rect 27712 18572 27764 18624
rect 30288 18640 30340 18692
rect 31484 18640 31536 18692
rect 32220 18751 32272 18760
rect 32220 18717 32229 18751
rect 32229 18717 32263 18751
rect 32263 18717 32272 18751
rect 32220 18708 32272 18717
rect 34520 18751 34572 18760
rect 34520 18717 34529 18751
rect 34529 18717 34563 18751
rect 34563 18717 34572 18751
rect 34520 18708 34572 18717
rect 34612 18640 34664 18692
rect 28908 18572 28960 18624
rect 31944 18615 31996 18624
rect 31944 18581 31953 18615
rect 31953 18581 31987 18615
rect 31987 18581 31996 18615
rect 31944 18572 31996 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 6368 18368 6420 18420
rect 9680 18368 9732 18420
rect 10324 18368 10376 18420
rect 10784 18368 10836 18420
rect 11612 18368 11664 18420
rect 12440 18368 12492 18420
rect 13084 18368 13136 18420
rect 13912 18368 13964 18420
rect 14004 18368 14056 18420
rect 14372 18368 14424 18420
rect 15108 18411 15160 18420
rect 15108 18377 15117 18411
rect 15117 18377 15151 18411
rect 15151 18377 15160 18411
rect 15108 18368 15160 18377
rect 1584 18300 1636 18352
rect 3424 18275 3476 18284
rect 3424 18241 3433 18275
rect 3433 18241 3467 18275
rect 3467 18241 3476 18275
rect 3424 18232 3476 18241
rect 9220 18232 9272 18284
rect 9588 18232 9640 18284
rect 11060 18232 11112 18284
rect 1400 18207 1452 18216
rect 1400 18173 1409 18207
rect 1409 18173 1443 18207
rect 1443 18173 1452 18207
rect 1400 18164 1452 18173
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 11796 18232 11848 18284
rect 12072 18232 12124 18284
rect 12808 18300 12860 18352
rect 13452 18300 13504 18352
rect 16580 18368 16632 18420
rect 18880 18411 18932 18420
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 12256 18164 12308 18216
rect 12900 18275 12952 18284
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 15292 18343 15344 18352
rect 15292 18309 15301 18343
rect 15301 18309 15335 18343
rect 15335 18309 15344 18343
rect 15292 18300 15344 18309
rect 13268 18164 13320 18216
rect 13728 18164 13780 18216
rect 13912 18164 13964 18216
rect 14464 18164 14516 18216
rect 14740 18232 14792 18284
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 15476 18275 15528 18284
rect 15476 18241 15485 18275
rect 15485 18241 15519 18275
rect 15519 18241 15528 18275
rect 15476 18232 15528 18241
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 17960 18232 18012 18284
rect 18144 18232 18196 18284
rect 12624 18096 12676 18148
rect 14832 18096 14884 18148
rect 15108 18096 15160 18148
rect 3148 18071 3200 18080
rect 3148 18037 3157 18071
rect 3157 18037 3191 18071
rect 3191 18037 3200 18071
rect 3148 18028 3200 18037
rect 3700 18071 3752 18080
rect 3700 18037 3709 18071
rect 3709 18037 3743 18071
rect 3743 18037 3752 18071
rect 3700 18028 3752 18037
rect 9864 18028 9916 18080
rect 11152 18028 11204 18080
rect 12440 18071 12492 18080
rect 12440 18037 12449 18071
rect 12449 18037 12483 18071
rect 12483 18037 12492 18071
rect 12440 18028 12492 18037
rect 12716 18071 12768 18080
rect 12716 18037 12725 18071
rect 12725 18037 12759 18071
rect 12759 18037 12768 18071
rect 12716 18028 12768 18037
rect 13176 18071 13228 18080
rect 13176 18037 13185 18071
rect 13185 18037 13219 18071
rect 13219 18037 13228 18071
rect 13176 18028 13228 18037
rect 13820 18028 13872 18080
rect 17040 18028 17092 18080
rect 17868 18028 17920 18080
rect 18880 18377 18889 18411
rect 18889 18377 18923 18411
rect 18923 18377 18932 18411
rect 18880 18368 18932 18377
rect 18972 18368 19024 18420
rect 22744 18368 22796 18420
rect 22836 18411 22888 18420
rect 22836 18377 22845 18411
rect 22845 18377 22879 18411
rect 22879 18377 22888 18411
rect 22836 18368 22888 18377
rect 30104 18411 30156 18420
rect 30104 18377 30113 18411
rect 30113 18377 30147 18411
rect 30147 18377 30156 18411
rect 30104 18368 30156 18377
rect 30288 18411 30340 18420
rect 30288 18377 30297 18411
rect 30297 18377 30331 18411
rect 30331 18377 30340 18411
rect 30288 18368 30340 18377
rect 31944 18368 31996 18420
rect 34520 18411 34572 18420
rect 34520 18377 34529 18411
rect 34529 18377 34563 18411
rect 34563 18377 34572 18411
rect 34520 18368 34572 18377
rect 18880 18275 18932 18284
rect 18880 18241 18889 18275
rect 18889 18241 18923 18275
rect 18923 18241 18932 18275
rect 18880 18232 18932 18241
rect 20076 18300 20128 18352
rect 19064 18232 19116 18284
rect 19248 18275 19300 18284
rect 19248 18241 19257 18275
rect 19257 18241 19291 18275
rect 19291 18241 19300 18275
rect 19248 18232 19300 18241
rect 19432 18232 19484 18284
rect 18420 18096 18472 18148
rect 19064 18028 19116 18080
rect 19156 18028 19208 18080
rect 21364 18028 21416 18080
rect 23204 18275 23256 18284
rect 22560 18164 22612 18216
rect 22652 18164 22704 18216
rect 23204 18241 23213 18275
rect 23213 18241 23247 18275
rect 23247 18241 23256 18275
rect 23204 18232 23256 18241
rect 27160 18232 27212 18284
rect 27896 18232 27948 18284
rect 33784 18300 33836 18352
rect 32772 18028 32824 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4068 17867 4120 17876
rect 4068 17833 4077 17867
rect 4077 17833 4111 17867
rect 4111 17833 4120 17867
rect 4068 17824 4120 17833
rect 4712 17824 4764 17876
rect 9680 17824 9732 17876
rect 11152 17824 11204 17876
rect 12716 17824 12768 17876
rect 12900 17824 12952 17876
rect 12992 17824 13044 17876
rect 14372 17867 14424 17876
rect 14372 17833 14381 17867
rect 14381 17833 14415 17867
rect 14415 17833 14424 17867
rect 14372 17824 14424 17833
rect 15108 17824 15160 17876
rect 19432 17824 19484 17876
rect 20720 17867 20772 17876
rect 20720 17833 20729 17867
rect 20729 17833 20763 17867
rect 20763 17833 20772 17867
rect 20720 17824 20772 17833
rect 11520 17799 11572 17808
rect 11520 17765 11529 17799
rect 11529 17765 11563 17799
rect 11563 17765 11572 17799
rect 11520 17756 11572 17765
rect 12532 17756 12584 17808
rect 14740 17799 14792 17808
rect 14740 17765 14749 17799
rect 14749 17765 14783 17799
rect 14783 17765 14792 17799
rect 14740 17756 14792 17765
rect 3608 17688 3660 17740
rect 5172 17688 5224 17740
rect 940 17620 992 17672
rect 3148 17620 3200 17672
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 4620 17620 4672 17672
rect 5264 17620 5316 17672
rect 6092 17620 6144 17672
rect 12072 17731 12124 17740
rect 12072 17697 12081 17731
rect 12081 17697 12115 17731
rect 12115 17697 12124 17731
rect 12072 17688 12124 17697
rect 12440 17688 12492 17740
rect 12900 17688 12952 17740
rect 20904 17756 20956 17808
rect 11060 17620 11112 17672
rect 12348 17620 12400 17672
rect 12624 17620 12676 17672
rect 1676 17484 1728 17536
rect 3976 17484 4028 17536
rect 6460 17527 6512 17536
rect 6460 17493 6469 17527
rect 6469 17493 6503 17527
rect 6503 17493 6512 17527
rect 6460 17484 6512 17493
rect 6736 17527 6788 17536
rect 6736 17493 6745 17527
rect 6745 17493 6779 17527
rect 6779 17493 6788 17527
rect 6736 17484 6788 17493
rect 9220 17484 9272 17536
rect 9864 17484 9916 17536
rect 10876 17484 10928 17536
rect 11980 17552 12032 17604
rect 13544 17663 13596 17672
rect 13544 17629 13553 17663
rect 13553 17629 13587 17663
rect 13587 17629 13596 17663
rect 13544 17620 13596 17629
rect 13636 17663 13688 17672
rect 13636 17629 13645 17663
rect 13645 17629 13679 17663
rect 13679 17629 13688 17663
rect 13636 17620 13688 17629
rect 13820 17620 13872 17672
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 12440 17527 12492 17536
rect 12440 17493 12449 17527
rect 12449 17493 12483 17527
rect 12483 17493 12492 17527
rect 12440 17484 12492 17493
rect 13728 17484 13780 17536
rect 16120 17484 16172 17536
rect 19340 17620 19392 17672
rect 21088 17688 21140 17740
rect 20076 17595 20128 17604
rect 20076 17561 20085 17595
rect 20085 17561 20119 17595
rect 20119 17561 20128 17595
rect 20076 17552 20128 17561
rect 20904 17620 20956 17672
rect 21180 17663 21232 17672
rect 21180 17629 21189 17663
rect 21189 17629 21223 17663
rect 21223 17629 21232 17663
rect 21180 17620 21232 17629
rect 21456 17663 21508 17672
rect 21456 17629 21465 17663
rect 21465 17629 21499 17663
rect 21499 17629 21508 17663
rect 21456 17620 21508 17629
rect 23020 17799 23072 17808
rect 23020 17765 23029 17799
rect 23029 17765 23063 17799
rect 23063 17765 23072 17799
rect 23020 17756 23072 17765
rect 21272 17552 21324 17604
rect 22744 17663 22796 17672
rect 22744 17629 22753 17663
rect 22753 17629 22787 17663
rect 22787 17629 22796 17663
rect 22744 17620 22796 17629
rect 27528 17824 27580 17876
rect 27712 17867 27764 17876
rect 27712 17833 27721 17867
rect 27721 17833 27755 17867
rect 27755 17833 27764 17867
rect 27712 17824 27764 17833
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 23480 17620 23532 17672
rect 23756 17663 23808 17672
rect 23756 17629 23765 17663
rect 23765 17629 23799 17663
rect 23799 17629 23808 17663
rect 23756 17620 23808 17629
rect 20720 17484 20772 17536
rect 20812 17527 20864 17536
rect 20812 17493 20821 17527
rect 20821 17493 20855 17527
rect 20855 17493 20864 17527
rect 20812 17484 20864 17493
rect 22560 17484 22612 17536
rect 22744 17484 22796 17536
rect 23664 17552 23716 17604
rect 27528 17620 27580 17672
rect 33784 17867 33836 17876
rect 33784 17833 33793 17867
rect 33793 17833 33827 17867
rect 33827 17833 33836 17867
rect 33784 17824 33836 17833
rect 28816 17799 28868 17808
rect 28816 17765 28825 17799
rect 28825 17765 28859 17799
rect 28859 17765 28868 17799
rect 28816 17756 28868 17765
rect 28724 17688 28776 17740
rect 27436 17552 27488 17604
rect 27896 17552 27948 17604
rect 28172 17552 28224 17604
rect 23112 17484 23164 17536
rect 26976 17484 27028 17536
rect 27620 17484 27672 17536
rect 27804 17484 27856 17536
rect 28448 17527 28500 17536
rect 28448 17493 28457 17527
rect 28457 17493 28491 17527
rect 28491 17493 28500 17527
rect 28448 17484 28500 17493
rect 28540 17484 28592 17536
rect 28908 17552 28960 17604
rect 33600 17527 33652 17536
rect 33600 17493 33609 17527
rect 33609 17493 33643 17527
rect 33643 17493 33652 17527
rect 33600 17484 33652 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 3240 17280 3292 17332
rect 6460 17280 6512 17332
rect 22928 17280 22980 17332
rect 23020 17280 23072 17332
rect 23112 17280 23164 17332
rect 23296 17280 23348 17332
rect 25872 17280 25924 17332
rect 27620 17280 27672 17332
rect 27804 17323 27856 17332
rect 27804 17289 27813 17323
rect 27813 17289 27847 17323
rect 27847 17289 27856 17323
rect 27804 17280 27856 17289
rect 28448 17280 28500 17332
rect 28816 17280 28868 17332
rect 29368 17280 29420 17332
rect 31484 17323 31536 17332
rect 31484 17289 31493 17323
rect 31493 17289 31527 17323
rect 31527 17289 31536 17323
rect 31484 17280 31536 17289
rect 3608 17144 3660 17196
rect 3884 17187 3936 17196
rect 3884 17153 3893 17187
rect 3893 17153 3927 17187
rect 3927 17153 3936 17187
rect 3884 17144 3936 17153
rect 6368 17144 6420 17196
rect 7564 17212 7616 17264
rect 10876 17255 10928 17264
rect 10876 17221 10885 17255
rect 10885 17221 10919 17255
rect 10919 17221 10928 17255
rect 10876 17212 10928 17221
rect 9220 17187 9272 17196
rect 3792 17119 3844 17128
rect 3792 17085 3801 17119
rect 3801 17085 3835 17119
rect 3835 17085 3844 17119
rect 3792 17076 3844 17085
rect 5080 17119 5132 17128
rect 5080 17085 5089 17119
rect 5089 17085 5123 17119
rect 5123 17085 5132 17119
rect 5080 17076 5132 17085
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 6828 17076 6880 17128
rect 7564 17076 7616 17128
rect 8760 17076 8812 17128
rect 11520 17144 11572 17196
rect 11980 17008 12032 17060
rect 12348 17144 12400 17196
rect 13268 17255 13320 17264
rect 13268 17221 13277 17255
rect 13277 17221 13311 17255
rect 13311 17221 13320 17255
rect 13268 17212 13320 17221
rect 13544 17255 13596 17264
rect 13544 17221 13553 17255
rect 13553 17221 13587 17255
rect 13587 17221 13596 17255
rect 13544 17212 13596 17221
rect 16580 17212 16632 17264
rect 18328 17255 18380 17264
rect 18328 17221 18337 17255
rect 18337 17221 18371 17255
rect 18371 17221 18380 17255
rect 18328 17212 18380 17221
rect 20812 17212 20864 17264
rect 21088 17255 21140 17264
rect 21088 17221 21097 17255
rect 21097 17221 21131 17255
rect 21131 17221 21140 17255
rect 21088 17212 21140 17221
rect 21272 17255 21324 17264
rect 21272 17221 21281 17255
rect 21281 17221 21315 17255
rect 21315 17221 21324 17255
rect 21272 17212 21324 17221
rect 21456 17255 21508 17264
rect 21456 17221 21465 17255
rect 21465 17221 21499 17255
rect 21499 17221 21508 17255
rect 21456 17212 21508 17221
rect 12440 17076 12492 17128
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 12992 17187 13044 17196
rect 12992 17153 13001 17187
rect 13001 17153 13035 17187
rect 13035 17153 13044 17187
rect 12992 17144 13044 17153
rect 15936 17144 15988 17196
rect 13912 17076 13964 17128
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 17960 17144 18012 17196
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 17408 17008 17460 17060
rect 20076 17144 20128 17196
rect 21180 17076 21232 17128
rect 22560 17076 22612 17128
rect 25228 17187 25280 17196
rect 25228 17153 25237 17187
rect 25237 17153 25271 17187
rect 25271 17153 25280 17187
rect 25228 17144 25280 17153
rect 25412 17144 25464 17196
rect 25044 17119 25096 17128
rect 25044 17085 25053 17119
rect 25053 17085 25087 17119
rect 25087 17085 25096 17119
rect 25044 17076 25096 17085
rect 25136 17119 25188 17128
rect 25136 17085 25145 17119
rect 25145 17085 25179 17119
rect 25179 17085 25188 17119
rect 25136 17076 25188 17085
rect 25872 17119 25924 17128
rect 25872 17085 25881 17119
rect 25881 17085 25915 17119
rect 25915 17085 25924 17119
rect 25872 17076 25924 17085
rect 6460 16940 6512 16992
rect 7012 16983 7064 16992
rect 7012 16949 7021 16983
rect 7021 16949 7055 16983
rect 7055 16949 7064 16983
rect 7012 16940 7064 16949
rect 9588 16940 9640 16992
rect 11704 16983 11756 16992
rect 11704 16949 11713 16983
rect 11713 16949 11747 16983
rect 11747 16949 11756 16983
rect 11704 16940 11756 16949
rect 16396 16983 16448 16992
rect 16396 16949 16405 16983
rect 16405 16949 16439 16983
rect 16439 16949 16448 16983
rect 16396 16940 16448 16949
rect 20444 17008 20496 17060
rect 20996 16940 21048 16992
rect 25596 16983 25648 16992
rect 25596 16949 25605 16983
rect 25605 16949 25639 16983
rect 25639 16949 25648 16983
rect 25596 16940 25648 16949
rect 25964 16940 26016 16992
rect 27528 17144 27580 17196
rect 27436 17076 27488 17128
rect 27804 17144 27856 17196
rect 30380 17212 30432 17264
rect 31760 17144 31812 17196
rect 31944 17144 31996 17196
rect 26240 16940 26292 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3240 16736 3292 16788
rect 3792 16779 3844 16788
rect 3792 16745 3801 16779
rect 3801 16745 3835 16779
rect 3835 16745 3844 16779
rect 3792 16736 3844 16745
rect 1676 16643 1728 16652
rect 1676 16609 1685 16643
rect 1685 16609 1719 16643
rect 1719 16609 1728 16643
rect 1676 16600 1728 16609
rect 1400 16575 1452 16584
rect 1400 16541 1409 16575
rect 1409 16541 1443 16575
rect 1443 16541 1452 16575
rect 1400 16532 1452 16541
rect 3976 16668 4028 16720
rect 4068 16643 4120 16652
rect 4068 16609 4077 16643
rect 4077 16609 4111 16643
rect 4111 16609 4120 16643
rect 4620 16668 4672 16720
rect 4068 16600 4120 16609
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 5080 16736 5132 16788
rect 5540 16668 5592 16720
rect 6828 16736 6880 16788
rect 8668 16779 8720 16788
rect 8668 16745 8677 16779
rect 8677 16745 8711 16779
rect 8711 16745 8720 16779
rect 8668 16736 8720 16745
rect 9864 16736 9916 16788
rect 12072 16736 12124 16788
rect 12992 16736 13044 16788
rect 15752 16736 15804 16788
rect 17408 16736 17460 16788
rect 18236 16736 18288 16788
rect 19984 16736 20036 16788
rect 20444 16779 20496 16788
rect 20444 16745 20453 16779
rect 20453 16745 20487 16779
rect 20487 16745 20496 16779
rect 20444 16736 20496 16745
rect 22376 16736 22428 16788
rect 22928 16736 22980 16788
rect 23572 16779 23624 16788
rect 23572 16745 23581 16779
rect 23581 16745 23615 16779
rect 23615 16745 23624 16779
rect 23572 16736 23624 16745
rect 25228 16736 25280 16788
rect 26240 16779 26292 16788
rect 26240 16745 26249 16779
rect 26249 16745 26283 16779
rect 26283 16745 26292 16779
rect 26240 16736 26292 16745
rect 30104 16736 30156 16788
rect 30380 16779 30432 16788
rect 30380 16745 30389 16779
rect 30389 16745 30423 16779
rect 30423 16745 30432 16779
rect 30380 16736 30432 16745
rect 4988 16532 5040 16584
rect 6460 16643 6512 16652
rect 6460 16609 6469 16643
rect 6469 16609 6503 16643
rect 6503 16609 6512 16643
rect 6460 16600 6512 16609
rect 9404 16600 9456 16652
rect 14188 16575 14240 16584
rect 14188 16541 14197 16575
rect 14197 16541 14231 16575
rect 14231 16541 14240 16575
rect 14188 16532 14240 16541
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 15936 16575 15988 16584
rect 15936 16541 15945 16575
rect 15945 16541 15979 16575
rect 15979 16541 15988 16575
rect 15936 16532 15988 16541
rect 16120 16575 16172 16584
rect 16120 16541 16129 16575
rect 16129 16541 16163 16575
rect 16163 16541 16172 16575
rect 16120 16532 16172 16541
rect 16396 16532 16448 16584
rect 16672 16575 16724 16584
rect 16672 16541 16681 16575
rect 16681 16541 16715 16575
rect 16715 16541 16724 16575
rect 16672 16532 16724 16541
rect 16856 16575 16908 16584
rect 16856 16541 16865 16575
rect 16865 16541 16899 16575
rect 16899 16541 16908 16575
rect 16856 16532 16908 16541
rect 19064 16600 19116 16652
rect 18328 16532 18380 16584
rect 18788 16532 18840 16584
rect 3148 16439 3200 16448
rect 3148 16405 3157 16439
rect 3157 16405 3191 16439
rect 3191 16405 3200 16439
rect 3148 16396 3200 16405
rect 4068 16396 4120 16448
rect 5264 16464 5316 16516
rect 7012 16464 7064 16516
rect 6736 16396 6788 16448
rect 10968 16396 11020 16448
rect 13360 16396 13412 16448
rect 18512 16439 18564 16448
rect 18512 16405 18521 16439
rect 18521 16405 18555 16439
rect 18555 16405 18564 16439
rect 18512 16396 18564 16405
rect 18696 16439 18748 16448
rect 18696 16405 18705 16439
rect 18705 16405 18739 16439
rect 18739 16405 18748 16439
rect 18696 16396 18748 16405
rect 22652 16668 22704 16720
rect 20812 16575 20864 16584
rect 20812 16541 20821 16575
rect 20821 16541 20855 16575
rect 20855 16541 20864 16575
rect 20812 16532 20864 16541
rect 23572 16600 23624 16652
rect 23664 16600 23716 16652
rect 23756 16532 23808 16584
rect 25412 16600 25464 16652
rect 25596 16600 25648 16652
rect 24768 16532 24820 16584
rect 24952 16532 25004 16584
rect 25872 16575 25924 16584
rect 25872 16541 25881 16575
rect 25881 16541 25915 16575
rect 25915 16541 25924 16575
rect 25872 16532 25924 16541
rect 26148 16532 26200 16584
rect 30656 16668 30708 16720
rect 32220 16736 32272 16788
rect 32680 16736 32732 16788
rect 33140 16668 33192 16720
rect 31392 16464 31444 16516
rect 32680 16600 32732 16652
rect 31760 16532 31812 16584
rect 34520 16575 34572 16584
rect 34520 16541 34529 16575
rect 34529 16541 34563 16575
rect 34563 16541 34572 16575
rect 34520 16532 34572 16541
rect 34612 16464 34664 16516
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 31944 16396 31996 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 3608 16192 3660 16244
rect 4160 16192 4212 16244
rect 10968 16235 11020 16244
rect 10968 16201 10977 16235
rect 10977 16201 11011 16235
rect 11011 16201 11020 16235
rect 10968 16192 11020 16201
rect 13912 16192 13964 16244
rect 14188 16192 14240 16244
rect 14372 16192 14424 16244
rect 16028 16192 16080 16244
rect 1400 15852 1452 15904
rect 3792 16124 3844 16176
rect 5540 16124 5592 16176
rect 11428 16124 11480 16176
rect 11520 16124 11572 16176
rect 6368 16099 6420 16108
rect 6368 16065 6377 16099
rect 6377 16065 6411 16099
rect 6411 16065 6420 16099
rect 6368 16056 6420 16065
rect 11060 16099 11112 16108
rect 11060 16065 11069 16099
rect 11069 16065 11103 16099
rect 11103 16065 11112 16099
rect 11060 16056 11112 16065
rect 11244 16056 11296 16108
rect 11888 16124 11940 16176
rect 12532 16167 12584 16176
rect 12532 16133 12541 16167
rect 12541 16133 12575 16167
rect 12575 16133 12584 16167
rect 12532 16124 12584 16133
rect 13360 16167 13412 16176
rect 13360 16133 13369 16167
rect 13369 16133 13403 16167
rect 13403 16133 13412 16167
rect 18696 16192 18748 16244
rect 13360 16124 13412 16133
rect 12440 16099 12492 16108
rect 12440 16065 12449 16099
rect 12449 16065 12483 16099
rect 12483 16065 12492 16099
rect 12440 16056 12492 16065
rect 12716 16099 12768 16108
rect 12716 16065 12725 16099
rect 12725 16065 12759 16099
rect 12759 16065 12768 16099
rect 12716 16056 12768 16065
rect 14096 16099 14148 16108
rect 14096 16065 14105 16099
rect 14105 16065 14139 16099
rect 14139 16065 14148 16099
rect 14096 16056 14148 16065
rect 14188 16056 14240 16108
rect 14280 16099 14332 16108
rect 14280 16065 14289 16099
rect 14289 16065 14323 16099
rect 14323 16065 14332 16099
rect 14280 16056 14332 16065
rect 16028 16056 16080 16108
rect 18880 16124 18932 16176
rect 15384 15988 15436 16040
rect 4068 15852 4120 15904
rect 6920 15852 6972 15904
rect 11796 15852 11848 15904
rect 11980 15895 12032 15904
rect 11980 15861 11989 15895
rect 11989 15861 12023 15895
rect 12023 15861 12032 15895
rect 11980 15852 12032 15861
rect 12164 15852 12216 15904
rect 12716 15852 12768 15904
rect 16764 15920 16816 15972
rect 17224 15920 17276 15972
rect 15660 15895 15712 15904
rect 15660 15861 15669 15895
rect 15669 15861 15703 15895
rect 15703 15861 15712 15895
rect 15660 15852 15712 15861
rect 17776 15852 17828 15904
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 19340 15988 19392 16040
rect 25136 16192 25188 16244
rect 27804 16235 27856 16244
rect 27804 16201 27813 16235
rect 27813 16201 27847 16235
rect 27847 16201 27856 16235
rect 27804 16192 27856 16201
rect 34520 16192 34572 16244
rect 22376 16056 22428 16108
rect 22560 16031 22612 16040
rect 22560 15997 22569 16031
rect 22569 15997 22603 16031
rect 22603 15997 22612 16031
rect 22560 15988 22612 15997
rect 22928 16099 22980 16108
rect 22928 16065 22937 16099
rect 22937 16065 22971 16099
rect 22971 16065 22980 16099
rect 22928 16056 22980 16065
rect 23112 16099 23164 16108
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 24124 16056 24176 16108
rect 24768 16099 24820 16108
rect 24768 16065 24777 16099
rect 24777 16065 24811 16099
rect 24811 16065 24820 16099
rect 24768 16056 24820 16065
rect 25964 16056 26016 16108
rect 27068 16056 27120 16108
rect 27160 16056 27212 16108
rect 27528 16056 27580 16108
rect 33140 16124 33192 16176
rect 33968 16124 34020 16176
rect 17960 15920 18012 15972
rect 21456 15920 21508 15972
rect 22652 15920 22704 15972
rect 18420 15852 18472 15904
rect 18788 15852 18840 15904
rect 20352 15852 20404 15904
rect 23940 15852 23992 15904
rect 25412 15852 25464 15904
rect 28356 15895 28408 15904
rect 28356 15861 28365 15895
rect 28365 15861 28399 15895
rect 28399 15861 28408 15895
rect 28356 15852 28408 15861
rect 32772 15895 32824 15904
rect 32772 15861 32781 15895
rect 32781 15861 32815 15895
rect 32815 15861 32824 15895
rect 32772 15852 32824 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3608 15691 3660 15700
rect 3608 15657 3617 15691
rect 3617 15657 3651 15691
rect 3651 15657 3660 15691
rect 3608 15648 3660 15657
rect 4620 15648 4672 15700
rect 8668 15648 8720 15700
rect 12440 15648 12492 15700
rect 1400 15580 1452 15632
rect 11060 15580 11112 15632
rect 15660 15648 15712 15700
rect 15936 15691 15988 15700
rect 15936 15657 15945 15691
rect 15945 15657 15979 15691
rect 15979 15657 15988 15691
rect 15936 15648 15988 15657
rect 18144 15648 18196 15700
rect 21456 15648 21508 15700
rect 3700 15512 3752 15564
rect 3884 15512 3936 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 11980 15512 12032 15564
rect 4068 15376 4120 15428
rect 4988 15444 5040 15496
rect 3608 15308 3660 15360
rect 3976 15308 4028 15360
rect 4804 15308 4856 15360
rect 4988 15351 5040 15360
rect 4988 15317 4997 15351
rect 4997 15317 5031 15351
rect 5031 15317 5040 15351
rect 4988 15308 5040 15317
rect 7472 15308 7524 15360
rect 8300 15308 8352 15360
rect 12532 15444 12584 15496
rect 8760 15308 8812 15360
rect 11244 15308 11296 15360
rect 11428 15308 11480 15360
rect 11520 15308 11572 15360
rect 12164 15308 12216 15360
rect 16948 15512 17000 15564
rect 14188 15487 14240 15496
rect 14188 15453 14197 15487
rect 14197 15453 14231 15487
rect 14231 15453 14240 15487
rect 14188 15444 14240 15453
rect 14372 15487 14424 15496
rect 14372 15453 14381 15487
rect 14381 15453 14415 15487
rect 14415 15453 14424 15487
rect 14372 15444 14424 15453
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 15752 15444 15804 15496
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 17040 15444 17092 15496
rect 17132 15487 17184 15496
rect 17132 15453 17141 15487
rect 17141 15453 17175 15487
rect 17175 15453 17184 15487
rect 17132 15444 17184 15453
rect 17224 15487 17276 15496
rect 17224 15453 17233 15487
rect 17233 15453 17267 15487
rect 17267 15453 17276 15487
rect 20260 15580 20312 15632
rect 20444 15623 20496 15632
rect 20444 15589 20453 15623
rect 20453 15589 20487 15623
rect 20487 15589 20496 15623
rect 22928 15648 22980 15700
rect 26976 15648 27028 15700
rect 20444 15580 20496 15589
rect 20076 15512 20128 15564
rect 17776 15487 17828 15496
rect 17224 15444 17276 15453
rect 17776 15453 17785 15487
rect 17785 15453 17819 15487
rect 17819 15453 17828 15487
rect 17776 15444 17828 15453
rect 18144 15487 18196 15496
rect 18144 15453 18153 15487
rect 18153 15453 18187 15487
rect 18187 15453 18196 15487
rect 18144 15444 18196 15453
rect 18512 15444 18564 15496
rect 20352 15487 20404 15496
rect 20352 15453 20361 15487
rect 20361 15453 20395 15487
rect 20395 15453 20404 15487
rect 20352 15444 20404 15453
rect 22284 15580 22336 15632
rect 33968 15691 34020 15700
rect 33968 15657 33977 15691
rect 33977 15657 34011 15691
rect 34011 15657 34020 15691
rect 33968 15648 34020 15657
rect 20996 15555 21048 15564
rect 20996 15521 21005 15555
rect 21005 15521 21039 15555
rect 21039 15521 21048 15555
rect 20996 15512 21048 15521
rect 12992 15308 13044 15360
rect 14280 15308 14332 15360
rect 15752 15308 15804 15360
rect 22376 15376 22428 15428
rect 16488 15308 16540 15360
rect 19064 15308 19116 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 22560 15308 22612 15360
rect 23664 15487 23716 15496
rect 23664 15453 23673 15487
rect 23673 15453 23707 15487
rect 23707 15453 23716 15487
rect 23664 15444 23716 15453
rect 23756 15487 23808 15496
rect 23756 15453 23771 15487
rect 23771 15453 23805 15487
rect 23805 15453 23808 15487
rect 23756 15444 23808 15453
rect 23940 15487 23992 15496
rect 23940 15453 23949 15487
rect 23949 15453 23983 15487
rect 23983 15453 23992 15487
rect 23940 15444 23992 15453
rect 23296 15376 23348 15428
rect 27160 15444 27212 15496
rect 28080 15555 28132 15564
rect 28080 15521 28089 15555
rect 28089 15521 28123 15555
rect 28123 15521 28132 15555
rect 28080 15512 28132 15521
rect 27896 15487 27948 15496
rect 27896 15453 27905 15487
rect 27905 15453 27939 15487
rect 27939 15453 27948 15487
rect 27896 15444 27948 15453
rect 28356 15512 28408 15564
rect 25596 15376 25648 15428
rect 26056 15351 26108 15360
rect 26056 15317 26065 15351
rect 26065 15317 26099 15351
rect 26099 15317 26108 15351
rect 26056 15308 26108 15317
rect 26240 15308 26292 15360
rect 27068 15351 27120 15360
rect 27068 15317 27077 15351
rect 27077 15317 27111 15351
rect 27111 15317 27120 15351
rect 27068 15308 27120 15317
rect 27252 15419 27304 15428
rect 27252 15385 27261 15419
rect 27261 15385 27295 15419
rect 27295 15385 27304 15419
rect 27252 15376 27304 15385
rect 27528 15376 27580 15428
rect 28356 15376 28408 15428
rect 28724 15376 28776 15428
rect 33600 15444 33652 15496
rect 27988 15308 28040 15360
rect 30196 15351 30248 15360
rect 30196 15317 30205 15351
rect 30205 15317 30239 15351
rect 30239 15317 30248 15351
rect 30196 15308 30248 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1492 15104 1544 15156
rect 3792 15147 3844 15156
rect 3792 15113 3801 15147
rect 3801 15113 3835 15147
rect 3835 15113 3844 15147
rect 3792 15104 3844 15113
rect 4804 15104 4856 15156
rect 6368 15104 6420 15156
rect 14372 15104 14424 15156
rect 15292 15104 15344 15156
rect 15384 15104 15436 15156
rect 1584 15036 1636 15088
rect 2320 15036 2372 15088
rect 5264 14968 5316 15020
rect 6920 15036 6972 15088
rect 8300 15036 8352 15088
rect 9864 15079 9916 15088
rect 9864 15045 9873 15079
rect 9873 15045 9907 15079
rect 9907 15045 9916 15079
rect 9864 15036 9916 15045
rect 8668 14968 8720 15020
rect 4988 14900 5040 14952
rect 8300 14900 8352 14952
rect 11244 14943 11296 14952
rect 11244 14909 11253 14943
rect 11253 14909 11287 14943
rect 11287 14909 11296 14943
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 12992 15036 13044 15088
rect 11796 14968 11848 14977
rect 12348 14968 12400 15020
rect 15108 15036 15160 15088
rect 16028 15104 16080 15156
rect 16672 15104 16724 15156
rect 20352 15104 20404 15156
rect 20812 15104 20864 15156
rect 21824 15104 21876 15156
rect 23756 15147 23808 15156
rect 23756 15113 23765 15147
rect 23765 15113 23799 15147
rect 23799 15113 23808 15147
rect 23756 15104 23808 15113
rect 26148 15104 26200 15156
rect 28080 15104 28132 15156
rect 28356 15147 28408 15156
rect 28356 15113 28365 15147
rect 28365 15113 28399 15147
rect 28399 15113 28408 15147
rect 28356 15104 28408 15113
rect 28724 15147 28776 15156
rect 28724 15113 28733 15147
rect 28733 15113 28767 15147
rect 28767 15113 28776 15147
rect 28724 15104 28776 15113
rect 29368 15104 29420 15156
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 15200 15011 15252 15020
rect 15200 14977 15209 15011
rect 15209 14977 15243 15011
rect 15243 14977 15252 15011
rect 15200 14968 15252 14977
rect 17040 15036 17092 15088
rect 18144 15079 18196 15088
rect 11244 14900 11296 14909
rect 14832 14900 14884 14952
rect 17132 15011 17184 15020
rect 17132 14977 17141 15011
rect 17141 14977 17175 15011
rect 17175 14977 17184 15011
rect 17132 14968 17184 14977
rect 18144 15045 18153 15079
rect 18153 15045 18187 15079
rect 18187 15045 18196 15079
rect 18144 15036 18196 15045
rect 18696 15036 18748 15088
rect 17040 14943 17092 14952
rect 17040 14909 17049 14943
rect 17049 14909 17083 14943
rect 17083 14909 17092 14943
rect 17040 14900 17092 14909
rect 17500 14943 17552 14952
rect 17500 14909 17509 14943
rect 17509 14909 17543 14943
rect 17543 14909 17552 14943
rect 17500 14900 17552 14909
rect 17684 14943 17736 14952
rect 17684 14909 17693 14943
rect 17693 14909 17727 14943
rect 17727 14909 17736 14943
rect 17684 14900 17736 14909
rect 17316 14832 17368 14884
rect 3332 14764 3384 14816
rect 3884 14764 3936 14816
rect 5172 14807 5224 14816
rect 5172 14773 5181 14807
rect 5181 14773 5215 14807
rect 5215 14773 5224 14807
rect 5172 14764 5224 14773
rect 11612 14807 11664 14816
rect 11612 14773 11621 14807
rect 11621 14773 11655 14807
rect 11655 14773 11664 14807
rect 11612 14764 11664 14773
rect 12532 14764 12584 14816
rect 15752 14764 15804 14816
rect 16212 14807 16264 14816
rect 16212 14773 16221 14807
rect 16221 14773 16255 14807
rect 16255 14773 16264 14807
rect 16212 14764 16264 14773
rect 18420 14968 18472 15020
rect 19432 15036 19484 15088
rect 20076 15036 20128 15088
rect 20260 15036 20312 15088
rect 21456 15036 21508 15088
rect 19248 14968 19300 15020
rect 20536 14968 20588 15020
rect 21364 14968 21416 15020
rect 22192 15036 22244 15088
rect 25136 15036 25188 15088
rect 23296 15011 23348 15020
rect 23296 14977 23305 15011
rect 23305 14977 23339 15011
rect 23339 14977 23348 15011
rect 23296 14968 23348 14977
rect 24032 14968 24084 15020
rect 25044 14968 25096 15020
rect 18144 14832 18196 14884
rect 19616 14900 19668 14952
rect 19340 14832 19392 14884
rect 25504 15011 25556 15020
rect 25504 14977 25513 15011
rect 25513 14977 25547 15011
rect 25547 14977 25556 15011
rect 25504 14968 25556 14977
rect 26056 15011 26108 15020
rect 26056 14977 26065 15011
rect 26065 14977 26099 15011
rect 26099 14977 26108 15011
rect 26056 14968 26108 14977
rect 26332 15011 26384 15020
rect 26332 14977 26341 15011
rect 26341 14977 26375 15011
rect 26375 14977 26384 15011
rect 26332 14968 26384 14977
rect 25412 14832 25464 14884
rect 25596 14832 25648 14884
rect 26148 14900 26200 14952
rect 27068 14968 27120 15020
rect 26240 14832 26292 14884
rect 27160 14900 27212 14952
rect 27988 14968 28040 15020
rect 28540 15011 28592 15020
rect 28540 14977 28549 15011
rect 28549 14977 28583 15011
rect 28583 14977 28592 15011
rect 28540 14968 28592 14977
rect 30196 15036 30248 15088
rect 30932 15036 30984 15088
rect 32772 14900 32824 14952
rect 19432 14764 19484 14816
rect 20076 14807 20128 14816
rect 20076 14773 20085 14807
rect 20085 14773 20119 14807
rect 20119 14773 20128 14807
rect 20076 14764 20128 14773
rect 25688 14764 25740 14816
rect 26332 14764 26384 14816
rect 31760 14807 31812 14816
rect 31760 14773 31769 14807
rect 31769 14773 31803 14807
rect 31803 14773 31812 14807
rect 31760 14764 31812 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3240 14560 3292 14612
rect 3608 14603 3660 14612
rect 3608 14569 3617 14603
rect 3617 14569 3651 14603
rect 3651 14569 3660 14603
rect 3608 14560 3660 14569
rect 3792 14560 3844 14612
rect 1492 14424 1544 14476
rect 2872 14424 2924 14476
rect 5172 14560 5224 14612
rect 8300 14603 8352 14612
rect 8300 14569 8309 14603
rect 8309 14569 8343 14603
rect 8343 14569 8352 14603
rect 8300 14560 8352 14569
rect 10968 14560 11020 14612
rect 11612 14560 11664 14612
rect 15936 14560 15988 14612
rect 16212 14560 16264 14612
rect 9588 14424 9640 14476
rect 6184 14399 6236 14408
rect 6184 14365 6193 14399
rect 6193 14365 6227 14399
rect 6227 14365 6236 14399
rect 6184 14356 6236 14365
rect 7472 14356 7524 14408
rect 1492 14288 1544 14340
rect 11060 14356 11112 14408
rect 17224 14560 17276 14612
rect 17592 14560 17644 14612
rect 18144 14603 18196 14612
rect 18144 14569 18153 14603
rect 18153 14569 18187 14603
rect 18187 14569 18196 14603
rect 18144 14560 18196 14569
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 20444 14560 20496 14612
rect 20996 14603 21048 14612
rect 20996 14569 21005 14603
rect 21005 14569 21039 14603
rect 21039 14569 21048 14603
rect 20996 14560 21048 14569
rect 25044 14560 25096 14612
rect 25412 14603 25464 14612
rect 25412 14569 25421 14603
rect 25421 14569 25455 14603
rect 25455 14569 25464 14603
rect 25412 14560 25464 14569
rect 30656 14603 30708 14612
rect 30656 14569 30665 14603
rect 30665 14569 30699 14603
rect 30699 14569 30708 14603
rect 30656 14560 30708 14569
rect 30932 14603 30984 14612
rect 30932 14569 30941 14603
rect 30941 14569 30975 14603
rect 30975 14569 30984 14603
rect 30932 14560 30984 14569
rect 11888 14288 11940 14340
rect 14372 14424 14424 14476
rect 15200 14424 15252 14476
rect 16764 14492 16816 14544
rect 21456 14535 21508 14544
rect 21456 14501 21465 14535
rect 21465 14501 21499 14535
rect 21499 14501 21508 14535
rect 21456 14492 21508 14501
rect 25688 14492 25740 14544
rect 17500 14424 17552 14476
rect 18696 14424 18748 14476
rect 14924 14399 14976 14408
rect 14924 14365 14939 14399
rect 14939 14365 14973 14399
rect 14973 14365 14976 14399
rect 14924 14356 14976 14365
rect 15660 14399 15712 14408
rect 15660 14365 15663 14399
rect 15663 14365 15697 14399
rect 15697 14365 15712 14399
rect 15660 14356 15712 14365
rect 15752 14356 15804 14408
rect 15936 14356 15988 14408
rect 15568 14288 15620 14340
rect 16028 14288 16080 14340
rect 16672 14399 16724 14408
rect 16672 14365 16681 14399
rect 16681 14365 16715 14399
rect 16715 14365 16724 14399
rect 16672 14356 16724 14365
rect 17684 14356 17736 14408
rect 17960 14399 18012 14408
rect 17960 14365 17969 14399
rect 17969 14365 18003 14399
rect 18003 14365 18012 14399
rect 17960 14356 18012 14365
rect 18144 14399 18196 14408
rect 18144 14365 18153 14399
rect 18153 14365 18187 14399
rect 18187 14365 18196 14399
rect 18144 14356 18196 14365
rect 18236 14356 18288 14408
rect 18512 14399 18564 14408
rect 18512 14365 18521 14399
rect 18521 14365 18555 14399
rect 18555 14365 18564 14399
rect 18512 14356 18564 14365
rect 19248 14399 19300 14408
rect 19248 14365 19257 14399
rect 19257 14365 19291 14399
rect 19291 14365 19300 14399
rect 19248 14356 19300 14365
rect 20076 14424 20128 14476
rect 20168 14399 20220 14408
rect 20168 14365 20177 14399
rect 20177 14365 20211 14399
rect 20211 14365 20220 14399
rect 20168 14356 20220 14365
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20260 14356 20312 14365
rect 20352 14399 20404 14408
rect 20352 14365 20361 14399
rect 20361 14365 20395 14399
rect 20395 14365 20404 14399
rect 20352 14356 20404 14365
rect 20536 14399 20588 14408
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 21364 14356 21416 14408
rect 21824 14399 21876 14408
rect 21824 14365 21833 14399
rect 21833 14365 21867 14399
rect 21867 14365 21876 14399
rect 21824 14356 21876 14365
rect 22468 14467 22520 14476
rect 22468 14433 22477 14467
rect 22477 14433 22511 14467
rect 22511 14433 22520 14467
rect 22468 14424 22520 14433
rect 25504 14424 25556 14476
rect 26148 14424 26200 14476
rect 23388 14399 23440 14408
rect 23388 14365 23397 14399
rect 23397 14365 23431 14399
rect 23431 14365 23440 14399
rect 23388 14356 23440 14365
rect 16948 14331 17000 14340
rect 16948 14297 16957 14331
rect 16957 14297 16991 14331
rect 16991 14297 17000 14331
rect 16948 14288 17000 14297
rect 10508 14263 10560 14272
rect 10508 14229 10517 14263
rect 10517 14229 10551 14263
rect 10551 14229 10560 14263
rect 10508 14220 10560 14229
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 15384 14220 15436 14272
rect 16488 14263 16540 14272
rect 16488 14229 16497 14263
rect 16497 14229 16531 14263
rect 16531 14229 16540 14263
rect 16488 14220 16540 14229
rect 16580 14220 16632 14272
rect 18052 14288 18104 14340
rect 19432 14288 19484 14340
rect 21088 14331 21140 14340
rect 21088 14297 21097 14331
rect 21097 14297 21131 14331
rect 21131 14297 21140 14331
rect 21088 14288 21140 14297
rect 22744 14288 22796 14340
rect 25136 14356 25188 14408
rect 25596 14399 25648 14408
rect 25596 14365 25605 14399
rect 25605 14365 25639 14399
rect 25639 14365 25648 14399
rect 25596 14356 25648 14365
rect 26056 14399 26108 14408
rect 26056 14365 26065 14399
rect 26065 14365 26099 14399
rect 26099 14365 26108 14399
rect 26056 14356 26108 14365
rect 26424 14356 26476 14408
rect 27160 14467 27212 14476
rect 27160 14433 27169 14467
rect 27169 14433 27203 14467
rect 27203 14433 27212 14467
rect 27160 14424 27212 14433
rect 34612 14288 34664 14340
rect 21272 14220 21324 14272
rect 23480 14220 23532 14272
rect 24676 14220 24728 14272
rect 25228 14263 25280 14272
rect 25228 14229 25237 14263
rect 25237 14229 25271 14263
rect 25271 14229 25280 14263
rect 25228 14220 25280 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 2320 14059 2372 14068
rect 2320 14025 2329 14059
rect 2329 14025 2363 14059
rect 2363 14025 2372 14059
rect 2320 14016 2372 14025
rect 8668 14016 8720 14068
rect 11612 14016 11664 14068
rect 14924 14016 14976 14068
rect 15568 14016 15620 14068
rect 15660 14016 15712 14068
rect 16212 14016 16264 14068
rect 16488 14016 16540 14068
rect 16764 14059 16816 14068
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 16856 14016 16908 14068
rect 17316 14016 17368 14068
rect 17960 14016 18012 14068
rect 18052 14059 18104 14068
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 18236 14016 18288 14068
rect 19524 14016 19576 14068
rect 3148 13880 3200 13932
rect 3976 13923 4028 13932
rect 3976 13889 3985 13923
rect 3985 13889 4019 13923
rect 4019 13889 4028 13923
rect 3976 13880 4028 13889
rect 4620 13812 4672 13864
rect 6184 13880 6236 13932
rect 8760 13880 8812 13932
rect 11888 13880 11940 13932
rect 13636 13880 13688 13932
rect 13912 13880 13964 13932
rect 11520 13812 11572 13864
rect 14556 13812 14608 13864
rect 16580 13812 16632 13864
rect 14188 13744 14240 13796
rect 15016 13744 15068 13796
rect 18420 13948 18472 14000
rect 20168 14016 20220 14068
rect 20260 14016 20312 14068
rect 20352 14016 20404 14068
rect 21640 14016 21692 14068
rect 22192 14059 22244 14068
rect 22192 14025 22201 14059
rect 22201 14025 22235 14059
rect 22235 14025 22244 14059
rect 22192 14016 22244 14025
rect 22284 14059 22336 14068
rect 22284 14025 22293 14059
rect 22293 14025 22327 14059
rect 22327 14025 22336 14059
rect 22284 14016 22336 14025
rect 22468 14059 22520 14068
rect 22468 14025 22477 14059
rect 22477 14025 22511 14059
rect 22511 14025 22520 14059
rect 22468 14016 22520 14025
rect 23112 14059 23164 14068
rect 23112 14025 23121 14059
rect 23121 14025 23155 14059
rect 23155 14025 23164 14059
rect 23112 14016 23164 14025
rect 24952 14016 25004 14068
rect 25688 14059 25740 14068
rect 25688 14025 25697 14059
rect 25697 14025 25731 14059
rect 25731 14025 25740 14059
rect 25688 14016 25740 14025
rect 31944 14059 31996 14068
rect 31944 14025 31953 14059
rect 31953 14025 31987 14059
rect 31987 14025 31996 14059
rect 31944 14016 31996 14025
rect 16948 13880 17000 13932
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 20536 13948 20588 14000
rect 24124 13991 24176 14000
rect 24124 13957 24133 13991
rect 24133 13957 24167 13991
rect 24167 13957 24176 13991
rect 24124 13948 24176 13957
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 22284 13880 22336 13932
rect 22560 13880 22612 13932
rect 20076 13812 20128 13864
rect 20260 13855 20312 13864
rect 20260 13821 20269 13855
rect 20269 13821 20303 13855
rect 20303 13821 20312 13855
rect 20260 13812 20312 13821
rect 20444 13812 20496 13864
rect 21916 13787 21968 13796
rect 21916 13753 21925 13787
rect 21925 13753 21959 13787
rect 21959 13753 21968 13787
rect 21916 13744 21968 13753
rect 3240 13676 3292 13728
rect 4068 13676 4120 13728
rect 4896 13676 4948 13728
rect 8760 13719 8812 13728
rect 8760 13685 8769 13719
rect 8769 13685 8803 13719
rect 8803 13685 8812 13719
rect 8760 13676 8812 13685
rect 12348 13676 12400 13728
rect 14648 13676 14700 13728
rect 14740 13719 14792 13728
rect 14740 13685 14749 13719
rect 14749 13685 14783 13719
rect 14783 13685 14792 13719
rect 14740 13676 14792 13685
rect 15200 13676 15252 13728
rect 19156 13676 19208 13728
rect 20352 13676 20404 13728
rect 23664 13812 23716 13864
rect 23940 13923 23992 13932
rect 23940 13889 23949 13923
rect 23949 13889 23983 13923
rect 23983 13889 23992 13923
rect 23940 13880 23992 13889
rect 24676 13923 24728 13932
rect 24676 13889 24685 13923
rect 24685 13889 24719 13923
rect 24719 13889 24728 13923
rect 24676 13880 24728 13889
rect 25044 13948 25096 14000
rect 34152 13948 34204 14000
rect 27804 13880 27856 13932
rect 24492 13855 24544 13864
rect 24492 13821 24501 13855
rect 24501 13821 24535 13855
rect 24535 13821 24544 13855
rect 24492 13812 24544 13821
rect 27988 13812 28040 13864
rect 31576 13923 31628 13932
rect 31576 13889 31585 13923
rect 31585 13889 31619 13923
rect 31619 13889 31628 13923
rect 31576 13880 31628 13889
rect 29828 13812 29880 13864
rect 31484 13812 31536 13864
rect 32220 13855 32272 13864
rect 32220 13821 32229 13855
rect 32229 13821 32263 13855
rect 32263 13821 32272 13855
rect 32220 13812 32272 13821
rect 32772 13812 32824 13864
rect 22560 13676 22612 13728
rect 23388 13676 23440 13728
rect 25228 13676 25280 13728
rect 29092 13676 29144 13728
rect 31760 13676 31812 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4620 13472 4672 13524
rect 1400 13379 1452 13388
rect 1400 13345 1409 13379
rect 1409 13345 1443 13379
rect 1443 13345 1452 13379
rect 1400 13336 1452 13345
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 2412 13200 2464 13252
rect 3148 13175 3200 13184
rect 3148 13141 3157 13175
rect 3157 13141 3191 13175
rect 3191 13141 3200 13175
rect 3148 13132 3200 13141
rect 4804 13404 4856 13456
rect 4896 13404 4948 13456
rect 4252 13268 4304 13320
rect 4344 13268 4396 13320
rect 3608 13200 3660 13252
rect 4068 13243 4120 13252
rect 4068 13209 4077 13243
rect 4077 13209 4111 13243
rect 4111 13209 4120 13243
rect 4068 13200 4120 13209
rect 3884 13132 3936 13184
rect 5080 13268 5132 13320
rect 5172 13311 5224 13320
rect 5172 13277 5181 13311
rect 5181 13277 5215 13311
rect 5215 13277 5224 13311
rect 5172 13268 5224 13277
rect 5264 13311 5316 13320
rect 5264 13277 5273 13311
rect 5273 13277 5307 13311
rect 5307 13277 5316 13311
rect 5264 13268 5316 13277
rect 5356 13311 5408 13320
rect 5356 13277 5365 13311
rect 5365 13277 5399 13311
rect 5399 13277 5408 13311
rect 5356 13268 5408 13277
rect 14648 13472 14700 13524
rect 14740 13472 14792 13524
rect 16120 13472 16172 13524
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 16948 13472 17000 13524
rect 17040 13472 17092 13524
rect 17592 13472 17644 13524
rect 18236 13472 18288 13524
rect 19248 13472 19300 13524
rect 19524 13515 19576 13524
rect 19524 13481 19533 13515
rect 19533 13481 19567 13515
rect 19567 13481 19576 13515
rect 19524 13472 19576 13481
rect 20444 13472 20496 13524
rect 20996 13472 21048 13524
rect 21640 13515 21692 13524
rect 21640 13481 21649 13515
rect 21649 13481 21683 13515
rect 21683 13481 21692 13515
rect 21640 13472 21692 13481
rect 15936 13404 15988 13456
rect 8668 13268 8720 13320
rect 8944 13311 8996 13320
rect 8944 13277 8953 13311
rect 8953 13277 8987 13311
rect 8987 13277 8996 13311
rect 8944 13268 8996 13277
rect 12164 13336 12216 13388
rect 11428 13311 11480 13320
rect 11428 13277 11437 13311
rect 11437 13277 11471 13311
rect 11471 13277 11480 13311
rect 11428 13268 11480 13277
rect 4620 13200 4672 13252
rect 9680 13200 9732 13252
rect 12440 13268 12492 13320
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 14648 13268 14700 13320
rect 15384 13336 15436 13388
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 16580 13311 16632 13320
rect 16580 13277 16589 13311
rect 16589 13277 16623 13311
rect 16623 13277 16632 13311
rect 16580 13268 16632 13277
rect 19432 13404 19484 13456
rect 17868 13336 17920 13388
rect 16948 13311 17000 13320
rect 16948 13277 16957 13311
rect 16957 13277 16991 13311
rect 16991 13277 17000 13311
rect 16948 13268 17000 13277
rect 17132 13311 17184 13320
rect 17132 13277 17141 13311
rect 17141 13277 17175 13311
rect 17175 13277 17184 13311
rect 17132 13268 17184 13277
rect 18052 13268 18104 13320
rect 18236 13268 18288 13320
rect 18420 13268 18472 13320
rect 19156 13336 19208 13388
rect 21916 13472 21968 13524
rect 22652 13472 22704 13524
rect 23112 13472 23164 13524
rect 23664 13515 23716 13524
rect 23664 13481 23673 13515
rect 23673 13481 23707 13515
rect 23707 13481 23716 13515
rect 23664 13472 23716 13481
rect 27252 13515 27304 13524
rect 27252 13481 27261 13515
rect 27261 13481 27295 13515
rect 27295 13481 27304 13515
rect 27252 13472 27304 13481
rect 28540 13515 28592 13524
rect 28540 13481 28549 13515
rect 28549 13481 28583 13515
rect 28583 13481 28592 13515
rect 28540 13472 28592 13481
rect 31484 13515 31536 13524
rect 31484 13481 31493 13515
rect 31493 13481 31527 13515
rect 31527 13481 31536 13515
rect 31484 13472 31536 13481
rect 32220 13472 32272 13524
rect 34152 13515 34204 13524
rect 34152 13481 34161 13515
rect 34161 13481 34195 13515
rect 34195 13481 34204 13515
rect 34152 13472 34204 13481
rect 22008 13404 22060 13456
rect 24492 13404 24544 13456
rect 29092 13379 29144 13388
rect 29092 13345 29101 13379
rect 29101 13345 29135 13379
rect 29135 13345 29144 13379
rect 29092 13336 29144 13345
rect 29368 13336 29420 13388
rect 18512 13243 18564 13252
rect 18512 13209 18521 13243
rect 18521 13209 18555 13243
rect 18555 13209 18564 13243
rect 18512 13200 18564 13209
rect 20536 13268 20588 13320
rect 5264 13132 5316 13184
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13084 13132 13136 13141
rect 17040 13132 17092 13184
rect 18144 13132 18196 13184
rect 19340 13200 19392 13252
rect 20260 13243 20312 13252
rect 20260 13209 20269 13243
rect 20269 13209 20303 13243
rect 20303 13209 20312 13243
rect 21364 13268 21416 13320
rect 23572 13268 23624 13320
rect 27436 13311 27488 13320
rect 27436 13277 27445 13311
rect 27445 13277 27479 13311
rect 27479 13277 27488 13311
rect 27436 13268 27488 13277
rect 20260 13200 20312 13209
rect 23940 13200 23992 13252
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 27988 13200 28040 13252
rect 28264 13311 28316 13320
rect 28264 13277 28273 13311
rect 28273 13277 28307 13311
rect 28307 13277 28316 13311
rect 28264 13268 28316 13277
rect 28356 13311 28408 13320
rect 28356 13277 28365 13311
rect 28365 13277 28399 13311
rect 28399 13277 28408 13311
rect 28356 13268 28408 13277
rect 29000 13311 29052 13320
rect 29000 13277 29009 13311
rect 29009 13277 29043 13311
rect 29043 13277 29052 13311
rect 29000 13268 29052 13277
rect 31760 13404 31812 13456
rect 31668 13268 31720 13320
rect 22560 13175 22612 13184
rect 22560 13141 22569 13175
rect 22569 13141 22603 13175
rect 22603 13141 22612 13175
rect 22560 13132 22612 13141
rect 23296 13175 23348 13184
rect 23296 13141 23305 13175
rect 23305 13141 23339 13175
rect 23339 13141 23348 13175
rect 23296 13132 23348 13141
rect 27252 13132 27304 13184
rect 28080 13132 28132 13184
rect 30748 13200 30800 13252
rect 31392 13132 31444 13184
rect 31944 13132 31996 13184
rect 34704 13132 34756 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 1676 12928 1728 12980
rect 2412 12971 2464 12980
rect 2412 12937 2421 12971
rect 2421 12937 2455 12971
rect 2455 12937 2464 12971
rect 2412 12928 2464 12937
rect 2872 12971 2924 12980
rect 940 12792 992 12844
rect 2872 12937 2881 12971
rect 2881 12937 2915 12971
rect 2915 12937 2924 12971
rect 2872 12928 2924 12937
rect 3332 12928 3384 12980
rect 3884 12971 3936 12980
rect 3884 12937 3893 12971
rect 3893 12937 3927 12971
rect 3927 12937 3936 12971
rect 3884 12928 3936 12937
rect 3976 12860 4028 12912
rect 5356 12928 5408 12980
rect 5172 12860 5224 12912
rect 3148 12792 3200 12844
rect 4252 12835 4304 12844
rect 4252 12801 4261 12835
rect 4261 12801 4295 12835
rect 4295 12801 4304 12835
rect 4252 12792 4304 12801
rect 4620 12792 4672 12844
rect 5264 12792 5316 12844
rect 8392 12860 8444 12912
rect 8944 12928 8996 12980
rect 9680 12928 9732 12980
rect 8944 12792 8996 12844
rect 10508 12903 10560 12912
rect 10508 12869 10517 12903
rect 10517 12869 10551 12903
rect 10551 12869 10560 12903
rect 10508 12860 10560 12869
rect 12532 12928 12584 12980
rect 4712 12656 4764 12708
rect 9588 12724 9640 12776
rect 4068 12588 4120 12640
rect 4344 12588 4396 12640
rect 5080 12588 5132 12640
rect 11520 12792 11572 12844
rect 14648 12928 14700 12980
rect 15292 12928 15344 12980
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 17500 12928 17552 12980
rect 17592 12928 17644 12980
rect 18512 12928 18564 12980
rect 19156 12971 19208 12980
rect 19156 12937 19165 12971
rect 19165 12937 19199 12971
rect 19199 12937 19208 12971
rect 19156 12928 19208 12937
rect 19248 12928 19300 12980
rect 19432 12928 19484 12980
rect 19800 12928 19852 12980
rect 21088 12928 21140 12980
rect 21364 12928 21416 12980
rect 22744 12971 22796 12980
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 13636 12835 13688 12844
rect 13636 12801 13645 12835
rect 13645 12801 13679 12835
rect 13679 12801 13688 12835
rect 13636 12792 13688 12801
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 12532 12767 12584 12776
rect 12532 12733 12541 12767
rect 12541 12733 12575 12767
rect 12575 12733 12584 12767
rect 12532 12724 12584 12733
rect 10048 12588 10100 12640
rect 14096 12835 14148 12844
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 15108 12792 15160 12844
rect 15936 12792 15988 12844
rect 14464 12656 14516 12708
rect 14648 12767 14700 12776
rect 14648 12733 14657 12767
rect 14657 12733 14691 12767
rect 14691 12733 14700 12767
rect 14648 12724 14700 12733
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 15752 12724 15804 12776
rect 16396 12835 16448 12844
rect 16396 12801 16405 12835
rect 16405 12801 16439 12835
rect 16439 12801 16448 12835
rect 16396 12792 16448 12801
rect 17040 12835 17092 12844
rect 17040 12801 17049 12835
rect 17049 12801 17083 12835
rect 17083 12801 17092 12835
rect 17040 12792 17092 12801
rect 17316 12835 17368 12844
rect 17316 12801 17325 12835
rect 17325 12801 17359 12835
rect 17359 12801 17368 12835
rect 17316 12792 17368 12801
rect 17868 12835 17920 12844
rect 17868 12801 17877 12835
rect 17877 12801 17911 12835
rect 17911 12801 17920 12835
rect 17868 12792 17920 12801
rect 18420 12792 18472 12844
rect 20996 12903 21048 12912
rect 20996 12869 21005 12903
rect 21005 12869 21039 12903
rect 21039 12869 21048 12903
rect 20996 12860 21048 12869
rect 18696 12724 18748 12776
rect 19064 12792 19116 12844
rect 19340 12792 19392 12844
rect 19984 12835 20036 12844
rect 19984 12801 19993 12835
rect 19993 12801 20027 12835
rect 20027 12801 20036 12835
rect 19984 12792 20036 12801
rect 22744 12937 22753 12971
rect 22753 12937 22787 12971
rect 22787 12937 22796 12971
rect 22744 12928 22796 12937
rect 23204 12928 23256 12980
rect 25228 12928 25280 12980
rect 27068 12928 27120 12980
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 15476 12656 15528 12708
rect 16488 12656 16540 12708
rect 19432 12656 19484 12708
rect 15016 12588 15068 12640
rect 15752 12588 15804 12640
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 18236 12588 18288 12640
rect 18328 12631 18380 12640
rect 18328 12597 18337 12631
rect 18337 12597 18371 12631
rect 18371 12597 18380 12631
rect 18328 12588 18380 12597
rect 22560 12792 22612 12844
rect 23664 12792 23716 12844
rect 22100 12767 22152 12776
rect 22100 12733 22109 12767
rect 22109 12733 22143 12767
rect 22143 12733 22152 12767
rect 22100 12724 22152 12733
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24492 12792 24544 12801
rect 25044 12835 25096 12844
rect 25044 12801 25053 12835
rect 25053 12801 25087 12835
rect 25087 12801 25096 12835
rect 25044 12792 25096 12801
rect 25136 12767 25188 12776
rect 25136 12733 25145 12767
rect 25145 12733 25179 12767
rect 25179 12733 25188 12767
rect 25136 12724 25188 12733
rect 22836 12656 22888 12708
rect 25872 12724 25924 12776
rect 26884 12860 26936 12912
rect 28264 12928 28316 12980
rect 29000 12928 29052 12980
rect 29368 12928 29420 12980
rect 29736 12928 29788 12980
rect 30656 12928 30708 12980
rect 30748 12971 30800 12980
rect 30748 12937 30757 12971
rect 30757 12937 30791 12971
rect 30791 12937 30800 12971
rect 30748 12928 30800 12937
rect 31392 12928 31444 12980
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 27252 12792 27304 12801
rect 27712 12860 27764 12912
rect 26792 12724 26844 12776
rect 28080 12724 28132 12776
rect 28356 12767 28408 12776
rect 28356 12733 28365 12767
rect 28365 12733 28399 12767
rect 28399 12733 28408 12767
rect 28356 12724 28408 12733
rect 27620 12656 27672 12708
rect 22192 12588 22244 12640
rect 22652 12588 22704 12640
rect 23388 12588 23440 12640
rect 23480 12631 23532 12640
rect 23480 12597 23489 12631
rect 23489 12597 23523 12631
rect 23523 12597 23532 12631
rect 23480 12588 23532 12597
rect 26056 12588 26108 12640
rect 26700 12588 26752 12640
rect 27252 12588 27304 12640
rect 31668 12860 31720 12912
rect 31760 12835 31812 12844
rect 31760 12801 31769 12835
rect 31769 12801 31803 12835
rect 31803 12801 31812 12835
rect 31760 12792 31812 12801
rect 31944 12835 31996 12844
rect 31944 12801 31953 12835
rect 31953 12801 31987 12835
rect 31987 12801 31996 12835
rect 31944 12792 31996 12801
rect 32680 12699 32732 12708
rect 32680 12665 32689 12699
rect 32689 12665 32723 12699
rect 32723 12665 32732 12699
rect 32680 12656 32732 12665
rect 34704 12588 34756 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 4068 12384 4120 12436
rect 8392 12384 8444 12436
rect 3332 12316 3384 12368
rect 1400 12291 1452 12300
rect 1400 12257 1409 12291
rect 1409 12257 1443 12291
rect 1443 12257 1452 12291
rect 1400 12248 1452 12257
rect 4620 12180 4672 12232
rect 1676 12155 1728 12164
rect 1676 12121 1685 12155
rect 1685 12121 1719 12155
rect 1719 12121 1728 12155
rect 1676 12112 1728 12121
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 8760 12384 8812 12436
rect 10048 12384 10100 12436
rect 11520 12427 11572 12436
rect 11520 12393 11529 12427
rect 11529 12393 11563 12427
rect 11563 12393 11572 12427
rect 11520 12384 11572 12393
rect 14096 12427 14148 12436
rect 14096 12393 14105 12427
rect 14105 12393 14139 12427
rect 14139 12393 14148 12427
rect 14096 12384 14148 12393
rect 15108 12384 15160 12436
rect 16212 12384 16264 12436
rect 14372 12316 14424 12368
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 13912 12180 13964 12232
rect 14464 12180 14516 12232
rect 14924 12291 14976 12300
rect 14924 12257 14933 12291
rect 14933 12257 14967 12291
rect 14967 12257 14976 12291
rect 14924 12248 14976 12257
rect 16580 12316 16632 12368
rect 14740 12180 14792 12232
rect 15568 12291 15620 12300
rect 15568 12257 15577 12291
rect 15577 12257 15611 12291
rect 15611 12257 15620 12291
rect 15568 12248 15620 12257
rect 15660 12291 15712 12300
rect 15660 12257 15669 12291
rect 15669 12257 15703 12291
rect 15703 12257 15712 12291
rect 15660 12248 15712 12257
rect 15752 12180 15804 12232
rect 15936 12180 15988 12232
rect 17500 12427 17552 12436
rect 17500 12393 17509 12427
rect 17509 12393 17543 12427
rect 17543 12393 17552 12427
rect 17500 12384 17552 12393
rect 17960 12384 18012 12436
rect 18420 12384 18472 12436
rect 19984 12384 20036 12436
rect 16856 12223 16908 12232
rect 16856 12189 16865 12223
rect 16865 12189 16899 12223
rect 16899 12189 16908 12223
rect 16856 12180 16908 12189
rect 17960 12248 18012 12300
rect 19800 12291 19852 12300
rect 7196 12087 7248 12096
rect 7196 12053 7205 12087
rect 7205 12053 7239 12087
rect 7239 12053 7248 12087
rect 7196 12044 7248 12053
rect 13636 12044 13688 12096
rect 16580 12112 16632 12164
rect 16764 12112 16816 12164
rect 17224 12180 17276 12232
rect 18512 12180 18564 12232
rect 18696 12223 18748 12232
rect 18696 12189 18705 12223
rect 18705 12189 18739 12223
rect 18739 12189 18748 12223
rect 18696 12180 18748 12189
rect 19800 12257 19809 12291
rect 19809 12257 19843 12291
rect 19843 12257 19852 12291
rect 19800 12248 19852 12257
rect 20076 12248 20128 12300
rect 18236 12112 18288 12164
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 21732 12180 21784 12232
rect 22836 12384 22888 12436
rect 23296 12384 23348 12436
rect 23388 12384 23440 12436
rect 22008 12180 22060 12232
rect 22468 12180 22520 12232
rect 22744 12223 22796 12232
rect 22744 12189 22753 12223
rect 22753 12189 22787 12223
rect 22787 12189 22796 12223
rect 22744 12180 22796 12189
rect 23204 12223 23256 12232
rect 23204 12189 23213 12223
rect 23213 12189 23247 12223
rect 23247 12189 23256 12223
rect 23204 12180 23256 12189
rect 22100 12112 22152 12164
rect 23848 12248 23900 12300
rect 23388 12223 23440 12232
rect 23388 12189 23397 12223
rect 23397 12189 23431 12223
rect 23431 12189 23440 12223
rect 23388 12180 23440 12189
rect 25228 12384 25280 12436
rect 25872 12316 25924 12368
rect 18788 12044 18840 12096
rect 19340 12044 19392 12096
rect 20260 12044 20312 12096
rect 21088 12044 21140 12096
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 22928 12044 22980 12096
rect 23572 12044 23624 12096
rect 23848 12087 23900 12096
rect 23848 12053 23857 12087
rect 23857 12053 23891 12087
rect 23891 12053 23900 12087
rect 23848 12044 23900 12053
rect 23940 12087 23992 12096
rect 23940 12053 23949 12087
rect 23949 12053 23983 12087
rect 23983 12053 23992 12087
rect 23940 12044 23992 12053
rect 24216 12112 24268 12164
rect 25688 12180 25740 12232
rect 25320 12155 25372 12164
rect 25320 12121 25329 12155
rect 25329 12121 25363 12155
rect 25363 12121 25372 12155
rect 26056 12223 26108 12232
rect 26056 12189 26065 12223
rect 26065 12189 26099 12223
rect 26099 12189 26108 12223
rect 26056 12180 26108 12189
rect 27436 12384 27488 12436
rect 32680 12384 32732 12436
rect 26792 12180 26844 12232
rect 26884 12223 26936 12232
rect 26884 12189 26893 12223
rect 26893 12189 26927 12223
rect 26927 12189 26936 12223
rect 26884 12180 26936 12189
rect 29828 12291 29880 12300
rect 29828 12257 29837 12291
rect 29837 12257 29871 12291
rect 29871 12257 29880 12291
rect 29828 12248 29880 12257
rect 27160 12180 27212 12232
rect 27528 12180 27580 12232
rect 25320 12112 25372 12121
rect 30932 12180 30984 12232
rect 32772 12223 32824 12232
rect 32772 12189 32781 12223
rect 32781 12189 32815 12223
rect 32815 12189 32824 12223
rect 32772 12180 32824 12189
rect 34704 12223 34756 12232
rect 34704 12189 34713 12223
rect 34713 12189 34747 12223
rect 34747 12189 34756 12223
rect 34704 12180 34756 12189
rect 26700 12044 26752 12096
rect 29736 12112 29788 12164
rect 27068 12044 27120 12096
rect 27712 12044 27764 12096
rect 31300 12087 31352 12096
rect 31300 12053 31309 12087
rect 31309 12053 31343 12087
rect 31343 12053 31352 12087
rect 31300 12044 31352 12053
rect 34520 12087 34572 12096
rect 34520 12053 34529 12087
rect 34529 12053 34563 12087
rect 34563 12053 34572 12087
rect 34520 12044 34572 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4620 11840 4672 11892
rect 7196 11840 7248 11892
rect 13084 11883 13136 11892
rect 13084 11849 13093 11883
rect 13093 11849 13127 11883
rect 13127 11849 13136 11883
rect 13084 11840 13136 11849
rect 13360 11883 13412 11892
rect 13360 11849 13369 11883
rect 13369 11849 13403 11883
rect 13403 11849 13412 11883
rect 13360 11840 13412 11849
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 12348 11772 12400 11824
rect 1400 11704 1452 11756
rect 3884 11704 3936 11756
rect 10048 11704 10100 11756
rect 2780 11679 2832 11688
rect 2780 11645 2789 11679
rect 2789 11645 2823 11679
rect 2823 11645 2832 11679
rect 2780 11636 2832 11645
rect 4620 11679 4672 11688
rect 4620 11645 4629 11679
rect 4629 11645 4663 11679
rect 4663 11645 4672 11679
rect 4620 11636 4672 11645
rect 15568 11704 15620 11756
rect 16028 11747 16080 11756
rect 16028 11713 16037 11747
rect 16037 11713 16071 11747
rect 16071 11713 16080 11747
rect 16028 11704 16080 11713
rect 16396 11704 16448 11756
rect 17868 11840 17920 11892
rect 19432 11840 19484 11892
rect 20628 11840 20680 11892
rect 20996 11772 21048 11824
rect 22192 11883 22244 11892
rect 22192 11849 22201 11883
rect 22201 11849 22235 11883
rect 22235 11849 22244 11883
rect 22192 11840 22244 11849
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 23204 11840 23256 11892
rect 23572 11840 23624 11892
rect 24768 11840 24820 11892
rect 26516 11840 26568 11892
rect 27068 11840 27120 11892
rect 27620 11883 27672 11892
rect 27620 11849 27629 11883
rect 27629 11849 27663 11883
rect 27663 11849 27672 11883
rect 27620 11840 27672 11849
rect 27712 11840 27764 11892
rect 27988 11840 28040 11892
rect 9588 11568 9640 11620
rect 10048 11543 10100 11552
rect 10048 11509 10057 11543
rect 10057 11509 10091 11543
rect 10091 11509 10100 11543
rect 10048 11500 10100 11509
rect 16120 11568 16172 11620
rect 18420 11747 18472 11756
rect 18420 11713 18429 11747
rect 18429 11713 18463 11747
rect 18463 11713 18472 11747
rect 18420 11704 18472 11713
rect 18512 11704 18564 11756
rect 20352 11704 20404 11756
rect 21088 11747 21140 11756
rect 21088 11713 21097 11747
rect 21097 11713 21131 11747
rect 21131 11713 21140 11747
rect 21088 11704 21140 11713
rect 21732 11704 21784 11756
rect 23940 11772 23992 11824
rect 26700 11772 26752 11824
rect 18788 11679 18840 11688
rect 18788 11645 18797 11679
rect 18797 11645 18831 11679
rect 18831 11645 18840 11679
rect 18788 11636 18840 11645
rect 20076 11568 20128 11620
rect 21364 11611 21416 11620
rect 21364 11577 21373 11611
rect 21373 11577 21407 11611
rect 21407 11577 21416 11611
rect 21364 11568 21416 11577
rect 22468 11679 22520 11688
rect 22468 11645 22477 11679
rect 22477 11645 22511 11679
rect 22511 11645 22520 11679
rect 22468 11636 22520 11645
rect 25964 11704 26016 11756
rect 27068 11704 27120 11756
rect 22836 11636 22888 11688
rect 25320 11636 25372 11688
rect 28080 11747 28132 11756
rect 28080 11713 28089 11747
rect 28089 11713 28123 11747
rect 28123 11713 28132 11747
rect 28080 11704 28132 11713
rect 29000 11840 29052 11892
rect 29736 11840 29788 11892
rect 30932 11883 30984 11892
rect 30932 11849 30941 11883
rect 30941 11849 30975 11883
rect 30975 11849 30984 11883
rect 30932 11840 30984 11849
rect 31944 11840 31996 11892
rect 34520 11840 34572 11892
rect 31300 11772 31352 11824
rect 31576 11772 31628 11824
rect 22928 11568 22980 11620
rect 18328 11543 18380 11552
rect 18328 11509 18337 11543
rect 18337 11509 18371 11543
rect 18371 11509 18380 11543
rect 18328 11500 18380 11509
rect 19340 11500 19392 11552
rect 20352 11543 20404 11552
rect 20352 11509 20361 11543
rect 20361 11509 20395 11543
rect 20395 11509 20404 11543
rect 20352 11500 20404 11509
rect 21180 11500 21232 11552
rect 22284 11500 22336 11552
rect 22744 11500 22796 11552
rect 23296 11500 23348 11552
rect 25688 11500 25740 11552
rect 26700 11500 26752 11552
rect 27252 11500 27304 11552
rect 27896 11636 27948 11688
rect 30380 11704 30432 11756
rect 27804 11568 27856 11620
rect 31484 11636 31536 11688
rect 34796 11704 34848 11756
rect 30472 11543 30524 11552
rect 30472 11509 30481 11543
rect 30481 11509 30515 11543
rect 30515 11509 30524 11543
rect 30472 11500 30524 11509
rect 31852 11543 31904 11552
rect 31852 11509 31861 11543
rect 31861 11509 31895 11543
rect 31895 11509 31904 11543
rect 31852 11500 31904 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 17960 11296 18012 11348
rect 18420 11296 18472 11348
rect 18512 11339 18564 11348
rect 18512 11305 18521 11339
rect 18521 11305 18555 11339
rect 18555 11305 18564 11339
rect 18512 11296 18564 11305
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 22192 11296 22244 11348
rect 22560 11296 22612 11348
rect 23940 11296 23992 11348
rect 24216 11339 24268 11348
rect 24216 11305 24225 11339
rect 24225 11305 24259 11339
rect 24259 11305 24268 11339
rect 24216 11296 24268 11305
rect 25320 11296 25372 11348
rect 27712 11296 27764 11348
rect 28356 11296 28408 11348
rect 29000 11296 29052 11348
rect 30472 11296 30524 11348
rect 31484 11339 31536 11348
rect 31484 11305 31493 11339
rect 31493 11305 31527 11339
rect 31527 11305 31536 11339
rect 31484 11296 31536 11305
rect 31760 11339 31812 11348
rect 31760 11305 31769 11339
rect 31769 11305 31803 11339
rect 31803 11305 31812 11339
rect 31760 11296 31812 11305
rect 31852 11296 31904 11348
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 21180 11228 21232 11280
rect 22100 11228 22152 11280
rect 22836 11228 22888 11280
rect 22008 11092 22060 11144
rect 22284 11135 22336 11144
rect 22284 11101 22293 11135
rect 22293 11101 22327 11135
rect 22327 11101 22336 11135
rect 22284 11092 22336 11101
rect 22376 11092 22428 11144
rect 22836 11092 22888 11144
rect 24676 11228 24728 11280
rect 27896 11228 27948 11280
rect 28080 11228 28132 11280
rect 9588 11067 9640 11076
rect 9588 11033 9597 11067
rect 9597 11033 9631 11067
rect 9631 11033 9640 11067
rect 9588 11024 9640 11033
rect 19340 11024 19392 11076
rect 20444 11067 20496 11076
rect 20444 11033 20453 11067
rect 20453 11033 20487 11067
rect 20487 11033 20496 11067
rect 20444 11024 20496 11033
rect 22652 11024 22704 11076
rect 23664 11092 23716 11144
rect 24032 11092 24084 11144
rect 24400 11135 24452 11144
rect 24400 11101 24409 11135
rect 24409 11101 24443 11135
rect 24443 11101 24452 11135
rect 24400 11092 24452 11101
rect 24492 11092 24544 11144
rect 23572 11024 23624 11076
rect 24768 11135 24820 11144
rect 24768 11101 24777 11135
rect 24777 11101 24811 11135
rect 24811 11101 24820 11135
rect 24768 11092 24820 11101
rect 25504 11135 25556 11144
rect 25504 11101 25513 11135
rect 25513 11101 25547 11135
rect 25547 11101 25556 11135
rect 25504 11092 25556 11101
rect 24676 11024 24728 11076
rect 26700 11092 26752 11144
rect 27252 11135 27304 11144
rect 27252 11101 27261 11135
rect 27261 11101 27295 11135
rect 27295 11101 27304 11135
rect 27252 11092 27304 11101
rect 27620 11135 27672 11144
rect 27620 11101 27629 11135
rect 27629 11101 27663 11135
rect 27663 11101 27672 11135
rect 27620 11092 27672 11101
rect 34612 11160 34664 11212
rect 31576 11135 31628 11144
rect 31576 11101 31585 11135
rect 31585 11101 31619 11135
rect 31619 11101 31628 11135
rect 31576 11092 31628 11101
rect 31760 11092 31812 11144
rect 32772 11135 32824 11144
rect 32772 11101 32781 11135
rect 32781 11101 32815 11135
rect 32815 11101 32824 11135
rect 32772 11092 32824 11101
rect 34704 11135 34756 11144
rect 34704 11101 34713 11135
rect 34713 11101 34747 11135
rect 34747 11101 34756 11135
rect 34704 11092 34756 11101
rect 30380 11067 30432 11076
rect 30380 11033 30389 11067
rect 30389 11033 30423 11067
rect 30423 11033 30432 11067
rect 30380 11024 30432 11033
rect 31116 11024 31168 11076
rect 19432 10956 19484 11008
rect 28908 10956 28960 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 10600 10795 10652 10804
rect 10600 10761 10609 10795
rect 10609 10761 10643 10795
rect 10643 10761 10652 10795
rect 10600 10752 10652 10761
rect 19340 10752 19392 10804
rect 20996 10752 21048 10804
rect 22100 10752 22152 10804
rect 19984 10684 20036 10736
rect 3240 10616 3292 10668
rect 18696 10659 18748 10668
rect 18696 10625 18705 10659
rect 18705 10625 18739 10659
rect 18739 10625 18748 10659
rect 18696 10616 18748 10625
rect 19248 10659 19300 10668
rect 19248 10625 19257 10659
rect 19257 10625 19291 10659
rect 19291 10625 19300 10659
rect 19248 10616 19300 10625
rect 20444 10659 20496 10668
rect 20444 10625 20453 10659
rect 20453 10625 20487 10659
rect 20487 10625 20496 10659
rect 20444 10616 20496 10625
rect 19984 10548 20036 10600
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 22652 10684 22704 10736
rect 21180 10591 21232 10600
rect 21180 10557 21189 10591
rect 21189 10557 21223 10591
rect 21223 10557 21232 10591
rect 21180 10548 21232 10557
rect 21272 10548 21324 10600
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 23020 10659 23072 10668
rect 23020 10625 23029 10659
rect 23029 10625 23063 10659
rect 23063 10625 23072 10659
rect 23020 10616 23072 10625
rect 23848 10752 23900 10804
rect 25504 10752 25556 10804
rect 25780 10752 25832 10804
rect 27528 10752 27580 10804
rect 29000 10752 29052 10804
rect 29368 10795 29420 10804
rect 29368 10761 29377 10795
rect 29377 10761 29411 10795
rect 29411 10761 29420 10795
rect 29368 10752 29420 10761
rect 24400 10684 24452 10736
rect 24492 10684 24544 10736
rect 22468 10548 22520 10600
rect 23572 10616 23624 10668
rect 24676 10659 24728 10668
rect 24676 10625 24685 10659
rect 24685 10625 24719 10659
rect 24719 10625 24728 10659
rect 24676 10616 24728 10625
rect 26516 10684 26568 10736
rect 23664 10548 23716 10600
rect 24216 10591 24268 10600
rect 24216 10557 24225 10591
rect 24225 10557 24259 10591
rect 24259 10557 24268 10591
rect 24216 10548 24268 10557
rect 22744 10480 22796 10532
rect 25044 10616 25096 10668
rect 25228 10591 25280 10600
rect 25228 10557 25237 10591
rect 25237 10557 25271 10591
rect 25271 10557 25280 10591
rect 25964 10659 26016 10668
rect 25964 10625 25973 10659
rect 25973 10625 26007 10659
rect 26007 10625 26016 10659
rect 25964 10616 26016 10625
rect 25228 10548 25280 10557
rect 17224 10412 17276 10464
rect 20536 10455 20588 10464
rect 20536 10421 20545 10455
rect 20545 10421 20579 10455
rect 20579 10421 20588 10455
rect 20536 10412 20588 10421
rect 20812 10455 20864 10464
rect 20812 10421 20821 10455
rect 20821 10421 20855 10455
rect 20855 10421 20864 10455
rect 20812 10412 20864 10421
rect 22284 10412 22336 10464
rect 25044 10455 25096 10464
rect 25044 10421 25053 10455
rect 25053 10421 25087 10455
rect 25087 10421 25096 10455
rect 25044 10412 25096 10421
rect 28908 10616 28960 10668
rect 31484 10616 31536 10668
rect 31576 10659 31628 10668
rect 31576 10625 31585 10659
rect 31585 10625 31619 10659
rect 31619 10625 31628 10659
rect 31576 10616 31628 10625
rect 31760 10659 31812 10668
rect 31760 10625 31769 10659
rect 31769 10625 31803 10659
rect 31803 10625 31812 10659
rect 31760 10616 31812 10625
rect 31944 10752 31996 10804
rect 32772 10752 32824 10804
rect 32220 10616 32272 10668
rect 26332 10523 26384 10532
rect 26332 10489 26341 10523
rect 26341 10489 26375 10523
rect 26375 10489 26384 10523
rect 26332 10480 26384 10489
rect 27252 10591 27304 10600
rect 27252 10557 27261 10591
rect 27261 10557 27295 10591
rect 27295 10557 27304 10591
rect 27252 10548 27304 10557
rect 31300 10480 31352 10532
rect 27528 10412 27580 10464
rect 30104 10455 30156 10464
rect 30104 10421 30113 10455
rect 30113 10421 30147 10455
rect 30147 10421 30156 10455
rect 30104 10412 30156 10421
rect 31392 10455 31444 10464
rect 31392 10421 31401 10455
rect 31401 10421 31435 10455
rect 31435 10421 31444 10455
rect 31392 10412 31444 10421
rect 34060 10412 34112 10464
rect 34704 10412 34756 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4620 10208 4672 10260
rect 18696 10251 18748 10260
rect 18696 10217 18705 10251
rect 18705 10217 18739 10251
rect 18739 10217 18748 10251
rect 18696 10208 18748 10217
rect 19248 10208 19300 10260
rect 19984 10251 20036 10260
rect 19984 10217 19993 10251
rect 19993 10217 20027 10251
rect 20027 10217 20036 10251
rect 19984 10208 20036 10217
rect 20536 10208 20588 10260
rect 20812 10208 20864 10260
rect 21272 10251 21324 10260
rect 21272 10217 21281 10251
rect 21281 10217 21315 10251
rect 21315 10217 21324 10251
rect 21272 10208 21324 10217
rect 22008 10251 22060 10260
rect 22008 10217 22017 10251
rect 22017 10217 22051 10251
rect 22051 10217 22060 10251
rect 22008 10208 22060 10217
rect 22836 10251 22888 10260
rect 22836 10217 22845 10251
rect 22845 10217 22879 10251
rect 22879 10217 22888 10251
rect 22836 10208 22888 10217
rect 23020 10208 23072 10260
rect 24032 10208 24084 10260
rect 24216 10208 24268 10260
rect 25228 10208 25280 10260
rect 26148 10208 26200 10260
rect 18328 10072 18380 10124
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 22560 10115 22612 10124
rect 22560 10081 22569 10115
rect 22569 10081 22603 10115
rect 22603 10081 22612 10115
rect 22560 10072 22612 10081
rect 23572 10072 23624 10124
rect 1400 9936 1452 9988
rect 2872 9936 2924 9988
rect 22008 10004 22060 10056
rect 22468 10047 22520 10056
rect 22468 10013 22477 10047
rect 22477 10013 22511 10047
rect 22511 10013 22520 10047
rect 22468 10004 22520 10013
rect 23664 10004 23716 10056
rect 24032 10004 24084 10056
rect 24124 10047 24176 10056
rect 24124 10013 24133 10047
rect 24133 10013 24167 10047
rect 24167 10013 24176 10047
rect 24124 10004 24176 10013
rect 25044 10004 25096 10056
rect 25780 10004 25832 10056
rect 18604 9868 18656 9920
rect 20352 9868 20404 9920
rect 21364 9868 21416 9920
rect 23940 9936 23992 9988
rect 22836 9868 22888 9920
rect 22928 9868 22980 9920
rect 24308 9868 24360 9920
rect 24492 9936 24544 9988
rect 25136 9936 25188 9988
rect 26148 9936 26200 9988
rect 25964 9868 26016 9920
rect 27252 10004 27304 10056
rect 28080 10115 28132 10124
rect 28080 10081 28089 10115
rect 28089 10081 28123 10115
rect 28123 10081 28132 10115
rect 28080 10072 28132 10081
rect 28908 10208 28960 10260
rect 31300 10251 31352 10260
rect 31300 10217 31309 10251
rect 31309 10217 31343 10251
rect 31343 10217 31352 10251
rect 31300 10208 31352 10217
rect 31392 10208 31444 10260
rect 31944 10208 31996 10260
rect 29368 10004 29420 10056
rect 31116 10004 31168 10056
rect 32220 10047 32272 10056
rect 32220 10013 32229 10047
rect 32229 10013 32263 10047
rect 32263 10013 32272 10047
rect 32220 10004 32272 10013
rect 32772 10047 32824 10056
rect 32772 10013 32781 10047
rect 32781 10013 32815 10047
rect 32815 10013 32824 10047
rect 32772 10004 32824 10013
rect 34060 10004 34112 10056
rect 30104 9936 30156 9988
rect 28540 9911 28592 9920
rect 28540 9877 28549 9911
rect 28549 9877 28583 9911
rect 28583 9877 28592 9911
rect 28540 9868 28592 9877
rect 29276 9911 29328 9920
rect 29276 9877 29285 9911
rect 29285 9877 29319 9911
rect 29319 9877 29328 9911
rect 29276 9868 29328 9877
rect 32220 9911 32272 9920
rect 32220 9877 32229 9911
rect 32229 9877 32263 9911
rect 32263 9877 32272 9911
rect 32220 9868 32272 9877
rect 32772 9868 32824 9920
rect 34520 9911 34572 9920
rect 34520 9877 34529 9911
rect 34529 9877 34563 9911
rect 34563 9877 34572 9911
rect 34520 9868 34572 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2872 9664 2924 9716
rect 3240 9707 3292 9716
rect 3240 9673 3249 9707
rect 3249 9673 3283 9707
rect 3283 9673 3292 9707
rect 3240 9664 3292 9673
rect 17224 9664 17276 9716
rect 22928 9664 22980 9716
rect 23020 9664 23072 9716
rect 24032 9707 24084 9716
rect 24032 9673 24041 9707
rect 24041 9673 24075 9707
rect 24075 9673 24084 9707
rect 24032 9664 24084 9673
rect 24124 9664 24176 9716
rect 18604 9596 18656 9648
rect 22100 9596 22152 9648
rect 22192 9528 22244 9580
rect 22468 9596 22520 9648
rect 23296 9596 23348 9648
rect 24308 9596 24360 9648
rect 26240 9664 26292 9716
rect 26608 9664 26660 9716
rect 28080 9664 28132 9716
rect 27160 9596 27212 9648
rect 23020 9528 23072 9580
rect 23940 9528 23992 9580
rect 24032 9528 24084 9580
rect 28540 9596 28592 9648
rect 29276 9596 29328 9648
rect 27528 9571 27580 9580
rect 27528 9537 27537 9571
rect 27537 9537 27571 9571
rect 27571 9537 27580 9571
rect 27528 9528 27580 9537
rect 31300 9528 31352 9580
rect 32772 9571 32824 9580
rect 32772 9537 32781 9571
rect 32781 9537 32815 9571
rect 32815 9537 32824 9571
rect 32772 9528 32824 9537
rect 34520 9528 34572 9580
rect 34796 9528 34848 9580
rect 29368 9460 29420 9512
rect 31116 9460 31168 9512
rect 32220 9503 32272 9512
rect 32220 9469 32229 9503
rect 32229 9469 32263 9503
rect 32263 9469 32272 9503
rect 32220 9460 32272 9469
rect 23756 9324 23808 9376
rect 32588 9367 32640 9376
rect 32588 9333 32597 9367
rect 32597 9333 32631 9367
rect 32631 9333 32640 9367
rect 32588 9324 32640 9333
rect 32956 9367 33008 9376
rect 32956 9333 32965 9367
rect 32965 9333 32999 9367
rect 32999 9333 33008 9367
rect 32956 9324 33008 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 1676 9120 1728 9172
rect 23020 9163 23072 9172
rect 23020 9129 23029 9163
rect 23029 9129 23063 9163
rect 23063 9129 23072 9163
rect 23020 9120 23072 9129
rect 23940 9120 23992 9172
rect 32956 9120 33008 9172
rect 10048 9052 10100 9104
rect 940 8916 992 8968
rect 23756 8916 23808 8968
rect 25044 8959 25096 8968
rect 25044 8925 25053 8959
rect 25053 8925 25087 8959
rect 25087 8925 25096 8959
rect 25044 8916 25096 8925
rect 26240 8916 26292 8968
rect 25964 8848 26016 8900
rect 34060 8916 34112 8968
rect 33048 8823 33100 8832
rect 33048 8789 33057 8823
rect 33057 8789 33091 8823
rect 33091 8789 33100 8823
rect 33048 8780 33100 8789
rect 33508 8823 33560 8832
rect 33508 8789 33517 8823
rect 33517 8789 33551 8823
rect 33551 8789 33560 8823
rect 33508 8780 33560 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 32588 8576 32640 8628
rect 26240 8508 26292 8560
rect 27804 8483 27856 8492
rect 27804 8449 27813 8483
rect 27813 8449 27847 8483
rect 27847 8449 27856 8483
rect 27804 8440 27856 8449
rect 32680 8508 32732 8560
rect 34060 8576 34112 8628
rect 33508 8508 33560 8560
rect 34244 8347 34296 8356
rect 34244 8313 34253 8347
rect 34253 8313 34287 8347
rect 34287 8313 34296 8347
rect 34244 8304 34296 8313
rect 34428 8279 34480 8288
rect 34428 8245 34437 8279
rect 34437 8245 34471 8279
rect 34471 8245 34480 8279
rect 34428 8236 34480 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 32680 8075 32732 8084
rect 32680 8041 32689 8075
rect 32689 8041 32723 8075
rect 32723 8041 32732 8075
rect 32680 8032 32732 8041
rect 33048 7939 33100 7948
rect 33048 7905 33057 7939
rect 33057 7905 33091 7939
rect 33091 7905 33100 7939
rect 33048 7896 33100 7905
rect 34428 7828 34480 7880
rect 34520 7735 34572 7744
rect 34520 7701 34529 7735
rect 34529 7701 34563 7735
rect 34563 7701 34572 7735
rect 34520 7692 34572 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 34612 7352 34664 7404
rect 34796 7352 34848 7404
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 940 6740 992 6792
rect 1492 6604 1544 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 34336 5695 34388 5704
rect 34336 5661 34345 5695
rect 34345 5661 34379 5695
rect 34379 5661 34388 5695
rect 34336 5652 34388 5661
rect 34060 5584 34112 5636
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2964 4768 3016 4820
rect 940 4564 992 4616
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 34520 3476 34572 3528
rect 34612 3408 34664 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1400 2592 1452 2644
rect 27804 2592 27856 2644
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 940 2388 992 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 952 36174 980 36751
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 940 36168 992 36174
rect 940 36110 992 36116
rect 33140 36168 33192 36174
rect 33140 36110 33192 36116
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 35894 1624 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 1596 35866 1716 35894
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 940 35080 992 35086
rect 940 35022 992 35028
rect 952 34649 980 35022
rect 938 34640 994 34649
rect 938 34575 994 34584
rect 940 32904 992 32910
rect 940 32846 992 32852
rect 952 32473 980 32846
rect 938 32464 994 32473
rect 938 32399 994 32408
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30297 1440 30670
rect 1398 30288 1454 30297
rect 1398 30223 1454 30232
rect 940 28552 992 28558
rect 940 28494 992 28500
rect 952 28121 980 28494
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 938 28112 994 28121
rect 938 28047 994 28056
rect 1596 25974 1624 28358
rect 1688 26450 1716 35866
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 1860 34944 1912 34950
rect 1860 34886 1912 34892
rect 1676 26444 1728 26450
rect 1676 26386 1728 26392
rect 1584 25968 1636 25974
rect 938 25936 994 25945
rect 1584 25910 1636 25916
rect 938 25871 940 25880
rect 992 25871 994 25880
rect 940 25842 992 25848
rect 1768 25696 1820 25702
rect 1768 25638 1820 25644
rect 940 24812 992 24818
rect 940 24754 992 24760
rect 952 23769 980 24754
rect 1584 24608 1636 24614
rect 1584 24550 1636 24556
rect 1400 24268 1452 24274
rect 1400 24210 1452 24216
rect 938 23760 994 23769
rect 938 23695 994 23704
rect 1412 23662 1440 24210
rect 1596 23866 1624 24550
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1780 22710 1808 25638
rect 1872 24274 1900 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 2872 30592 2924 30598
rect 2872 30534 2924 30540
rect 2884 27674 2912 30534
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 3608 27328 3660 27334
rect 3608 27270 3660 27276
rect 3620 26790 3648 27270
rect 3608 26784 3660 26790
rect 3608 26726 3660 26732
rect 3620 26450 3648 26726
rect 3608 26444 3660 26450
rect 3608 26386 3660 26392
rect 4080 26314 4108 32710
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19904 28614 20116 28642
rect 19904 28422 19932 28614
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19996 28422 20024 28494
rect 19340 28416 19392 28422
rect 19340 28358 19392 28364
rect 19892 28416 19944 28422
rect 19892 28358 19944 28364
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 19352 28082 19380 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19340 28076 19392 28082
rect 19340 28018 19392 28024
rect 19432 28008 19484 28014
rect 19432 27950 19484 27956
rect 19524 28008 19576 28014
rect 19524 27950 19576 27956
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 14924 27532 14976 27538
rect 14924 27474 14976 27480
rect 16764 27532 16816 27538
rect 16764 27474 16816 27480
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 4160 27396 4212 27402
rect 4160 27338 4212 27344
rect 4172 27130 4200 27338
rect 5540 27328 5592 27334
rect 5540 27270 5592 27276
rect 5816 27328 5868 27334
rect 5816 27270 5868 27276
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 5552 26738 5580 27270
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 2136 26308 2188 26314
rect 2136 26250 2188 26256
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 4068 26308 4120 26314
rect 4068 26250 4120 26256
rect 4712 26308 4764 26314
rect 4712 26250 4764 26256
rect 2044 26240 2096 26246
rect 2044 26182 2096 26188
rect 2056 25838 2084 26182
rect 2148 26042 2176 26250
rect 2136 26036 2188 26042
rect 2136 25978 2188 25984
rect 2044 25832 2096 25838
rect 2044 25774 2096 25780
rect 2056 24410 2084 25774
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2884 25158 2912 25638
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 3608 25152 3660 25158
rect 3608 25094 3660 25100
rect 2044 24404 2096 24410
rect 2044 24346 2096 24352
rect 1860 24268 1912 24274
rect 1860 24210 1912 24216
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2792 23322 2820 23666
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2884 23118 2912 25094
rect 3620 24614 3648 25094
rect 3988 24886 4016 26250
rect 4724 26042 4752 26250
rect 4712 26036 4764 26042
rect 4712 25978 4764 25984
rect 4620 25764 4672 25770
rect 4620 25706 4672 25712
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4160 25152 4212 25158
rect 4160 25094 4212 25100
rect 3976 24880 4028 24886
rect 4172 24834 4200 25094
rect 3976 24822 4028 24828
rect 4080 24818 4200 24834
rect 4632 24818 4660 25706
rect 4068 24812 4200 24818
rect 4120 24806 4200 24812
rect 4252 24812 4304 24818
rect 4068 24754 4120 24760
rect 4252 24754 4304 24760
rect 4620 24812 4672 24818
rect 4620 24754 4672 24760
rect 4264 24698 4292 24754
rect 4080 24670 4292 24698
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3620 24410 3648 24550
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 3620 23526 3648 24346
rect 4080 24290 4108 24670
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4632 24410 4660 24754
rect 4712 24608 4764 24614
rect 4712 24550 4764 24556
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4724 24290 4752 24550
rect 4080 24262 4200 24290
rect 4172 24206 4200 24262
rect 4632 24262 4752 24290
rect 4160 24200 4212 24206
rect 4160 24142 4212 24148
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4080 23866 4108 24006
rect 3792 23860 3844 23866
rect 3792 23802 3844 23808
rect 4068 23860 4120 23866
rect 4068 23802 4120 23808
rect 3608 23520 3660 23526
rect 3608 23462 3660 23468
rect 2872 23112 2924 23118
rect 2872 23054 2924 23060
rect 3620 22982 3648 23462
rect 3424 22976 3476 22982
rect 3424 22918 3476 22924
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 1768 22704 1820 22710
rect 1768 22646 1820 22652
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 2320 22432 2372 22438
rect 2320 22374 2372 22380
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21593 980 21966
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1596 21690 1624 21830
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 938 21584 994 21593
rect 2332 21554 2360 22374
rect 2884 22234 2912 22646
rect 2872 22228 2924 22234
rect 2872 22170 2924 22176
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 938 21519 994 21528
rect 2320 21548 2372 21554
rect 2320 21490 2372 21496
rect 3160 21146 3188 22034
rect 3332 21616 3384 21622
rect 3332 21558 3384 21564
rect 3344 21146 3372 21558
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3332 21140 3384 21146
rect 3332 21082 3384 21088
rect 3240 20936 3292 20942
rect 3240 20878 3292 20884
rect 940 19848 992 19854
rect 940 19790 992 19796
rect 952 19417 980 19790
rect 1584 19712 1636 19718
rect 1584 19654 1636 19660
rect 938 19408 994 19417
rect 938 19343 994 19352
rect 1596 18358 1624 19654
rect 1584 18352 1636 18358
rect 1584 18294 1636 18300
rect 1400 18216 1452 18222
rect 1400 18158 1452 18164
rect 940 17672 992 17678
rect 940 17614 992 17620
rect 952 17241 980 17614
rect 938 17232 994 17241
rect 938 17167 994 17176
rect 1412 16590 1440 18158
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3160 17678 3188 18022
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1688 16658 1716 17478
rect 3252 17338 3280 20878
rect 3436 18290 3464 22918
rect 3804 22098 3832 23802
rect 4172 23610 4200 24142
rect 4632 24070 4660 24262
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4080 23594 4200 23610
rect 4068 23588 4200 23594
rect 4120 23582 4200 23588
rect 4068 23530 4120 23536
rect 4080 23202 4108 23530
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4080 23174 4200 23202
rect 4172 23118 4200 23174
rect 4344 23180 4396 23186
rect 4344 23122 4396 23128
rect 4160 23112 4212 23118
rect 4160 23054 4212 23060
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 3976 22568 4028 22574
rect 3976 22510 4028 22516
rect 3988 22234 4016 22510
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3792 22092 3844 22098
rect 4080 22094 4108 22918
rect 4356 22778 4384 23122
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4632 22642 4660 24006
rect 4908 23322 4936 24142
rect 5000 23866 5028 26726
rect 5552 26710 5764 26738
rect 5540 26240 5592 26246
rect 5540 26182 5592 26188
rect 5552 25430 5580 26182
rect 5540 25424 5592 25430
rect 5540 25366 5592 25372
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 5092 24206 5120 25094
rect 5552 24818 5580 25366
rect 5632 25152 5684 25158
rect 5632 25094 5684 25100
rect 5356 24812 5408 24818
rect 5356 24754 5408 24760
rect 5540 24812 5592 24818
rect 5540 24754 5592 24760
rect 5368 24410 5396 24754
rect 5356 24404 5408 24410
rect 5356 24346 5408 24352
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 5092 24070 5120 24142
rect 5080 24064 5132 24070
rect 5080 24006 5132 24012
rect 4988 23860 5040 23866
rect 4988 23802 5040 23808
rect 5092 23526 5120 24006
rect 5080 23520 5132 23526
rect 5080 23462 5132 23468
rect 4896 23316 4948 23322
rect 4896 23258 4948 23264
rect 4620 22636 4672 22642
rect 4620 22578 4672 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4528 22228 4580 22234
rect 4528 22170 4580 22176
rect 3792 22034 3844 22040
rect 3988 22066 4108 22094
rect 3988 21894 4016 22066
rect 3976 21888 4028 21894
rect 3976 21830 4028 21836
rect 3988 21486 4016 21830
rect 4436 21548 4488 21554
rect 4540 21536 4568 22170
rect 4632 22094 4660 22578
rect 4712 22500 4764 22506
rect 4712 22442 4764 22448
rect 4724 22234 4752 22442
rect 4712 22228 4764 22234
rect 4712 22170 4764 22176
rect 4632 22066 4752 22094
rect 4620 21548 4672 21554
rect 4540 21508 4620 21536
rect 4436 21490 4488 21496
rect 4620 21490 4672 21496
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 4448 21350 4476 21490
rect 4436 21344 4488 21350
rect 4436 21286 4488 21292
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3700 18080 3752 18086
rect 3700 18022 3752 18028
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 3240 17332 3292 17338
rect 3240 17274 3292 17280
rect 3252 16794 3280 17274
rect 3620 17202 3648 17682
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 1676 16652 1728 16658
rect 1676 16594 1728 16600
rect 1400 16584 1452 16590
rect 1400 16526 1452 16532
rect 1412 15910 1440 16526
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 1400 15904 1452 15910
rect 1400 15846 1452 15852
rect 1412 15638 1440 15846
rect 1400 15632 1452 15638
rect 1452 15580 1532 15586
rect 1400 15574 1532 15580
rect 1412 15558 1532 15574
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15201 1440 15438
rect 1398 15192 1454 15201
rect 1504 15162 1532 15558
rect 1398 15127 1454 15136
rect 1492 15156 1544 15162
rect 1492 15098 1544 15104
rect 1504 14498 1532 15098
rect 1584 15088 1636 15094
rect 1584 15030 1636 15036
rect 2320 15088 2372 15094
rect 2320 15030 2372 15036
rect 1412 14482 1532 14498
rect 1412 14476 1544 14482
rect 1412 14470 1492 14476
rect 1412 13394 1440 14470
rect 1492 14418 1544 14424
rect 1492 14340 1544 14346
rect 1492 14282 1544 14288
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 938 12880 994 12889
rect 938 12815 940 12824
rect 992 12815 994 12824
rect 940 12786 992 12792
rect 1412 12306 1440 13330
rect 1400 12300 1452 12306
rect 1400 12242 1452 12248
rect 1412 11762 1440 12242
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1400 9988 1452 9994
rect 1400 9930 1452 9936
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 952 8537 980 8910
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 952 6361 980 6734
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1412 2650 1440 9930
rect 1504 6662 1532 14282
rect 1596 11354 1624 15030
rect 2332 14074 2360 15030
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 2320 14068 2372 14074
rect 2320 14010 2372 14016
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 2412 13252 2464 13258
rect 2412 13194 2464 13200
rect 1688 12986 1716 13194
rect 2424 12986 2452 13194
rect 2884 12986 2912 14418
rect 3160 13938 3188 16390
rect 3252 14618 3280 16730
rect 3620 16250 3648 17138
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3620 15706 3648 16186
rect 3608 15700 3660 15706
rect 3608 15642 3660 15648
rect 3712 15570 3740 18022
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4724 17882 4752 22066
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4816 21690 4844 21830
rect 4804 21684 4856 21690
rect 4804 21626 4856 21632
rect 4816 20806 4844 21626
rect 4908 21350 4936 23258
rect 5092 23050 5120 23462
rect 5080 23044 5132 23050
rect 5080 22986 5132 22992
rect 5172 23044 5224 23050
rect 5172 22986 5224 22992
rect 5092 22574 5120 22986
rect 5184 22778 5212 22986
rect 5264 22976 5316 22982
rect 5264 22918 5316 22924
rect 5172 22772 5224 22778
rect 5172 22714 5224 22720
rect 5276 22642 5304 22918
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5092 22438 5120 22510
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 5172 22432 5224 22438
rect 5172 22374 5224 22380
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 21486 5028 21830
rect 4988 21480 5040 21486
rect 4988 21422 5040 21428
rect 4896 21344 4948 21350
rect 4896 21286 4948 21292
rect 5000 20942 5028 21422
rect 5092 21146 5120 22374
rect 5184 22114 5212 22374
rect 5276 22234 5304 22578
rect 5368 22506 5396 24346
rect 5644 24206 5672 25094
rect 5736 24834 5764 26710
rect 5828 26586 5856 27270
rect 14844 26586 14872 27406
rect 14936 26994 14964 27474
rect 15108 27464 15160 27470
rect 15160 27412 15332 27418
rect 15108 27406 15332 27412
rect 15120 27390 15332 27406
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 5816 26580 5868 26586
rect 5816 26522 5868 26528
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 5828 25378 5856 26522
rect 9312 26444 9364 26450
rect 9312 26386 9364 26392
rect 9772 26444 9824 26450
rect 9772 26386 9824 26392
rect 12992 26444 13044 26450
rect 12992 26386 13044 26392
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 6840 26042 6868 26318
rect 9324 26314 9352 26386
rect 8300 26308 8352 26314
rect 8300 26250 8352 26256
rect 9312 26308 9364 26314
rect 9312 26250 9364 26256
rect 9680 26308 9732 26314
rect 9680 26250 9732 26256
rect 6828 26036 6880 26042
rect 6828 25978 6880 25984
rect 5908 25900 5960 25906
rect 5908 25842 5960 25848
rect 5920 25498 5948 25842
rect 6000 25832 6052 25838
rect 6000 25774 6052 25780
rect 5908 25492 5960 25498
rect 5908 25434 5960 25440
rect 5828 25350 5948 25378
rect 5736 24806 5856 24834
rect 5920 24818 5948 25350
rect 6012 24886 6040 25774
rect 8312 25498 8340 26250
rect 9692 26042 9720 26250
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9784 25922 9812 26386
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 9600 25894 9812 25922
rect 8300 25492 8352 25498
rect 8300 25434 8352 25440
rect 6000 24880 6052 24886
rect 6000 24822 6052 24828
rect 8312 24818 8340 25434
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 5724 24744 5776 24750
rect 5724 24686 5776 24692
rect 5736 24410 5764 24686
rect 5724 24404 5776 24410
rect 5724 24346 5776 24352
rect 5632 24200 5684 24206
rect 5632 24142 5684 24148
rect 5828 23338 5856 24806
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 8300 24812 8352 24818
rect 8300 24754 8352 24760
rect 7944 24410 7972 24754
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 8312 23798 8340 24754
rect 9416 24410 9444 24822
rect 9600 24410 9628 25894
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9404 24404 9456 24410
rect 9404 24346 9456 24352
rect 9588 24404 9640 24410
rect 9588 24346 9640 24352
rect 9876 24070 9904 25638
rect 10704 25498 10732 26250
rect 12912 25906 12940 26318
rect 13004 25974 13032 26386
rect 14936 26382 14964 26930
rect 15304 26790 15332 27390
rect 15660 27328 15712 27334
rect 15660 27270 15712 27276
rect 15936 27328 15988 27334
rect 15936 27270 15988 27276
rect 15672 27130 15700 27270
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15948 27062 15976 27270
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 16304 26988 16356 26994
rect 16304 26930 16356 26936
rect 15844 26852 15896 26858
rect 15844 26794 15896 26800
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15384 26784 15436 26790
rect 15384 26726 15436 26732
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 14924 26376 14976 26382
rect 14924 26318 14976 26324
rect 13268 26240 13320 26246
rect 13268 26182 13320 26188
rect 12992 25968 13044 25974
rect 12992 25910 13044 25916
rect 12900 25900 12952 25906
rect 12900 25842 12952 25848
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10704 24886 10732 25434
rect 12912 25362 12940 25842
rect 13004 25362 13032 25910
rect 13280 25838 13308 26182
rect 13648 26042 13676 26318
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13268 25832 13320 25838
rect 13268 25774 13320 25780
rect 14648 25696 14700 25702
rect 14648 25638 14700 25644
rect 11244 25356 11296 25362
rect 11244 25298 11296 25304
rect 12900 25356 12952 25362
rect 12900 25298 12952 25304
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 11152 25288 11204 25294
rect 11152 25230 11204 25236
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 10692 24880 10744 24886
rect 10692 24822 10744 24828
rect 11072 24800 11100 25162
rect 11164 24954 11192 25230
rect 11256 24954 11284 25298
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 12452 24954 12480 25230
rect 12532 25220 12584 25226
rect 12532 25162 12584 25168
rect 12544 24954 12572 25162
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 11244 24948 11296 24954
rect 11244 24890 11296 24896
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 11152 24812 11204 24818
rect 11072 24772 11152 24800
rect 11152 24754 11204 24760
rect 11428 24812 11480 24818
rect 11428 24754 11480 24760
rect 11704 24812 11756 24818
rect 11704 24754 11756 24760
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12348 24812 12400 24818
rect 12348 24754 12400 24760
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 10152 24410 10180 24550
rect 10140 24404 10192 24410
rect 10140 24346 10192 24352
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 8852 23792 8904 23798
rect 8852 23734 8904 23740
rect 6368 23724 6420 23730
rect 6368 23666 6420 23672
rect 5644 23310 5856 23338
rect 6380 23322 6408 23666
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 6368 23316 6420 23322
rect 5644 23118 5672 23310
rect 6368 23258 6420 23264
rect 7024 23186 7052 23462
rect 5724 23180 5776 23186
rect 5724 23122 5776 23128
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 5632 23112 5684 23118
rect 5632 23054 5684 23060
rect 5644 22778 5672 23054
rect 5736 22778 5764 23122
rect 8772 23118 8800 23462
rect 8864 23118 8892 23734
rect 9036 23724 9088 23730
rect 9036 23666 9088 23672
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 9048 23322 9076 23666
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 6368 23112 6420 23118
rect 6368 23054 6420 23060
rect 8760 23112 8812 23118
rect 8760 23054 8812 23060
rect 8852 23112 8904 23118
rect 8852 23054 8904 23060
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5724 22772 5776 22778
rect 5724 22714 5776 22720
rect 5356 22500 5408 22506
rect 5356 22442 5408 22448
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5356 22160 5408 22166
rect 5184 22086 5304 22114
rect 5356 22102 5408 22108
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5184 21146 5212 21286
rect 5080 21140 5132 21146
rect 5080 21082 5132 21088
rect 5172 21140 5224 21146
rect 5172 21082 5224 21088
rect 4988 20936 5040 20942
rect 4988 20878 5040 20884
rect 4804 20800 4856 20806
rect 4804 20742 4856 20748
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3896 17202 3924 17614
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3884 17196 3936 17202
rect 3884 17138 3936 17144
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3804 16794 3832 17070
rect 3792 16788 3844 16794
rect 3792 16730 3844 16736
rect 3988 16726 4016 17478
rect 3976 16720 4028 16726
rect 3976 16662 4028 16668
rect 3792 16176 3844 16182
rect 3792 16118 3844 16124
rect 3700 15564 3752 15570
rect 3700 15506 3752 15512
rect 3608 15360 3660 15366
rect 3608 15302 3660 15308
rect 3332 14816 3384 14822
rect 3332 14758 3384 14764
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3148 13932 3200 13938
rect 3148 13874 3200 13880
rect 3240 13728 3292 13734
rect 3344 13716 3372 14758
rect 3620 14618 3648 15302
rect 3804 15162 3832 16118
rect 3884 15564 3936 15570
rect 3884 15506 3936 15512
rect 3792 15156 3844 15162
rect 3792 15098 3844 15104
rect 3804 14618 3832 15098
rect 3896 14822 3924 15506
rect 3988 15366 4016 16662
rect 4080 16658 4108 17818
rect 4816 17762 4844 20742
rect 4724 17734 4844 17762
rect 5184 17746 5212 21082
rect 5172 17740 5224 17746
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16726 4660 17614
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 15910 4108 16390
rect 4172 16250 4200 16526
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4080 15434 4108 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15706 4660 16662
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3792 14612 3844 14618
rect 3792 14554 3844 14560
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3292 13688 3372 13716
rect 3240 13670 3292 13676
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 2412 12980 2464 12986
rect 2412 12922 2464 12928
rect 2872 12980 2924 12986
rect 2872 12922 2924 12928
rect 3160 12850 3188 13126
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 1676 12164 1728 12170
rect 1676 12106 1728 12112
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1688 9178 1716 12106
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 1676 9172 1728 9178
rect 1676 9114 1728 9120
rect 2792 6914 2820 11630
rect 3252 10674 3280 13670
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3332 12980 3384 12986
rect 3332 12922 3384 12928
rect 3344 12374 3372 12922
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2884 9722 2912 9930
rect 3252 9722 3280 10610
rect 3620 10062 3648 13194
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3896 12986 3924 13126
rect 3884 12980 3936 12986
rect 3884 12922 3936 12928
rect 3988 12918 4016 13874
rect 4080 13734 4108 15370
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13258 4108 13670
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 13806
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4068 13252 4120 13258
rect 4068 13194 4120 13200
rect 3976 12912 4028 12918
rect 3976 12854 4028 12860
rect 4264 12850 4292 13262
rect 4252 12844 4304 12850
rect 4252 12786 4304 12792
rect 4356 12646 4384 13262
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 4632 12850 4660 13194
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4344 12640 4396 12646
rect 4344 12582 4396 12588
rect 4080 12442 4108 12582
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4632 12238 4660 12786
rect 4724 12714 4752 17734
rect 5172 17682 5224 17688
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5092 16794 5120 17070
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 15502 5028 16526
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4988 15360 5040 15366
rect 4988 15302 5040 15308
rect 4816 15162 4844 15302
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 5000 14958 5028 15302
rect 4988 14952 5040 14958
rect 5184 14940 5212 17682
rect 5276 17678 5304 22086
rect 5368 21554 5396 22102
rect 5356 21548 5408 21554
rect 5356 21490 5408 21496
rect 5828 21146 5856 23054
rect 6380 22574 6408 23054
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22642 8432 22918
rect 8392 22636 8444 22642
rect 8392 22578 8444 22584
rect 6368 22568 6420 22574
rect 6368 22510 6420 22516
rect 6380 21894 6408 22510
rect 8300 21956 8352 21962
rect 8300 21898 8352 21904
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 6380 21486 6408 21830
rect 7380 21616 7432 21622
rect 7380 21558 7432 21564
rect 6368 21480 6420 21486
rect 6368 21422 6420 21428
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 6000 21004 6052 21010
rect 6000 20946 6052 20952
rect 6012 20534 6040 20946
rect 6092 20868 6144 20874
rect 6092 20810 6144 20816
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 6104 17678 6132 20810
rect 6380 20466 6408 21422
rect 7392 21146 7420 21558
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7564 20800 7616 20806
rect 7564 20742 7616 20748
rect 7380 20528 7432 20534
rect 7380 20470 7432 20476
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6380 18426 6408 20402
rect 7392 20058 7420 20470
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 7576 19718 7604 20742
rect 8312 20058 8340 21898
rect 8404 21894 8432 22578
rect 8864 22506 8892 23054
rect 9784 22574 9812 23666
rect 9876 23526 9904 24006
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 9956 23044 10008 23050
rect 9956 22986 10008 22992
rect 9968 22778 9996 22986
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9772 22568 9824 22574
rect 9772 22510 9824 22516
rect 8852 22500 8904 22506
rect 8852 22442 8904 22448
rect 8864 22234 8892 22442
rect 8852 22228 8904 22234
rect 8852 22170 8904 22176
rect 8392 21888 8444 21894
rect 8392 21830 8444 21836
rect 9404 21888 9456 21894
rect 9404 21830 9456 21836
rect 8404 20942 8432 21830
rect 9416 21350 9444 21830
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 8392 20936 8444 20942
rect 8392 20878 8444 20884
rect 9416 20874 9444 21286
rect 9692 21078 9720 21490
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9404 20868 9456 20874
rect 9404 20810 9456 20816
rect 8300 20052 8352 20058
rect 8300 19994 8352 20000
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 6368 18420 6420 18426
rect 6368 18362 6420 18368
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 6092 17672 6144 17678
rect 6092 17614 6144 17620
rect 6380 17202 6408 18362
rect 6460 17536 6512 17542
rect 6460 17478 6512 17484
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6472 17338 6500 17478
rect 6460 17332 6512 17338
rect 6460 17274 6512 17280
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 5540 16720 5592 16726
rect 5540 16662 5592 16668
rect 5264 16516 5316 16522
rect 5264 16458 5316 16464
rect 5276 15026 5304 16458
rect 5552 16182 5580 16662
rect 6472 16658 6500 16934
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6748 16454 6776 17478
rect 7576 17270 7604 19654
rect 9220 19168 9272 19174
rect 9220 19110 9272 19116
rect 9232 18290 9260 19110
rect 9220 18284 9272 18290
rect 9220 18226 9272 18232
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7576 17134 7604 17206
rect 9232 17202 9260 17478
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 8760 17128 8812 17134
rect 8760 17070 8812 17076
rect 6840 16794 6868 17070
rect 7012 16992 7064 16998
rect 7012 16934 7064 16940
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 7024 16522 7052 16934
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 5540 16176 5592 16182
rect 5540 16118 5592 16124
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6380 15162 6408 16050
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6932 15094 6960 15846
rect 8680 15706 8708 16730
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 4988 14894 5040 14900
rect 5092 14912 5212 14940
rect 5092 14804 5120 14912
rect 4816 14776 5120 14804
rect 5172 14816 5224 14822
rect 4816 13462 4844 14776
rect 5172 14758 5224 14764
rect 5184 14618 5212 14758
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 7484 14414 7512 15302
rect 8312 15094 8340 15302
rect 8300 15088 8352 15094
rect 8300 15030 8352 15036
rect 8680 15026 8708 15642
rect 8772 15366 8800 17070
rect 9416 16658 9444 20810
rect 9588 20800 9640 20806
rect 9588 20742 9640 20748
rect 9600 20330 9628 20742
rect 9692 20602 9720 21014
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9588 20324 9640 20330
rect 9588 20266 9640 20272
rect 9784 19514 9812 22510
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10508 21344 10560 21350
rect 10508 21286 10560 21292
rect 10428 21146 10456 21286
rect 10520 21146 10548 21286
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 10508 21140 10560 21146
rect 10508 21082 10560 21088
rect 10428 20466 10456 21082
rect 10416 20460 10468 20466
rect 10416 20402 10468 20408
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10060 19514 10088 20334
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 10048 19508 10100 19514
rect 10048 19450 10100 19456
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9692 18766 9720 19178
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9692 18426 9720 18702
rect 9876 18630 9904 19314
rect 10324 18760 10376 18766
rect 10324 18702 10376 18708
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9600 16998 9628 18226
rect 9692 17882 9720 18362
rect 9876 18086 9904 18566
rect 10336 18426 10364 18702
rect 10324 18420 10376 18426
rect 10324 18362 10376 18368
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9876 17542 9904 18022
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8312 14618 8340 14894
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 6184 14408 6236 14414
rect 6184 14350 6236 14356
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 6196 13938 6224 14350
rect 8680 14074 8708 14962
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 6184 13932 6236 13938
rect 6184 13874 6236 13880
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4908 13462 4936 13670
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4896 13456 4948 13462
rect 4896 13398 4948 13404
rect 4816 13172 4844 13398
rect 8680 13326 8708 14010
rect 8772 13938 8800 15302
rect 9600 14482 9628 16934
rect 9876 16794 9904 17478
rect 9864 16788 9916 16794
rect 9864 16730 9916 16736
rect 9876 15094 9904 16730
rect 9864 15088 9916 15094
rect 9864 15030 9916 15036
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 10508 14272 10560 14278
rect 10508 14214 10560 14220
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13734 8800 13874
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 5172 13320 5224 13326
rect 5172 13262 5224 13268
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 8668 13320 8720 13326
rect 8668 13262 8720 13268
rect 5092 13172 5120 13262
rect 4816 13144 5120 13172
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 5092 12646 5120 13144
rect 5184 12918 5212 13262
rect 5276 13190 5304 13262
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5276 12850 5304 13126
rect 5368 12986 5396 13262
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 8392 12912 8444 12918
rect 8392 12854 8444 12860
rect 5264 12844 5316 12850
rect 5264 12786 5316 12792
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 8404 12442 8432 12854
rect 8772 12442 8800 13670
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8956 12986 8984 13262
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9692 12986 9720 13194
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 8956 12850 8984 12922
rect 10520 12918 10548 14214
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 8392 12436 8444 12442
rect 8392 12378 8444 12384
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11762 3924 12038
rect 4632 11898 4660 12174
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7208 11898 7236 12038
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4632 10266 4660 11630
rect 9600 11626 9628 12718
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 12442 10088 12582
rect 10048 12436 10100 12442
rect 10048 12378 10100 12384
rect 10060 11762 10088 12378
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9588 11620 9640 11626
rect 9588 11562 9640 11568
rect 9600 11082 9628 11562
rect 10060 11558 10088 11698
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 4620 10260 4672 10266
rect 4620 10202 4672 10208
rect 3608 10056 3660 10062
rect 3608 9998 3660 10004
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2792 6886 3004 6914
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 2976 4826 3004 6886
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1400 2644 1452 2650
rect 1400 2586 1452 2592
rect 9600 2514 9628 11018
rect 10060 9110 10088 11494
rect 10612 10810 10640 23462
rect 11164 22642 11192 24754
rect 11440 24070 11468 24754
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23866 11468 24006
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11716 23594 11744 24754
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11704 23588 11756 23594
rect 11704 23530 11756 23536
rect 11992 23526 12020 24550
rect 12176 24206 12204 24754
rect 12164 24200 12216 24206
rect 12164 24142 12216 24148
rect 12360 23730 12388 24754
rect 12452 23798 12480 24754
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13556 24138 13584 24550
rect 14108 24206 14136 24550
rect 14200 24206 14228 24754
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 14096 24200 14148 24206
rect 14188 24200 14240 24206
rect 14096 24142 14148 24148
rect 14186 24168 14188 24177
rect 14280 24200 14332 24206
rect 14240 24168 14242 24177
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12622 24032 12678 24041
rect 12440 23792 12492 23798
rect 12440 23734 12492 23740
rect 12348 23724 12400 23730
rect 12348 23666 12400 23672
rect 11244 23520 11296 23526
rect 11244 23462 11296 23468
rect 11980 23520 12032 23526
rect 11980 23462 12032 23468
rect 11256 23118 11284 23462
rect 11992 23322 12020 23462
rect 11980 23316 12032 23322
rect 11980 23258 12032 23264
rect 11244 23112 11296 23118
rect 11244 23054 11296 23060
rect 11888 23044 11940 23050
rect 11992 23032 12020 23258
rect 11940 23004 12020 23032
rect 12348 23044 12400 23050
rect 11888 22986 11940 22992
rect 12348 22986 12400 22992
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11164 21690 11192 22578
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11624 21690 11652 21830
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11244 21616 11296 21622
rect 11244 21558 11296 21564
rect 10784 21480 10836 21486
rect 10784 21422 10836 21428
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10796 20942 10824 21422
rect 10876 21072 10928 21078
rect 10876 21014 10928 21020
rect 10692 20936 10744 20942
rect 10692 20878 10744 20884
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10704 20398 10732 20878
rect 10692 20392 10744 20398
rect 10692 20334 10744 20340
rect 10796 19990 10824 20878
rect 10888 20806 10916 21014
rect 10980 20942 11008 21422
rect 11256 20942 11284 21558
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 10968 20936 11020 20942
rect 10968 20878 11020 20884
rect 11152 20936 11204 20942
rect 11152 20878 11204 20884
rect 11244 20936 11296 20942
rect 11244 20878 11296 20884
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10888 20602 10916 20742
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10784 19984 10836 19990
rect 10784 19926 10836 19932
rect 10796 18426 10824 19926
rect 10980 19310 11008 20742
rect 11164 20602 11192 20878
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 11152 20596 11204 20602
rect 11152 20538 11204 20544
rect 11072 20058 11100 20538
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11072 19922 11100 19994
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10968 19304 11020 19310
rect 10968 19246 11020 19252
rect 10980 18698 11008 19246
rect 11152 19168 11204 19174
rect 11440 19156 11468 20810
rect 11532 19310 11560 21490
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11808 20942 11836 21286
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 20466 11744 20742
rect 11612 20460 11664 20466
rect 11612 20402 11664 20408
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11624 19786 11652 20402
rect 11808 19854 11836 20878
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11612 19304 11664 19310
rect 11612 19246 11664 19252
rect 11796 19304 11848 19310
rect 11796 19246 11848 19252
rect 11624 19156 11652 19246
rect 11440 19128 11652 19156
rect 11152 19110 11204 19116
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 11060 18284 11112 18290
rect 11060 18226 11112 18232
rect 11072 17678 11100 18226
rect 11164 18086 11192 19110
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11164 17882 11192 18022
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11532 17814 11560 18770
rect 11624 18426 11652 19128
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11612 18420 11664 18426
rect 11612 18362 11664 18368
rect 11716 18290 11744 18566
rect 11808 18290 11836 19246
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11796 18284 11848 18290
rect 11796 18226 11848 18232
rect 11520 17808 11572 17814
rect 11520 17750 11572 17756
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 10888 17270 10916 17478
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 11532 17202 11560 17750
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11716 16998 11744 18226
rect 11704 16992 11756 16998
rect 11704 16934 11756 16940
rect 10968 16448 11020 16454
rect 10968 16390 11020 16396
rect 10980 16250 11008 16390
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 10980 14618 11008 16186
rect 11900 16182 11928 22986
rect 11978 21720 12034 21729
rect 11978 21655 11980 21664
rect 12032 21655 12034 21664
rect 11980 21626 12032 21632
rect 12360 21486 12388 22986
rect 12544 22642 12572 24006
rect 12622 23967 12678 23976
rect 12636 23594 12664 23967
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12728 23730 12756 23802
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12900 23724 12952 23730
rect 13004 23712 13032 24074
rect 13924 24070 13952 24142
rect 14384 24188 14412 25094
rect 14568 24954 14596 25230
rect 14556 24948 14608 24954
rect 14556 24890 14608 24896
rect 14464 24676 14516 24682
rect 14464 24618 14516 24624
rect 14332 24160 14412 24188
rect 14280 24142 14332 24148
rect 14186 24103 14242 24112
rect 13912 24064 13964 24070
rect 13964 24012 14136 24018
rect 13912 24006 14136 24012
rect 13924 23990 14136 24006
rect 12952 23684 13032 23712
rect 12900 23666 12952 23672
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12728 22982 12756 23666
rect 13004 23118 13032 23684
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13832 23322 13860 23666
rect 14108 23322 14136 23990
rect 14292 23730 14320 24142
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23866 14412 24006
rect 14372 23860 14424 23866
rect 14372 23802 14424 23808
rect 14280 23724 14332 23730
rect 14332 23684 14412 23712
rect 14280 23666 14332 23672
rect 13820 23316 13872 23322
rect 13820 23258 13872 23264
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 12992 23112 13044 23118
rect 12992 23054 13044 23060
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12348 21480 12400 21486
rect 12348 21422 12400 21428
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 12912 20602 12940 20742
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12532 20528 12584 20534
rect 12584 20476 12940 20482
rect 12532 20470 12940 20476
rect 12544 20466 12940 20470
rect 12544 20460 12952 20466
rect 12544 20454 12900 20460
rect 12900 20402 12952 20408
rect 12532 20324 12584 20330
rect 13004 20312 13032 23054
rect 13268 22568 13320 22574
rect 13268 22510 13320 22516
rect 13280 21894 13308 22510
rect 13820 22500 13872 22506
rect 13820 22442 13872 22448
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13280 21690 13308 21830
rect 13268 21684 13320 21690
rect 13268 21626 13320 21632
rect 13452 21684 13504 21690
rect 13452 21626 13504 21632
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13280 20602 13308 21490
rect 13268 20596 13320 20602
rect 13268 20538 13320 20544
rect 13280 20466 13308 20538
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13188 20312 13216 20402
rect 12584 20284 13216 20312
rect 12532 20266 12584 20272
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11992 19514 12020 19790
rect 12084 19514 12112 19926
rect 12624 19712 12676 19718
rect 12346 19680 12402 19689
rect 12624 19654 12676 19660
rect 12346 19615 12402 19624
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 11992 17610 12020 19450
rect 12084 18970 12112 19450
rect 12176 19310 12204 19450
rect 12360 19310 12388 19615
rect 12636 19378 12664 19654
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 12072 18964 12124 18970
rect 12072 18906 12124 18912
rect 12176 18850 12204 19246
rect 12176 18834 12388 18850
rect 12176 18828 12400 18834
rect 12176 18822 12348 18828
rect 12348 18770 12400 18776
rect 12256 18692 12308 18698
rect 12256 18634 12308 18640
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 12084 17746 12112 18226
rect 12268 18222 12296 18634
rect 12348 18624 12400 18630
rect 12348 18566 12400 18572
rect 12360 18290 12388 18566
rect 12452 18426 12480 19314
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12348 18284 12400 18290
rect 12348 18226 12400 18232
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12452 17746 12480 18022
rect 12544 17814 12572 19178
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18154 12664 19110
rect 12728 18970 12756 19314
rect 13188 19258 13216 20284
rect 13280 19990 13308 20402
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 13372 19514 13400 20402
rect 13464 19854 13492 21626
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13556 20466 13584 21490
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13648 20330 13676 21830
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13648 19938 13676 20266
rect 13740 20058 13768 20402
rect 13832 20330 13860 22442
rect 14108 22094 14136 23258
rect 14384 23118 14412 23684
rect 14372 23112 14424 23118
rect 14372 23054 14424 23060
rect 14476 22506 14504 24618
rect 14660 24614 14688 25638
rect 14936 24954 14964 26318
rect 15108 25696 15160 25702
rect 15108 25638 15160 25644
rect 14924 24948 14976 24954
rect 14924 24890 14976 24896
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24342 14688 24550
rect 14844 24410 14872 24754
rect 15028 24410 15056 24822
rect 15120 24562 15148 25638
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15212 24682 15240 25162
rect 15304 24936 15332 26726
rect 15396 26314 15424 26726
rect 15856 26450 15884 26794
rect 15844 26444 15896 26450
rect 15844 26386 15896 26392
rect 16316 26382 16344 26930
rect 16776 26586 16804 27474
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16868 26858 16896 27270
rect 17328 26994 17356 27406
rect 17500 27328 17552 27334
rect 17500 27270 17552 27276
rect 17960 27328 18012 27334
rect 17960 27270 18012 27276
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18696 27328 18748 27334
rect 18696 27270 18748 27276
rect 17512 26994 17540 27270
rect 17316 26988 17368 26994
rect 17316 26930 17368 26936
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 16856 26852 16908 26858
rect 16856 26794 16908 26800
rect 16868 26586 16896 26794
rect 16764 26580 16816 26586
rect 16764 26522 16816 26528
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 15384 26308 15436 26314
rect 15384 26250 15436 26256
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 15660 25968 15712 25974
rect 15660 25910 15712 25916
rect 15672 25430 15700 25910
rect 15948 25838 15976 26250
rect 16396 26240 16448 26246
rect 16316 26188 16396 26194
rect 16316 26182 16448 26188
rect 16316 26166 16436 26182
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 15936 25832 15988 25838
rect 15936 25774 15988 25780
rect 16132 25498 16160 25842
rect 16316 25702 16344 26166
rect 16764 25900 16816 25906
rect 16764 25842 16816 25848
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16304 25696 16356 25702
rect 16304 25638 16356 25644
rect 16120 25492 16172 25498
rect 16120 25434 16172 25440
rect 15660 25424 15712 25430
rect 15660 25366 15712 25372
rect 15384 24948 15436 24954
rect 15304 24908 15384 24936
rect 15384 24890 15436 24896
rect 15672 24886 15700 25366
rect 16316 25294 16344 25638
rect 16592 25362 16620 25774
rect 16776 25498 16804 25842
rect 17132 25696 17184 25702
rect 17132 25638 17184 25644
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 16304 25288 16356 25294
rect 16304 25230 16356 25236
rect 15568 24880 15620 24886
rect 15568 24822 15620 24828
rect 15660 24880 15712 24886
rect 15660 24822 15712 24828
rect 15200 24676 15252 24682
rect 15200 24618 15252 24624
rect 15476 24608 15528 24614
rect 15120 24556 15476 24562
rect 15120 24550 15528 24556
rect 15120 24534 15516 24550
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 15016 24404 15068 24410
rect 15016 24346 15068 24352
rect 14648 24336 14700 24342
rect 14648 24278 14700 24284
rect 14556 24064 14608 24070
rect 14556 24006 14608 24012
rect 14568 23866 14596 24006
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14568 23594 14596 23666
rect 15028 23594 15056 24346
rect 15108 24200 15160 24206
rect 15108 24142 15160 24148
rect 15198 24168 15254 24177
rect 15120 24070 15148 24142
rect 15198 24103 15254 24112
rect 15108 24064 15160 24070
rect 15108 24006 15160 24012
rect 15120 23866 15148 24006
rect 15108 23860 15160 23866
rect 15108 23802 15160 23808
rect 15212 23662 15240 24103
rect 15488 24070 15516 24534
rect 15580 24410 15608 24822
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15672 24342 15700 24822
rect 16040 24410 16068 25230
rect 16120 25152 16172 25158
rect 16120 25094 16172 25100
rect 16132 24682 16160 25094
rect 16592 24954 16620 25298
rect 16764 25152 16816 25158
rect 16764 25094 16816 25100
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16396 24812 16448 24818
rect 16396 24754 16448 24760
rect 16120 24676 16172 24682
rect 16120 24618 16172 24624
rect 16028 24404 16080 24410
rect 16028 24346 16080 24352
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15108 23656 15160 23662
rect 15108 23598 15160 23604
rect 15200 23656 15252 23662
rect 15200 23598 15252 23604
rect 14556 23588 14608 23594
rect 14556 23530 14608 23536
rect 15016 23588 15068 23594
rect 15016 23530 15068 23536
rect 15028 23186 15056 23530
rect 15120 23322 15148 23598
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15488 23254 15516 24006
rect 15476 23248 15528 23254
rect 15476 23190 15528 23196
rect 15580 23186 15608 24142
rect 15672 23322 15700 24278
rect 16040 24206 16068 24346
rect 16028 24200 16080 24206
rect 16028 24142 16080 24148
rect 16132 24052 16160 24618
rect 16212 24064 16264 24070
rect 16132 24024 16212 24052
rect 15752 23656 15804 23662
rect 15752 23598 15804 23604
rect 15660 23316 15712 23322
rect 15660 23258 15712 23264
rect 15016 23180 15068 23186
rect 15016 23122 15068 23128
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15660 22636 15712 22642
rect 15660 22578 15712 22584
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14924 22432 14976 22438
rect 14924 22374 14976 22380
rect 14016 22066 14136 22094
rect 14016 22030 14044 22066
rect 14936 22030 14964 22374
rect 15396 22234 15424 22578
rect 15568 22432 15620 22438
rect 15488 22392 15568 22420
rect 15384 22228 15436 22234
rect 15384 22170 15436 22176
rect 15488 22030 15516 22392
rect 15568 22374 15620 22380
rect 15672 22234 15700 22578
rect 15660 22228 15712 22234
rect 15660 22170 15712 22176
rect 15764 22030 15792 23598
rect 16028 23316 16080 23322
rect 16028 23258 16080 23264
rect 14004 22024 14056 22030
rect 14004 21966 14056 21972
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15568 22024 15620 22030
rect 15752 22024 15804 22030
rect 15620 21984 15700 22012
rect 15568 21966 15620 21972
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 13924 21554 13952 21830
rect 14016 21554 14044 21966
rect 13912 21548 13964 21554
rect 13912 21490 13964 21496
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 14372 21344 14424 21350
rect 14372 21286 14424 21292
rect 13924 21010 13952 21286
rect 13912 21004 13964 21010
rect 13912 20946 13964 20952
rect 14384 20942 14412 21286
rect 14568 20942 14596 21966
rect 15488 21350 15516 21966
rect 15672 21350 15700 21984
rect 15752 21966 15804 21972
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14292 20602 14320 20878
rect 14384 20806 14412 20878
rect 14372 20800 14424 20806
rect 14372 20742 14424 20748
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 13820 20324 13872 20330
rect 13820 20266 13872 20272
rect 14108 20058 14136 20402
rect 14292 20058 14320 20402
rect 14384 20058 14412 20742
rect 14568 20466 14596 20878
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14372 20052 14424 20058
rect 14372 19994 14424 20000
rect 14292 19938 14320 19994
rect 13648 19910 14320 19938
rect 13452 19848 13504 19854
rect 13452 19790 13504 19796
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13360 19508 13412 19514
rect 13360 19450 13412 19456
rect 13188 19230 13308 19258
rect 13280 19174 13308 19230
rect 13268 19168 13320 19174
rect 13268 19110 13320 19116
rect 13280 18970 13308 19110
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 13268 18964 13320 18970
rect 13268 18906 13320 18912
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13084 18624 13136 18630
rect 13084 18566 13136 18572
rect 13452 18624 13504 18630
rect 13452 18566 13504 18572
rect 13096 18426 13124 18566
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13464 18358 13492 18566
rect 12808 18352 12860 18358
rect 12808 18294 12860 18300
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17882 12756 18022
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12532 17808 12584 17814
rect 12532 17750 12584 17756
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 17066 12020 17546
rect 11980 17060 12032 17066
rect 11980 17002 12032 17008
rect 12084 16794 12112 17682
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12624 17672 12676 17678
rect 12820 17660 12848 18294
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12912 17882 12940 18226
rect 13004 17882 13032 18226
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13176 18080 13228 18086
rect 13174 18048 13176 18057
rect 13228 18048 13230 18057
rect 13174 17983 13230 17992
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 12900 17740 12952 17746
rect 12900 17682 12952 17688
rect 12676 17632 12848 17660
rect 12624 17614 12676 17620
rect 12360 17202 12388 17614
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12452 17134 12480 17478
rect 12912 17202 12940 17682
rect 13280 17270 13308 18158
rect 13556 17678 13584 18906
rect 13648 17678 13676 19722
rect 13740 18222 13768 19910
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13832 19514 13860 19790
rect 14384 19718 14412 19994
rect 14372 19712 14424 19718
rect 15028 19689 15056 21286
rect 15672 20942 15700 21286
rect 15764 21146 15792 21966
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15200 20936 15252 20942
rect 15200 20878 15252 20884
rect 15476 20936 15528 20942
rect 15476 20878 15528 20884
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15212 20602 15240 20878
rect 15488 20806 15516 20878
rect 15568 20868 15620 20874
rect 15568 20810 15620 20816
rect 15384 20800 15436 20806
rect 15384 20742 15436 20748
rect 15476 20800 15528 20806
rect 15476 20742 15528 20748
rect 15200 20596 15252 20602
rect 15200 20538 15252 20544
rect 14372 19654 14424 19660
rect 15014 19680 15070 19689
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 14384 18698 14412 19654
rect 15014 19615 15070 19624
rect 15200 19440 15252 19446
rect 15200 19382 15252 19388
rect 15212 19174 15240 19382
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 14740 19168 14792 19174
rect 14740 19110 14792 19116
rect 15200 19168 15252 19174
rect 15200 19110 15252 19116
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14372 18692 14424 18698
rect 14372 18634 14424 18640
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18426 13952 18566
rect 14384 18426 14412 18634
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 14004 18420 14056 18426
rect 14004 18362 14056 18368
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14016 18306 14044 18362
rect 13924 18278 14044 18306
rect 13924 18222 13952 18278
rect 13728 18216 13780 18222
rect 13728 18158 13780 18164
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13636 17672 13688 17678
rect 13636 17614 13688 17620
rect 13556 17270 13584 17614
rect 13740 17542 13768 18158
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17678 13860 18022
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13268 17264 13320 17270
rect 13268 17206 13320 17212
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 12992 17196 13044 17202
rect 12992 17138 13044 17144
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 13004 16794 13032 17138
rect 13924 17134 13952 18158
rect 14384 17882 14412 18362
rect 14476 18222 14504 18906
rect 14752 18630 14780 19110
rect 15212 18766 15240 19110
rect 15304 18834 15332 19314
rect 15396 19310 15424 20742
rect 15580 20602 15608 20810
rect 15752 20800 15804 20806
rect 15752 20742 15804 20748
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15764 20466 15792 20742
rect 15752 20460 15804 20466
rect 15752 20402 15804 20408
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15488 20058 15516 20334
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15292 18828 15344 18834
rect 15292 18770 15344 18776
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 14740 18624 14792 18630
rect 14740 18566 14792 18572
rect 14752 18290 14780 18566
rect 15120 18426 15148 18634
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15304 18358 15332 18770
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15488 18290 15516 19994
rect 15568 19712 15620 19718
rect 15764 19700 15792 20402
rect 15844 20256 15896 20262
rect 15844 20198 15896 20204
rect 15856 19854 15884 20198
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15620 19672 15792 19700
rect 15568 19654 15620 19660
rect 15580 19514 15608 19654
rect 15568 19508 15620 19514
rect 15568 19450 15620 19456
rect 15580 18970 15608 19450
rect 15752 19372 15804 19378
rect 15752 19314 15804 19320
rect 15660 19304 15712 19310
rect 15660 19246 15712 19252
rect 15672 18970 15700 19246
rect 15764 18970 15792 19314
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 18290 15792 18566
rect 15856 18290 15884 19790
rect 15936 19168 15988 19174
rect 15936 19110 15988 19116
rect 15948 18766 15976 19110
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15476 18284 15528 18290
rect 15476 18226 15528 18232
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 14464 18216 14516 18222
rect 14464 18158 14516 18164
rect 14372 17876 14424 17882
rect 14372 17818 14424 17824
rect 14752 17814 14780 18226
rect 14844 18154 14872 18226
rect 14832 18148 14884 18154
rect 14832 18090 14884 18096
rect 15108 18148 15160 18154
rect 15108 18090 15160 18096
rect 15120 17882 15148 18090
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 14740 17808 14792 17814
rect 14740 17750 14792 17756
rect 15936 17196 15988 17202
rect 15936 17138 15988 17144
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15764 16794 15792 17070
rect 12072 16788 12124 16794
rect 12072 16730 12124 16736
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15948 16590 15976 17138
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16182 13400 16390
rect 14200 16250 14228 16526
rect 14384 16250 14412 16526
rect 13912 16244 13964 16250
rect 14188 16244 14240 16250
rect 13964 16204 14136 16232
rect 13912 16186 13964 16192
rect 11428 16176 11480 16182
rect 11428 16118 11480 16124
rect 11520 16176 11572 16182
rect 11520 16118 11572 16124
rect 11888 16176 11940 16182
rect 11888 16118 11940 16124
rect 12532 16176 12584 16182
rect 12532 16118 12584 16124
rect 13360 16176 13412 16182
rect 13360 16118 13412 16124
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11072 15638 11100 16050
rect 11060 15632 11112 15638
rect 11060 15574 11112 15580
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11072 14414 11100 15574
rect 11256 15366 11284 16050
rect 11440 15366 11468 16118
rect 11532 15366 11560 16118
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 11796 15904 11848 15910
rect 11796 15846 11848 15852
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11520 15360 11572 15366
rect 11520 15302 11572 15308
rect 11256 14958 11284 15302
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11440 13326 11468 15302
rect 11532 13870 11560 15302
rect 11808 15026 11836 15846
rect 11992 15570 12020 15846
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 12176 15366 12204 15846
rect 12452 15706 12480 16050
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12544 15502 12572 16118
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15910 12756 16050
rect 12716 15904 12768 15910
rect 12716 15846 12768 15852
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11624 14618 11652 14758
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11624 14074 11652 14554
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11612 14068 11664 14074
rect 11612 14010 11664 14016
rect 11900 13938 11928 14282
rect 11888 13932 11940 13938
rect 11888 13874 11940 13880
rect 11520 13864 11572 13870
rect 11520 13806 11572 13812
rect 11428 13320 11480 13326
rect 11428 13262 11480 13268
rect 11532 12850 11560 13806
rect 12176 13394 12204 15302
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12360 13734 12388 14962
rect 12544 14822 12572 15438
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 15094 13032 15302
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 12532 14816 12584 14822
rect 12532 14758 12584 14764
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12164 13388 12216 13394
rect 12164 13330 12216 13336
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12442 11560 12786
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 12360 11830 12388 13670
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12452 12850 12480 13262
rect 12544 12986 12572 14758
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12452 12238 12480 12786
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12544 12434 12572 12718
rect 12544 12406 12664 12434
rect 12636 12238 12664 12406
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 13096 11898 13124 13126
rect 13372 11898 13400 16118
rect 14108 16114 14136 16204
rect 14188 16186 14240 16192
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14186 16144 14242 16153
rect 14096 16108 14148 16114
rect 14186 16079 14188 16088
rect 14096 16050 14148 16056
rect 14240 16079 14242 16088
rect 14280 16108 14332 16114
rect 14188 16050 14240 16056
rect 14280 16050 14332 16056
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 13648 12850 13676 13874
rect 13924 12850 13952 13874
rect 14200 13802 14228 15438
rect 14292 15366 14320 16050
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14384 15162 14412 15438
rect 15304 15162 15332 15438
rect 15396 15162 15424 15982
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15672 15706 15700 15846
rect 15948 15706 15976 16526
rect 16040 16250 16068 23258
rect 16132 20806 16160 24024
rect 16212 24006 16264 24012
rect 16408 23866 16436 24754
rect 16776 24750 16804 25094
rect 17144 24954 17172 25638
rect 17132 24948 17184 24954
rect 17132 24890 17184 24896
rect 17224 24880 17276 24886
rect 17224 24822 17276 24828
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16776 23662 16804 24686
rect 17052 24206 17080 24754
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 17236 24070 17264 24822
rect 17328 24342 17356 26930
rect 17512 26586 17540 26930
rect 17500 26580 17552 26586
rect 17500 26522 17552 26528
rect 17972 25838 18000 27270
rect 18524 26994 18552 27270
rect 18708 26994 18736 27270
rect 19352 27062 19380 27814
rect 19444 27674 19472 27950
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19536 27606 19564 27950
rect 19524 27600 19576 27606
rect 19524 27542 19576 27548
rect 19536 27418 19564 27542
rect 19444 27390 19564 27418
rect 19340 27056 19392 27062
rect 19340 26998 19392 27004
rect 18420 26988 18472 26994
rect 18420 26930 18472 26936
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18788 26988 18840 26994
rect 19444 26976 19472 27390
rect 19812 27316 19840 28154
rect 19996 27554 20024 28358
rect 20088 28150 20116 28614
rect 20352 28620 20404 28626
rect 20352 28562 20404 28568
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 20076 28144 20128 28150
rect 20076 28086 20128 28092
rect 20180 28014 20208 28426
rect 20076 28008 20128 28014
rect 20076 27950 20128 27956
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 20088 27674 20116 27950
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 19996 27526 20116 27554
rect 19812 27288 20024 27316
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19524 26988 19576 26994
rect 19444 26948 19524 26976
rect 18788 26930 18840 26936
rect 19524 26930 19576 26936
rect 18432 26586 18460 26930
rect 18420 26580 18472 26586
rect 18420 26522 18472 26528
rect 18052 26376 18104 26382
rect 18052 26318 18104 26324
rect 18236 26376 18288 26382
rect 18236 26318 18288 26324
rect 18064 26042 18092 26318
rect 18052 26036 18104 26042
rect 18052 25978 18104 25984
rect 18248 25974 18276 26318
rect 18708 26042 18736 26930
rect 18800 26382 18828 26930
rect 19340 26920 19392 26926
rect 19392 26880 19472 26908
rect 19340 26862 19392 26868
rect 19340 26784 19392 26790
rect 19340 26726 19392 26732
rect 19352 26586 19380 26726
rect 19340 26580 19392 26586
rect 19340 26522 19392 26528
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18236 25968 18288 25974
rect 18236 25910 18288 25916
rect 17868 25832 17920 25838
rect 17868 25774 17920 25780
rect 17960 25832 18012 25838
rect 17960 25774 18012 25780
rect 17684 25152 17736 25158
rect 17684 25094 17736 25100
rect 17316 24336 17368 24342
rect 17316 24278 17368 24284
rect 17408 24336 17460 24342
rect 17408 24278 17460 24284
rect 17316 24200 17368 24206
rect 17316 24142 17368 24148
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17144 23798 17172 24006
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17328 23662 17356 24142
rect 17420 24041 17448 24278
rect 17696 24138 17724 25094
rect 17880 24206 17908 25774
rect 17972 25158 18000 25774
rect 18248 25498 18276 25910
rect 18236 25492 18288 25498
rect 18236 25434 18288 25440
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 18800 24818 18828 26318
rect 18880 25968 18932 25974
rect 18880 25910 18932 25916
rect 18892 25294 18920 25910
rect 19444 25906 19472 26880
rect 19536 26450 19564 26930
rect 19524 26444 19576 26450
rect 19524 26386 19576 26392
rect 19996 26382 20024 27288
rect 20088 27130 20116 27526
rect 20180 27470 20208 27950
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 20076 27124 20128 27130
rect 20076 27066 20128 27072
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20088 26586 20116 26930
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 19984 26376 20036 26382
rect 19984 26318 20036 26324
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19892 26036 19944 26042
rect 19996 26024 20024 26318
rect 19944 25996 20024 26024
rect 19892 25978 19944 25984
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 18972 25696 19024 25702
rect 18972 25638 19024 25644
rect 18984 25498 19012 25638
rect 18972 25492 19024 25498
rect 18972 25434 19024 25440
rect 20088 25362 20116 25842
rect 20272 25498 20300 26930
rect 20364 26586 20392 28562
rect 33048 28484 33100 28490
rect 33048 28426 33100 28432
rect 21548 28416 21600 28422
rect 21548 28358 21600 28364
rect 32588 28416 32640 28422
rect 32588 28358 32640 28364
rect 21560 28218 21588 28358
rect 21456 28212 21508 28218
rect 21456 28154 21508 28160
rect 21548 28212 21600 28218
rect 21548 28154 21600 28160
rect 21088 28076 21140 28082
rect 21088 28018 21140 28024
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20720 26988 20772 26994
rect 20548 26948 20720 26976
rect 20352 26580 20404 26586
rect 20352 26522 20404 26528
rect 20364 25906 20392 26522
rect 20444 26376 20496 26382
rect 20548 26364 20576 26948
rect 20720 26930 20772 26936
rect 20824 26926 20852 27814
rect 20812 26920 20864 26926
rect 20812 26862 20864 26868
rect 20496 26336 20576 26364
rect 20444 26318 20496 26324
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20364 25378 20392 25842
rect 20456 25838 20484 26182
rect 20548 25906 20576 26336
rect 21100 26042 21128 28018
rect 21468 27674 21496 28154
rect 22560 28076 22612 28082
rect 22560 28018 22612 28024
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21456 27328 21508 27334
rect 21456 27270 21508 27276
rect 21468 26586 21496 27270
rect 22572 27130 22600 28018
rect 32600 27878 32628 28358
rect 32956 28008 33008 28014
rect 32956 27950 33008 27956
rect 22836 27872 22888 27878
rect 22836 27814 22888 27820
rect 30656 27872 30708 27878
rect 30656 27814 30708 27820
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 31024 27872 31076 27878
rect 31024 27814 31076 27820
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 32588 27872 32640 27878
rect 32588 27814 32640 27820
rect 22848 27674 22876 27814
rect 22836 27668 22888 27674
rect 22836 27610 22888 27616
rect 23664 27532 23716 27538
rect 23664 27474 23716 27480
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23480 27464 23532 27470
rect 23480 27406 23532 27412
rect 22560 27124 22612 27130
rect 22560 27066 22612 27072
rect 23400 27062 23428 27406
rect 23492 27130 23520 27406
rect 23676 27130 23704 27474
rect 30668 27470 30696 27814
rect 30840 27532 30892 27538
rect 30840 27474 30892 27480
rect 29736 27464 29788 27470
rect 29736 27406 29788 27412
rect 30656 27464 30708 27470
rect 30852 27418 30880 27474
rect 30708 27412 30880 27418
rect 30656 27406 30880 27412
rect 25964 27396 26016 27402
rect 25964 27338 26016 27344
rect 25976 27130 26004 27338
rect 26700 27328 26752 27334
rect 26700 27270 26752 27276
rect 27068 27328 27120 27334
rect 27068 27270 27120 27276
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 26712 27130 26740 27270
rect 27080 27130 27108 27270
rect 27264 27130 27292 27270
rect 29748 27130 29776 27406
rect 30668 27390 30880 27406
rect 30012 27328 30064 27334
rect 30012 27270 30064 27276
rect 23480 27124 23532 27130
rect 23480 27066 23532 27072
rect 23664 27124 23716 27130
rect 23664 27066 23716 27072
rect 25964 27124 26016 27130
rect 25964 27066 26016 27072
rect 26700 27124 26752 27130
rect 26700 27066 26752 27072
rect 27068 27124 27120 27130
rect 27068 27066 27120 27072
rect 27252 27124 27304 27130
rect 27252 27066 27304 27072
rect 29736 27124 29788 27130
rect 29736 27066 29788 27072
rect 21640 27056 21692 27062
rect 21640 26998 21692 27004
rect 23388 27056 23440 27062
rect 23388 26998 23440 27004
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21652 26450 21680 26998
rect 26712 26994 26740 27066
rect 21824 26988 21876 26994
rect 21824 26930 21876 26936
rect 22284 26988 22336 26994
rect 22284 26930 22336 26936
rect 24860 26988 24912 26994
rect 24860 26930 24912 26936
rect 26700 26988 26752 26994
rect 26700 26930 26752 26936
rect 26884 26988 26936 26994
rect 26884 26930 26936 26936
rect 21836 26586 21864 26930
rect 22296 26586 22324 26930
rect 22376 26852 22428 26858
rect 22376 26794 22428 26800
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 21824 26580 21876 26586
rect 21824 26522 21876 26528
rect 22100 26580 22152 26586
rect 22100 26522 22152 26528
rect 22284 26580 22336 26586
rect 22284 26522 22336 26528
rect 21640 26444 21692 26450
rect 21640 26386 21692 26392
rect 21548 26376 21600 26382
rect 21548 26318 21600 26324
rect 21560 26042 21588 26318
rect 21088 26036 21140 26042
rect 21088 25978 21140 25984
rect 21548 26036 21600 26042
rect 21548 25978 21600 25984
rect 20536 25900 20588 25906
rect 20536 25842 20588 25848
rect 20444 25832 20496 25838
rect 20444 25774 20496 25780
rect 21272 25832 21324 25838
rect 21272 25774 21324 25780
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 20272 25350 20392 25378
rect 20272 25294 20300 25350
rect 20732 25294 20760 25638
rect 21284 25498 21312 25774
rect 21272 25492 21324 25498
rect 21272 25434 21324 25440
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 18236 24812 18288 24818
rect 18236 24754 18288 24760
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 18248 24614 18276 24754
rect 18892 24682 18920 25230
rect 18880 24676 18932 24682
rect 18880 24618 18932 24624
rect 19248 24676 19300 24682
rect 19248 24618 19300 24624
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18328 24608 18380 24614
rect 18328 24550 18380 24556
rect 18248 24410 18276 24550
rect 18236 24404 18288 24410
rect 18236 24346 18288 24352
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17406 24032 17462 24041
rect 17406 23967 17462 23976
rect 16764 23656 16816 23662
rect 16764 23598 16816 23604
rect 17316 23656 17368 23662
rect 17316 23598 17368 23604
rect 16212 22024 16264 22030
rect 16212 21966 16264 21972
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16224 21690 16252 21966
rect 16316 21894 16344 21966
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16316 21729 16344 21830
rect 16302 21720 16358 21729
rect 16212 21684 16264 21690
rect 16500 21690 16528 21966
rect 16302 21655 16358 21664
rect 16488 21684 16540 21690
rect 16212 21626 16264 21632
rect 16488 21626 16540 21632
rect 16304 20868 16356 20874
rect 16304 20810 16356 20816
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16316 20398 16344 20810
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16316 20058 16344 20334
rect 16304 20052 16356 20058
rect 16304 19994 16356 20000
rect 16580 19712 16632 19718
rect 16578 19680 16580 19689
rect 16632 19680 16634 19689
rect 16578 19615 16634 19624
rect 16578 19544 16634 19553
rect 16120 19508 16172 19514
rect 16578 19479 16580 19488
rect 16120 19450 16172 19456
rect 16632 19479 16634 19488
rect 16672 19508 16724 19514
rect 16580 19450 16632 19456
rect 16672 19450 16724 19456
rect 16132 18290 16160 19450
rect 16684 19378 16712 19450
rect 16672 19372 16724 19378
rect 16672 19314 16724 19320
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16592 18902 16620 19246
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16580 18692 16632 18698
rect 16580 18634 16632 18640
rect 16592 18426 16620 18634
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 16132 16590 16160 17478
rect 16592 17270 16620 17614
rect 16580 17264 16632 17270
rect 16580 17206 16632 17212
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 16590 16436 16934
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16040 16114 16068 16186
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15660 15700 15712 15706
rect 15936 15700 15988 15706
rect 15712 15660 15792 15688
rect 15660 15642 15712 15648
rect 15764 15502 15792 15660
rect 15936 15642 15988 15648
rect 16040 15502 16068 16050
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 14372 15156 14424 15162
rect 14372 15098 14424 15104
rect 15292 15156 15344 15162
rect 15292 15098 15344 15104
rect 15384 15156 15436 15162
rect 15384 15098 15436 15104
rect 15108 15088 15160 15094
rect 15108 15030 15160 15036
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 13636 12844 13688 12850
rect 13636 12786 13688 12792
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13648 12102 13676 12786
rect 14108 12442 14136 12786
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14384 12374 14412 14418
rect 14556 13864 14608 13870
rect 14556 13806 14608 13812
rect 14568 13326 14596 13806
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14660 13530 14688 13670
rect 14752 13530 14780 13670
rect 14648 13524 14700 13530
rect 14648 13466 14700 13472
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14568 12764 14596 13262
rect 14660 12986 14688 13262
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14648 12776 14700 12782
rect 14568 12736 14648 12764
rect 14648 12718 14700 12724
rect 14464 12708 14516 12714
rect 14464 12650 14516 12656
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14476 12238 14504 12650
rect 14752 12238 14780 13466
rect 14844 12782 14872 14894
rect 14936 14414 14964 14962
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14936 14074 14964 14350
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15028 13802 15056 14214
rect 15016 13796 15068 13802
rect 15016 13738 15068 13744
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15028 12646 15056 13738
rect 15120 12850 15148 15030
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15212 14482 15240 14962
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15672 14414 15700 15438
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 14822 15792 15302
rect 16040 15162 16068 15438
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15764 14414 15792 14758
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15948 14414 15976 14554
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 13326 15240 13670
rect 15396 13394 15424 14214
rect 15580 14074 15608 14282
rect 15672 14074 15700 14350
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15936 13456 15988 13462
rect 15936 13398 15988 13404
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15304 12986 15332 13262
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15120 12442 15148 12786
rect 15488 12714 15516 13262
rect 15948 12986 15976 13398
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15764 12646 15792 12718
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15014 12336 15070 12345
rect 14924 12300 14976 12306
rect 14976 12280 15014 12288
rect 15658 12336 15714 12345
rect 14976 12271 15070 12280
rect 15568 12300 15620 12306
rect 14976 12260 15056 12271
rect 14924 12242 14976 12248
rect 15658 12271 15660 12280
rect 15568 12242 15620 12248
rect 15712 12271 15714 12280
rect 15660 12242 15712 12248
rect 13912 12232 13964 12238
rect 13912 12174 13964 12180
rect 14464 12232 14516 12238
rect 14464 12174 14516 12180
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13924 11898 13952 12174
rect 13084 11892 13136 11898
rect 13084 11834 13136 11840
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 12348 11824 12400 11830
rect 12348 11766 12400 11772
rect 15580 11762 15608 12242
rect 15764 12238 15792 12582
rect 15948 12238 15976 12786
rect 15752 12232 15804 12238
rect 15936 12232 15988 12238
rect 15752 12174 15804 12180
rect 15934 12200 15936 12209
rect 15988 12200 15990 12209
rect 15934 12135 15990 12144
rect 16040 11762 16068 14282
rect 16132 13530 16160 16526
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16212 14816 16264 14822
rect 16212 14758 16264 14764
rect 16224 14618 16252 14758
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 16224 14074 16252 14554
rect 16500 14362 16528 15302
rect 16684 15162 16712 16526
rect 16776 15978 16804 23598
rect 17696 23526 17724 24074
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 16868 22506 16896 23462
rect 18248 23186 18276 24346
rect 18340 24206 18368 24550
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18340 23798 18368 24142
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18616 23730 18644 24346
rect 19260 24206 19288 24618
rect 19352 24410 19380 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19616 24608 19668 24614
rect 19616 24550 19668 24556
rect 19628 24410 19656 24550
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19616 24404 19668 24410
rect 19616 24346 19668 24352
rect 19248 24200 19300 24206
rect 19248 24142 19300 24148
rect 19984 24200 20036 24206
rect 19984 24142 20036 24148
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 18420 23724 18472 23730
rect 18420 23666 18472 23672
rect 18604 23724 18656 23730
rect 18604 23666 18656 23672
rect 18432 23322 18460 23666
rect 19996 23662 20024 24142
rect 20272 23798 20300 25230
rect 21548 24676 21600 24682
rect 21548 24618 21600 24624
rect 20996 24336 21048 24342
rect 20996 24278 21048 24284
rect 20548 24138 20852 24154
rect 20548 24132 20864 24138
rect 20548 24126 20812 24132
rect 20260 23792 20312 23798
rect 20260 23734 20312 23740
rect 20444 23724 20496 23730
rect 20548 23712 20576 24126
rect 20812 24074 20864 24080
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20496 23684 20576 23712
rect 20626 23760 20682 23769
rect 20626 23695 20682 23704
rect 20444 23666 20496 23672
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 18420 23316 18472 23322
rect 18420 23258 18472 23264
rect 18236 23180 18288 23186
rect 18236 23122 18288 23128
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 18236 23044 18288 23050
rect 18236 22986 18288 22992
rect 18248 22642 18276 22986
rect 18512 22976 18564 22982
rect 18512 22918 18564 22924
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 17684 22636 17736 22642
rect 17684 22578 17736 22584
rect 17868 22636 17920 22642
rect 17868 22578 17920 22584
rect 18052 22636 18104 22642
rect 18052 22578 18104 22584
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 16856 22500 16908 22506
rect 16856 22442 16908 22448
rect 16960 22234 16988 22578
rect 17040 22432 17092 22438
rect 17040 22374 17092 22380
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 16856 22024 16908 22030
rect 16856 21966 16908 21972
rect 16960 21978 16988 22170
rect 17052 22098 17080 22374
rect 17040 22092 17092 22098
rect 17040 22034 17092 22040
rect 16868 21894 16896 21966
rect 16960 21962 17632 21978
rect 16960 21956 17644 21962
rect 16960 21950 17592 21956
rect 17592 21898 17644 21904
rect 16856 21888 16908 21894
rect 16856 21830 16908 21836
rect 17224 21888 17276 21894
rect 17224 21830 17276 21836
rect 17236 21690 17264 21830
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17500 21548 17552 21554
rect 17500 21490 17552 21496
rect 17512 21146 17540 21490
rect 17224 21140 17276 21146
rect 17224 21082 17276 21088
rect 17500 21140 17552 21146
rect 17500 21082 17552 21088
rect 17040 20528 17092 20534
rect 17040 20470 17092 20476
rect 17052 20262 17080 20470
rect 17236 20466 17264 21082
rect 17316 20936 17368 20942
rect 17316 20878 17368 20884
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17040 20256 17092 20262
rect 17040 20198 17092 20204
rect 17052 18766 17080 20198
rect 17236 18766 17264 20402
rect 17328 20330 17356 20878
rect 17316 20324 17368 20330
rect 17316 20266 17368 20272
rect 17328 19174 17356 20266
rect 17604 20058 17632 21898
rect 17696 21690 17724 22578
rect 17776 22160 17828 22166
rect 17776 22102 17828 22108
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17696 20602 17724 21626
rect 17788 21554 17816 22102
rect 17880 22030 17908 22578
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17880 21554 17908 21966
rect 18064 21690 18092 22578
rect 18524 22506 18552 22918
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 18052 21684 18104 21690
rect 18052 21626 18104 21632
rect 17972 21570 18000 21626
rect 17972 21554 18092 21570
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17868 21548 17920 21554
rect 17972 21548 18104 21554
rect 17972 21542 18052 21548
rect 17868 21490 17920 21496
rect 18052 21490 18104 21496
rect 17868 21412 17920 21418
rect 17868 21354 17920 21360
rect 17880 21146 17908 21354
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17972 20398 18000 20878
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17592 20052 17644 20058
rect 17592 19994 17644 20000
rect 17788 19922 17816 20198
rect 18524 19990 18552 22442
rect 18696 22024 18748 22030
rect 18696 21966 18748 21972
rect 18708 21350 18736 21966
rect 18696 21344 18748 21350
rect 18696 21286 18748 21292
rect 18512 19984 18564 19990
rect 18512 19926 18564 19932
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17512 19514 17540 19654
rect 17500 19508 17552 19514
rect 17500 19450 17552 19456
rect 17788 19310 17816 19858
rect 17958 19544 18014 19553
rect 17958 19479 17960 19488
rect 18012 19479 18014 19488
rect 17960 19450 18012 19456
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17776 19304 17828 19310
rect 17776 19246 17828 19252
rect 17316 19168 17368 19174
rect 17316 19110 17368 19116
rect 17696 18970 17724 19246
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17972 18834 18000 19314
rect 18064 18970 18092 19314
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17052 18086 17080 18702
rect 17960 18624 18012 18630
rect 18156 18612 18184 19246
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18420 19168 18472 19174
rect 18420 19110 18472 19116
rect 18340 18766 18368 19110
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18432 18630 18460 19110
rect 18012 18584 18184 18612
rect 18420 18624 18472 18630
rect 17960 18566 18012 18572
rect 18420 18566 18472 18572
rect 17972 18290 18000 18566
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 17040 18080 17092 18086
rect 17040 18022 17092 18028
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17408 17060 17460 17066
rect 17408 17002 17460 17008
rect 17420 16794 17448 17002
rect 17408 16788 17460 16794
rect 17408 16730 17460 16736
rect 16856 16584 16908 16590
rect 16856 16526 16908 16532
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16684 14414 16712 15098
rect 16764 14544 16816 14550
rect 16764 14486 16816 14492
rect 16672 14408 16724 14414
rect 16408 14334 16620 14362
rect 16672 14350 16724 14356
rect 16212 14068 16264 14074
rect 16212 14010 16264 14016
rect 16408 13530 16436 14334
rect 16592 14278 16620 14334
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16580 14272 16632 14278
rect 16580 14214 16632 14220
rect 16500 14074 16528 14214
rect 16776 14074 16804 14486
rect 16868 14074 16896 16526
rect 17880 15994 17908 18022
rect 17972 17202 18000 18226
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 17880 15978 18000 15994
rect 17224 15972 17276 15978
rect 17880 15972 18012 15978
rect 17880 15966 17960 15972
rect 17224 15914 17276 15920
rect 17960 15914 18012 15920
rect 16948 15564 17000 15570
rect 16948 15506 17000 15512
rect 16960 14346 16988 15506
rect 17236 15502 17264 15914
rect 17776 15904 17828 15910
rect 17776 15846 17828 15852
rect 17788 15502 17816 15846
rect 18156 15706 18184 18226
rect 18432 18154 18460 18566
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18328 17264 18380 17270
rect 18328 17206 18380 17212
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18248 16794 18276 17070
rect 18236 16788 18288 16794
rect 18236 16730 18288 16736
rect 18340 16590 18368 17206
rect 18800 16674 18828 23054
rect 19996 22982 20024 23598
rect 20456 23118 20484 23666
rect 20640 23662 20668 23695
rect 20628 23656 20680 23662
rect 20628 23598 20680 23604
rect 20812 23656 20864 23662
rect 20812 23598 20864 23604
rect 20824 23322 20852 23598
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20916 23118 20944 24074
rect 21008 23866 21036 24278
rect 21088 24268 21140 24274
rect 21088 24210 21140 24216
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 21100 23322 21128 24210
rect 21180 24064 21232 24070
rect 21180 24006 21232 24012
rect 21192 23798 21220 24006
rect 21180 23792 21232 23798
rect 21180 23734 21232 23740
rect 21088 23316 21140 23322
rect 21088 23258 21140 23264
rect 21192 23254 21220 23734
rect 21272 23724 21324 23730
rect 21456 23724 21508 23730
rect 21324 23684 21404 23712
rect 21272 23666 21324 23672
rect 21180 23248 21232 23254
rect 21180 23190 21232 23196
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20628 23112 20680 23118
rect 20904 23112 20956 23118
rect 20680 23072 20760 23100
rect 20628 23054 20680 23060
rect 19984 22976 20036 22982
rect 19984 22918 20036 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19536 19922 19564 20198
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18892 18426 18920 19314
rect 18972 19304 19024 19310
rect 19024 19264 19196 19292
rect 18972 19246 19024 19252
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18984 18698 19012 18838
rect 19076 18698 19104 18906
rect 18972 18692 19024 18698
rect 18972 18634 19024 18640
rect 19064 18692 19116 18698
rect 19064 18634 19116 18640
rect 18984 18426 19012 18634
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18880 18284 18932 18290
rect 18984 18272 19012 18362
rect 18932 18244 19012 18272
rect 19064 18284 19116 18290
rect 18880 18226 18932 18232
rect 19064 18226 19116 18232
rect 19076 18086 19104 18226
rect 19168 18086 19196 19264
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19260 18970 19288 19110
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19340 18828 19392 18834
rect 19260 18788 19340 18816
rect 19260 18290 19288 18788
rect 19340 18770 19392 18776
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19444 18630 19472 18702
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 18290 19472 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19248 18284 19300 18290
rect 19248 18226 19300 18232
rect 19432 18284 19484 18290
rect 19432 18226 19484 18232
rect 19064 18080 19116 18086
rect 19064 18022 19116 18028
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19338 18048 19394 18057
rect 19338 17983 19394 17992
rect 19352 17678 19380 17983
rect 19444 17882 19472 18226
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 16794 20024 22918
rect 20456 22710 20484 23054
rect 20732 22778 20760 23072
rect 20904 23054 20956 23060
rect 21376 22982 21404 23684
rect 21456 23666 21508 23672
rect 21468 23322 21496 23666
rect 21456 23316 21508 23322
rect 21456 23258 21508 23264
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20732 22234 20760 22714
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 21180 22160 21232 22166
rect 21180 22102 21232 22108
rect 21192 22030 21220 22102
rect 21284 22098 21312 22578
rect 21376 22234 21404 22918
rect 21364 22228 21416 22234
rect 21364 22170 21416 22176
rect 21272 22092 21324 22098
rect 21272 22034 21324 22040
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20904 21888 20956 21894
rect 20904 21830 20956 21836
rect 20364 21010 20392 21830
rect 20916 21554 20944 21830
rect 21192 21690 21220 21966
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 20444 21548 20496 21554
rect 20444 21490 20496 21496
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20364 20466 20392 20946
rect 20456 20602 20484 21490
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20352 20324 20404 20330
rect 20352 20266 20404 20272
rect 20364 19802 20392 20266
rect 20456 20058 20484 20538
rect 20548 20466 20576 21490
rect 20732 20942 20760 21490
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20482 20760 20878
rect 20916 20602 20944 21490
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20536 20460 20588 20466
rect 20732 20454 20852 20482
rect 20536 20402 20588 20408
rect 20824 20398 20852 20454
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20628 20324 20680 20330
rect 20628 20266 20680 20272
rect 20444 20052 20496 20058
rect 20444 19994 20496 20000
rect 20640 19990 20668 20266
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20628 19848 20680 19854
rect 20364 19786 20484 19802
rect 20628 19790 20680 19796
rect 20364 19780 20496 19786
rect 20364 19774 20444 19780
rect 20444 19722 20496 19728
rect 20352 19712 20404 19718
rect 20352 19654 20404 19660
rect 20364 19514 20392 19654
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20088 18358 20116 19314
rect 20364 18902 20392 19450
rect 20456 19378 20484 19722
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20640 19174 20668 19790
rect 20628 19168 20680 19174
rect 20628 19110 20680 19116
rect 20352 18896 20404 18902
rect 20352 18838 20404 18844
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20076 18352 20128 18358
rect 20076 18294 20128 18300
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 20088 17202 20116 17546
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20456 17066 20484 18566
rect 20444 17060 20496 17066
rect 20444 17002 20496 17008
rect 20456 16794 20484 17002
rect 19984 16788 20036 16794
rect 19984 16730 20036 16736
rect 20444 16788 20496 16794
rect 20444 16730 20496 16736
rect 18800 16646 18920 16674
rect 18328 16584 18380 16590
rect 18328 16526 18380 16532
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18144 15700 18196 15706
rect 18144 15642 18196 15648
rect 17040 15496 17092 15502
rect 17040 15438 17092 15444
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17224 15496 17276 15502
rect 17224 15438 17276 15444
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17052 15094 17080 15438
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 17144 15026 17172 15438
rect 17132 15020 17184 15026
rect 17132 14962 17184 14968
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16856 14068 16908 14074
rect 16856 14010 16908 14016
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16592 13326 16620 13806
rect 16580 13320 16632 13326
rect 16776 13308 16804 14010
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16960 13530 16988 13874
rect 17052 13530 17080 14894
rect 17236 14618 17264 15438
rect 18156 15094 18184 15438
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 17500 14952 17552 14958
rect 17500 14894 17552 14900
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17316 14884 17368 14890
rect 17316 14826 17368 14832
rect 17224 14612 17276 14618
rect 17224 14554 17276 14560
rect 17328 14074 17356 14826
rect 17512 14482 17540 14894
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17316 14068 17368 14074
rect 17316 14010 17368 14016
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 13320 17000 13326
rect 16776 13280 16948 13308
rect 16580 13262 16632 13268
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16120 12640 16172 12646
rect 16408 12628 16436 12786
rect 16488 12708 16540 12714
rect 16488 12650 16540 12656
rect 16120 12582 16172 12588
rect 16224 12600 16436 12628
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 16028 11756 16080 11762
rect 16028 11698 16080 11704
rect 16132 11626 16160 12582
rect 16224 12442 16252 12600
rect 16500 12458 16528 12650
rect 16212 12436 16264 12442
rect 16316 12430 16528 12458
rect 16316 12406 16436 12430
rect 16212 12378 16264 12384
rect 16408 11762 16436 12406
rect 16580 12368 16632 12374
rect 16632 12328 16804 12356
rect 16580 12310 16632 12316
rect 16776 12170 16804 12328
rect 16868 12238 16896 13280
rect 16948 13262 17000 13268
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 17040 13184 17092 13190
rect 17040 13126 17092 13132
rect 17052 12850 17080 13126
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16592 12050 16620 12106
rect 17144 12050 17172 13262
rect 17328 12850 17356 14010
rect 17604 13530 17632 14554
rect 17696 14414 17724 14894
rect 18156 14890 18184 15030
rect 18432 15026 18460 15846
rect 18524 15502 18552 16390
rect 18708 16250 18736 16390
rect 18696 16244 18748 16250
rect 18696 16186 18748 16192
rect 18800 15910 18828 16526
rect 18892 16182 18920 16646
rect 19064 16652 19116 16658
rect 19064 16594 19116 16600
rect 18880 16176 18932 16182
rect 18878 16144 18880 16153
rect 18932 16144 18934 16153
rect 18878 16079 18934 16088
rect 18788 15904 18840 15910
rect 18788 15846 18840 15852
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18144 14884 18196 14890
rect 18144 14826 18196 14832
rect 18156 14618 18184 14826
rect 18144 14612 18196 14618
rect 18144 14554 18196 14560
rect 18524 14414 18552 15438
rect 19076 15366 19104 16594
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19064 15360 19116 15366
rect 19064 15302 19116 15308
rect 18696 15088 18748 15094
rect 18696 15030 18748 15036
rect 18708 14482 18736 15030
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 17972 14074 18000 14350
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 14074 18092 14282
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 17592 13524 17644 13530
rect 17592 13466 17644 13472
rect 17604 12986 17632 13466
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17512 12442 17540 12922
rect 17880 12850 17908 13330
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17500 12436 17552 12442
rect 17500 12378 17552 12384
rect 17224 12232 17276 12238
rect 17222 12200 17224 12209
rect 17276 12200 17278 12209
rect 17222 12135 17278 12144
rect 16592 12022 17172 12050
rect 17880 11898 17908 12786
rect 17972 12442 18000 14010
rect 18064 13326 18092 14010
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18156 13190 18184 14350
rect 18248 14074 18276 14350
rect 18236 14068 18288 14074
rect 18236 14010 18288 14016
rect 18248 13530 18276 14010
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18236 13524 18288 13530
rect 18236 13466 18288 13472
rect 18248 13326 18276 13466
rect 18432 13326 18460 13942
rect 18236 13320 18288 13326
rect 18236 13262 18288 13268
rect 18420 13320 18472 13326
rect 18420 13262 18472 13268
rect 18144 13184 18196 13190
rect 18144 13126 18196 13132
rect 18248 12646 18276 13262
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18524 12986 18552 13194
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 19076 12850 19104 15302
rect 19260 15026 19288 16050
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19248 15020 19300 15026
rect 19248 14962 19300 14968
rect 19352 14890 19380 15982
rect 20352 15904 20404 15910
rect 20352 15846 20404 15852
rect 20260 15632 20312 15638
rect 20260 15574 20312 15580
rect 20076 15564 20128 15570
rect 20076 15506 20128 15512
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15094 19472 15302
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15094 20116 15506
rect 20272 15094 20300 15574
rect 20364 15502 20392 15846
rect 20444 15632 20496 15638
rect 20444 15574 20496 15580
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20364 15162 20392 15438
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 20076 15088 20128 15094
rect 20076 15030 20128 15036
rect 20260 15088 20312 15094
rect 20260 15030 20312 15036
rect 19616 14952 19668 14958
rect 19616 14894 19668 14900
rect 19340 14884 19392 14890
rect 19340 14826 19392 14832
rect 19248 14408 19300 14414
rect 19248 14350 19300 14356
rect 19156 13728 19208 13734
rect 19156 13670 19208 13676
rect 19168 13394 19196 13670
rect 19260 13530 19288 14350
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12986 19196 13330
rect 19260 12986 19288 13466
rect 19352 13258 19380 14826
rect 19432 14816 19484 14822
rect 19432 14758 19484 14764
rect 19444 14346 19472 14758
rect 19628 14618 19656 14894
rect 20088 14822 20116 15030
rect 20076 14816 20128 14822
rect 20076 14758 20128 14764
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 20088 14482 20116 14758
rect 20364 14498 20392 15098
rect 20456 14618 20484 15574
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20076 14476 20128 14482
rect 20364 14470 20484 14498
rect 20076 14418 20128 14424
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19524 14068 19576 14074
rect 19524 14010 19576 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19444 13462 19472 13874
rect 19536 13530 19564 14010
rect 20088 13870 20116 14418
rect 20168 14408 20220 14414
rect 20168 14350 20220 14356
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20180 14074 20208 14350
rect 20272 14074 20300 14350
rect 20364 14074 20392 14350
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20456 13870 20484 14470
rect 20548 14414 20576 14962
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20548 14006 20576 14350
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20444 13864 20496 13870
rect 20444 13806 20496 13812
rect 19524 13524 19576 13530
rect 19524 13466 19576 13472
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19156 12980 19208 12986
rect 19156 12922 19208 12928
rect 19248 12980 19300 12986
rect 19248 12922 19300 12928
rect 19352 12850 19380 13194
rect 19444 12986 19472 13398
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19800 12980 19852 12986
rect 19800 12922 19852 12928
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 19064 12844 19116 12850
rect 19064 12786 19116 12792
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 18236 12640 18288 12646
rect 18236 12582 18288 12588
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 17972 12306 18000 12378
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17868 11892 17920 11898
rect 17868 11834 17920 11840
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 17972 11354 18000 12242
rect 18236 12164 18288 12170
rect 18340 12152 18368 12582
rect 18432 12442 18460 12786
rect 18696 12776 18748 12782
rect 18696 12718 18748 12724
rect 18420 12436 18472 12442
rect 18420 12378 18472 12384
rect 18288 12124 18368 12152
rect 18236 12106 18288 12112
rect 18432 11762 18460 12378
rect 18708 12238 18736 12718
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19444 12238 19472 12650
rect 19812 12306 19840 12922
rect 19984 12844 20036 12850
rect 19984 12786 20036 12792
rect 19996 12442 20024 12786
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20088 12306 20116 13806
rect 20272 13258 20300 13806
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20364 12434 20392 13670
rect 20456 13530 20484 13806
rect 20444 13524 20496 13530
rect 20444 13466 20496 13472
rect 20548 13326 20576 13942
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20272 12406 20392 12434
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18696 12232 18748 12238
rect 18696 12174 18748 12180
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 18524 11762 18552 12174
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18420 11756 18472 11762
rect 18420 11698 18472 11704
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 17960 11348 18012 11354
rect 17960 11290 18012 11296
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 17224 10464 17276 10470
rect 17224 10406 17276 10412
rect 17236 9722 17264 10406
rect 18340 10130 18368 11494
rect 18432 11354 18460 11698
rect 18524 11354 18552 11698
rect 18800 11694 18828 12038
rect 18788 11688 18840 11694
rect 18788 11630 18840 11636
rect 19352 11558 19380 12038
rect 19444 11898 19472 12174
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 20088 11626 20116 12242
rect 20272 12102 20300 12406
rect 20352 12232 20404 12238
rect 20548 12220 20576 12718
rect 20404 12192 20576 12220
rect 20352 12174 20404 12180
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 19340 11552 19392 11558
rect 20272 11540 20300 12038
rect 20364 11762 20392 12174
rect 20640 11898 20668 19110
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 17882 20760 18702
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20824 17762 20852 20334
rect 20732 17734 20852 17762
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20732 17542 20760 17734
rect 20916 17678 20944 17750
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20812 17536 20864 17542
rect 20812 17478 20864 17484
rect 20824 17270 20852 17478
rect 20812 17264 20864 17270
rect 20812 17206 20864 17212
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20824 15162 20852 16526
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20916 14600 20944 17614
rect 21008 16998 21036 21490
rect 21284 21486 21312 22034
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21284 19446 21312 20402
rect 21560 20058 21588 24618
rect 21652 23866 21680 26386
rect 22112 25906 22140 26522
rect 22388 26382 22416 26794
rect 23400 26586 23428 26794
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 21916 25832 21968 25838
rect 21916 25774 21968 25780
rect 21928 25294 21956 25774
rect 22204 25430 22232 25978
rect 22388 25770 22416 26318
rect 22664 26042 22692 26318
rect 22652 26036 22704 26042
rect 22652 25978 22704 25984
rect 23400 25906 23428 26522
rect 24320 26518 24348 26726
rect 24872 26586 24900 26930
rect 26896 26586 26924 26930
rect 24860 26580 24912 26586
rect 24860 26522 24912 26528
rect 26884 26580 26936 26586
rect 26884 26522 26936 26528
rect 24308 26512 24360 26518
rect 24308 26454 24360 26460
rect 26700 26512 26752 26518
rect 26700 26454 26752 26460
rect 26712 25974 26740 26454
rect 26700 25968 26752 25974
rect 26700 25910 26752 25916
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 22376 25764 22428 25770
rect 22376 25706 22428 25712
rect 22388 25498 22416 25706
rect 23400 25498 23428 25842
rect 26896 25702 26924 26522
rect 26884 25696 26936 25702
rect 26884 25638 26936 25644
rect 26896 25498 26924 25638
rect 22376 25492 22428 25498
rect 22376 25434 22428 25440
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 26884 25492 26936 25498
rect 26884 25434 26936 25440
rect 22192 25424 22244 25430
rect 22192 25366 22244 25372
rect 23388 25356 23440 25362
rect 23388 25298 23440 25304
rect 21916 25288 21968 25294
rect 21916 25230 21968 25236
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 23216 24954 23244 25230
rect 23204 24948 23256 24954
rect 23204 24890 23256 24896
rect 23400 24818 23428 25298
rect 23940 25288 23992 25294
rect 23940 25230 23992 25236
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 25412 25288 25464 25294
rect 25412 25230 25464 25236
rect 23952 24954 23980 25230
rect 24596 24954 24624 25230
rect 25424 24954 25452 25230
rect 23940 24948 23992 24954
rect 23940 24890 23992 24896
rect 24584 24948 24636 24954
rect 24584 24890 24636 24896
rect 25412 24948 25464 24954
rect 25412 24890 25464 24896
rect 23388 24812 23440 24818
rect 23388 24754 23440 24760
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 25228 24812 25280 24818
rect 25228 24754 25280 24760
rect 26608 24812 26660 24818
rect 26608 24754 26660 24760
rect 23952 24614 23980 24754
rect 24032 24744 24084 24750
rect 24504 24698 24532 24754
rect 24860 24744 24912 24750
rect 24084 24692 24860 24698
rect 24032 24686 24912 24692
rect 24044 24670 24900 24686
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23940 24608 23992 24614
rect 23940 24550 23992 24556
rect 23124 24274 23152 24550
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 22848 23820 23152 23848
rect 22652 23792 22704 23798
rect 22650 23760 22652 23769
rect 22704 23760 22706 23769
rect 21916 23724 21968 23730
rect 21916 23666 21968 23672
rect 22560 23724 22612 23730
rect 22848 23730 22876 23820
rect 22650 23695 22706 23704
rect 22836 23724 22888 23730
rect 22560 23666 22612 23672
rect 22836 23666 22888 23672
rect 21928 22778 21956 23666
rect 22008 23044 22060 23050
rect 22008 22986 22060 22992
rect 21916 22772 21968 22778
rect 21916 22714 21968 22720
rect 22020 22710 22048 22986
rect 22008 22704 22060 22710
rect 22008 22646 22060 22652
rect 22020 22094 22048 22646
rect 22572 22234 22600 23666
rect 23020 23656 23072 23662
rect 23020 23598 23072 23604
rect 22928 23520 22980 23526
rect 22928 23462 22980 23468
rect 22940 23186 22968 23462
rect 23032 23322 23060 23598
rect 23124 23526 23152 23820
rect 23216 23730 23244 24550
rect 23952 23866 23980 24550
rect 23940 23860 23992 23866
rect 23940 23802 23992 23808
rect 23204 23724 23256 23730
rect 23204 23666 23256 23672
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 23584 23322 23612 23598
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 23572 23316 23624 23322
rect 23572 23258 23624 23264
rect 22928 23180 22980 23186
rect 22928 23122 22980 23128
rect 23388 23180 23440 23186
rect 23388 23122 23440 23128
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22664 22574 22692 22918
rect 23308 22778 23336 22986
rect 23400 22778 23428 23122
rect 24504 23118 24532 23666
rect 24780 23594 24808 24670
rect 25044 24268 25096 24274
rect 25044 24210 25096 24216
rect 24768 23588 24820 23594
rect 24768 23530 24820 23536
rect 24780 23254 24808 23530
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24584 23044 24636 23050
rect 24584 22986 24636 22992
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 24308 22772 24360 22778
rect 24308 22714 24360 22720
rect 22652 22568 22704 22574
rect 22652 22510 22704 22516
rect 22744 22432 22796 22438
rect 22744 22374 22796 22380
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 21928 22066 22048 22094
rect 21928 22030 21956 22066
rect 22756 22030 22784 22374
rect 23308 22094 23336 22714
rect 23848 22568 23900 22574
rect 23848 22510 23900 22516
rect 23388 22500 23440 22506
rect 23388 22442 23440 22448
rect 23032 22066 23336 22094
rect 23032 22030 23060 22066
rect 23400 22030 23428 22442
rect 23664 22228 23716 22234
rect 23664 22170 23716 22176
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 23020 22024 23072 22030
rect 23020 21966 23072 21972
rect 23388 22024 23440 22030
rect 23388 21966 23440 21972
rect 21928 21554 21956 21966
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22204 21622 22232 21898
rect 22192 21616 22244 21622
rect 22192 21558 22244 21564
rect 21916 21548 21968 21554
rect 21916 21490 21968 21496
rect 23032 21146 23060 21966
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23216 21690 23244 21830
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23584 21554 23612 21830
rect 23676 21690 23704 22170
rect 23860 22094 23888 22510
rect 24320 22506 24348 22714
rect 24412 22710 24440 22986
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24308 22500 24360 22506
rect 24308 22442 24360 22448
rect 23940 22432 23992 22438
rect 23940 22374 23992 22380
rect 23952 22234 23980 22374
rect 23940 22228 23992 22234
rect 23940 22170 23992 22176
rect 23768 22066 23888 22094
rect 23768 22030 23796 22066
rect 23756 22024 23808 22030
rect 23756 21966 23808 21972
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 23768 21418 23796 21966
rect 23756 21412 23808 21418
rect 23756 21354 23808 21360
rect 23020 21140 23072 21146
rect 23020 21082 23072 21088
rect 21732 20936 21784 20942
rect 21732 20878 21784 20884
rect 21744 20534 21772 20878
rect 24596 20602 24624 22986
rect 24952 22636 25004 22642
rect 24952 22578 25004 22584
rect 24964 21554 24992 22578
rect 24952 21548 25004 21554
rect 24952 21490 25004 21496
rect 24860 21480 24912 21486
rect 24860 21422 24912 21428
rect 24872 20942 24900 21422
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 22652 20596 22704 20602
rect 22652 20538 22704 20544
rect 24584 20596 24636 20602
rect 24584 20538 24636 20544
rect 21732 20528 21784 20534
rect 21732 20470 21784 20476
rect 22468 20256 22520 20262
rect 22468 20198 22520 20204
rect 22560 20256 22612 20262
rect 22560 20198 22612 20204
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 22192 19916 22244 19922
rect 22192 19858 22244 19864
rect 22204 19514 22232 19858
rect 22376 19848 22428 19854
rect 22376 19790 22428 19796
rect 22480 19802 22508 20198
rect 22572 19990 22600 20198
rect 22560 19984 22612 19990
rect 22560 19926 22612 19932
rect 22664 19854 22692 20538
rect 24676 20460 24728 20466
rect 24676 20402 24728 20408
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23756 20256 23808 20262
rect 23756 20198 23808 20204
rect 23032 20058 23060 20198
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22652 19848 22704 19854
rect 22192 19508 22244 19514
rect 22192 19450 22244 19456
rect 21272 19440 21324 19446
rect 21272 19382 21324 19388
rect 21364 18080 21416 18086
rect 21364 18022 21416 18028
rect 21088 17740 21140 17746
rect 21088 17682 21140 17688
rect 21100 17270 21128 17682
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17264 21140 17270
rect 21088 17206 21140 17212
rect 21192 17134 21220 17614
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21284 17270 21312 17546
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 15570 21036 16390
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 21376 15026 21404 18022
rect 21456 17672 21508 17678
rect 21456 17614 21508 17620
rect 21468 17270 21496 17614
rect 21456 17264 21508 17270
rect 21456 17206 21508 17212
rect 22388 16794 22416 19790
rect 22480 19774 22600 19802
rect 22652 19790 22704 19796
rect 22572 18766 22600 19774
rect 22664 19174 22692 19790
rect 23768 19786 23796 20198
rect 23756 19780 23808 19786
rect 23756 19722 23808 19728
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 23204 19168 23256 19174
rect 23204 19110 23256 19116
rect 22560 18760 22612 18766
rect 22560 18702 22612 18708
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22572 18222 22600 18702
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22756 18426 22784 18566
rect 22848 18426 22876 18702
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22836 18420 22888 18426
rect 22836 18362 22888 18368
rect 23216 18290 23244 19110
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 22560 18216 22612 18222
rect 22560 18158 22612 18164
rect 22652 18216 22704 18222
rect 22652 18158 22704 18164
rect 22560 17536 22612 17542
rect 22560 17478 22612 17484
rect 22572 17134 22600 17478
rect 22560 17128 22612 17134
rect 22560 17070 22612 17076
rect 22376 16788 22428 16794
rect 22376 16730 22428 16736
rect 22388 16114 22416 16730
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 21456 15972 21508 15978
rect 21456 15914 21508 15920
rect 21468 15706 21496 15914
rect 21456 15700 21508 15706
rect 21456 15642 21508 15648
rect 22284 15632 22336 15638
rect 22284 15574 22336 15580
rect 21824 15156 21876 15162
rect 21824 15098 21876 15104
rect 21456 15088 21508 15094
rect 21456 15030 21508 15036
rect 21364 15020 21416 15026
rect 21364 14962 21416 14968
rect 20996 14612 21048 14618
rect 20916 14572 20996 14600
rect 20996 14554 21048 14560
rect 21376 14414 21404 14962
rect 21468 14550 21496 15030
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21836 14414 21864 15098
rect 22192 15088 22244 15094
rect 22192 15030 22244 15036
rect 21364 14408 21416 14414
rect 21364 14350 21416 14356
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 21088 14340 21140 14346
rect 21088 14282 21140 14288
rect 20996 13524 21048 13530
rect 20996 13466 21048 13472
rect 21008 12918 21036 13466
rect 21100 12986 21128 14282
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 13938 21312 14214
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21376 13326 21404 14350
rect 22204 14074 22232 15030
rect 22296 14074 22324 15574
rect 22388 15434 22416 16050
rect 22572 16046 22600 17070
rect 22664 16726 22692 18158
rect 23020 17808 23072 17814
rect 23020 17750 23072 17756
rect 22744 17672 22796 17678
rect 22744 17614 22796 17620
rect 22756 17542 22784 17614
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 23032 17338 23060 17750
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23480 17672 23532 17678
rect 23480 17614 23532 17620
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23124 17338 23152 17478
rect 23308 17338 23336 17614
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 23020 17332 23072 17338
rect 23020 17274 23072 17280
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 22940 16794 22968 17274
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22652 16720 22704 16726
rect 22652 16662 22704 16668
rect 22928 16108 22980 16114
rect 22928 16050 22980 16056
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 22560 16040 22612 16046
rect 22560 15982 22612 15988
rect 22652 15972 22704 15978
rect 22652 15914 22704 15920
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22560 15360 22612 15366
rect 22664 15348 22692 15914
rect 22940 15706 22968 16050
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22612 15320 22692 15348
rect 22560 15302 22612 15308
rect 22468 14476 22520 14482
rect 22468 14418 22520 14424
rect 22480 14074 22508 14418
rect 21640 14068 21692 14074
rect 21640 14010 21692 14016
rect 22192 14068 22244 14074
rect 22192 14010 22244 14016
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 21652 13530 21680 14010
rect 21916 13796 21968 13802
rect 21916 13738 21968 13744
rect 21928 13530 21956 13738
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 22008 13456 22060 13462
rect 22008 13398 22060 13404
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21376 12986 21404 13262
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 22020 12238 22048 13398
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 22204 12730 22232 14010
rect 22296 13938 22324 14010
rect 22572 13938 22600 15302
rect 22744 14340 22796 14346
rect 22744 14282 22796 14288
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22572 13734 22600 13874
rect 22560 13728 22612 13734
rect 22560 13670 22612 13676
rect 22572 13190 22600 13670
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 22560 13184 22612 13190
rect 22560 13126 22612 13132
rect 22572 12850 22600 13126
rect 22560 12844 22612 12850
rect 22560 12786 22612 12792
rect 21732 12232 21784 12238
rect 21732 12174 21784 12180
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20996 11824 21048 11830
rect 20996 11766 21048 11772
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20352 11552 20404 11558
rect 20272 11512 20352 11540
rect 19340 11494 19392 11500
rect 20352 11494 20404 11500
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18512 11348 18564 11354
rect 18512 11290 18564 11296
rect 19352 11082 19380 11494
rect 19340 11076 19392 11082
rect 19340 11018 19392 11024
rect 19432 11008 19484 11014
rect 19352 10956 19432 10962
rect 19352 10950 19484 10956
rect 19352 10934 19472 10950
rect 19352 10810 19380 10934
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19984 10736 20036 10742
rect 19982 10704 19984 10713
rect 20036 10704 20038 10713
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 19248 10668 19300 10674
rect 19982 10639 20038 10648
rect 19248 10610 19300 10616
rect 18708 10266 18736 10610
rect 19260 10266 19288 10610
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19996 10266 20024 10542
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 18328 10124 18380 10130
rect 18328 10066 18380 10072
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18616 9926 18644 9998
rect 20364 9926 20392 11494
rect 21008 11354 21036 11766
rect 21100 11762 21128 12038
rect 21744 11762 21772 12174
rect 22112 12170 22140 12718
rect 22204 12702 22416 12730
rect 22192 12640 22244 12646
rect 22192 12582 22244 12588
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22204 11898 22232 12582
rect 22192 11892 22244 11898
rect 22192 11834 22244 11840
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 21088 11756 21140 11762
rect 21088 11698 21140 11704
rect 21732 11756 21784 11762
rect 21732 11698 21784 11704
rect 21362 11656 21418 11665
rect 21362 11591 21364 11600
rect 21416 11591 21418 11600
rect 21364 11562 21416 11568
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20456 10674 20484 11018
rect 21008 10810 21036 11290
rect 21192 11286 21220 11494
rect 22204 11354 22232 11834
rect 22296 11558 22324 11834
rect 22284 11552 22336 11558
rect 22284 11494 22336 11500
rect 22192 11348 22244 11354
rect 22192 11290 22244 11296
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 20444 10668 20496 10674
rect 20444 10610 20496 10616
rect 21192 10606 21220 11222
rect 22008 11144 22060 11150
rect 22008 11086 22060 11092
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21272 10600 21324 10606
rect 21272 10542 21324 10548
rect 20536 10464 20588 10470
rect 20536 10406 20588 10412
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20548 10266 20576 10406
rect 20824 10266 20852 10406
rect 21284 10266 21312 10542
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 9926 21404 10610
rect 22020 10266 22048 11086
rect 22112 10810 22140 11222
rect 22388 11150 22416 12702
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22480 11694 22508 12174
rect 22468 11688 22520 11694
rect 22468 11630 22520 11636
rect 22284 11144 22336 11150
rect 22284 11086 22336 11092
rect 22376 11144 22428 11150
rect 22376 11086 22428 11092
rect 22100 10804 22152 10810
rect 22152 10764 22232 10792
rect 22100 10746 22152 10752
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22020 10062 22048 10202
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 20352 9920 20404 9926
rect 20352 9862 20404 9868
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 18616 9654 18644 9862
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 22020 9674 22048 9998
rect 22020 9654 22140 9674
rect 18604 9648 18656 9654
rect 22020 9648 22152 9654
rect 22020 9646 22100 9648
rect 18604 9590 18656 9596
rect 22100 9590 22152 9596
rect 22204 9586 22232 10764
rect 22296 10470 22324 11086
rect 22480 10606 22508 11630
rect 22572 11354 22600 12786
rect 22664 12646 22692 13466
rect 22756 12986 22784 14282
rect 23124 14074 23152 16050
rect 23296 15428 23348 15434
rect 23296 15370 23348 15376
rect 23308 15026 23336 15370
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23388 14408 23440 14414
rect 23388 14350 23440 14356
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23124 13530 23152 14010
rect 23400 13734 23428 14350
rect 23492 14278 23520 17614
rect 23584 16794 23612 19450
rect 23664 18692 23716 18698
rect 23664 18634 23716 18640
rect 23676 17610 23704 18634
rect 23768 17678 23796 19722
rect 24688 19310 24716 20402
rect 24872 20330 24900 20878
rect 24964 20602 24992 21490
rect 25056 20942 25084 24210
rect 25240 23254 25268 24754
rect 26240 23724 26292 23730
rect 26240 23666 26292 23672
rect 26148 23656 26200 23662
rect 26148 23598 26200 23604
rect 25228 23248 25280 23254
rect 25228 23190 25280 23196
rect 26160 23118 26188 23598
rect 26252 23322 26280 23666
rect 26240 23316 26292 23322
rect 26240 23258 26292 23264
rect 25136 23112 25188 23118
rect 25136 23054 25188 23060
rect 26056 23112 26108 23118
rect 26056 23054 26108 23060
rect 26148 23112 26200 23118
rect 26148 23054 26200 23060
rect 25148 21010 25176 23054
rect 25320 22976 25372 22982
rect 25320 22918 25372 22924
rect 25332 22642 25360 22918
rect 25320 22636 25372 22642
rect 25320 22578 25372 22584
rect 25872 22568 25924 22574
rect 25872 22510 25924 22516
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25884 20942 25912 22510
rect 26068 22506 26096 23054
rect 26056 22500 26108 22506
rect 26056 22442 26108 22448
rect 26160 22166 26188 23054
rect 26148 22160 26200 22166
rect 26148 22102 26200 22108
rect 26424 21548 26476 21554
rect 26424 21490 26476 21496
rect 26436 21146 26464 21490
rect 26424 21140 26476 21146
rect 26424 21082 26476 21088
rect 25044 20936 25096 20942
rect 25044 20878 25096 20884
rect 25504 20936 25556 20942
rect 25504 20878 25556 20884
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 24952 20596 25004 20602
rect 24952 20538 25004 20544
rect 25136 20460 25188 20466
rect 25136 20402 25188 20408
rect 24860 20324 24912 20330
rect 24860 20266 24912 20272
rect 24872 19922 24900 20266
rect 25148 20058 25176 20402
rect 25136 20052 25188 20058
rect 25136 19994 25188 20000
rect 24860 19916 24912 19922
rect 24860 19858 24912 19864
rect 25320 19780 25372 19786
rect 25320 19722 25372 19728
rect 25228 19712 25280 19718
rect 25228 19654 25280 19660
rect 25240 19394 25268 19654
rect 25332 19514 25360 19722
rect 25516 19514 25544 20878
rect 25792 20466 25820 20878
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25596 20324 25648 20330
rect 25596 20266 25648 20272
rect 25608 19854 25636 20266
rect 25792 19922 25820 20402
rect 25884 20058 25912 20878
rect 26332 20868 26384 20874
rect 26332 20810 26384 20816
rect 26344 20466 26372 20810
rect 26332 20460 26384 20466
rect 26332 20402 26384 20408
rect 26516 20256 26568 20262
rect 26516 20198 26568 20204
rect 26528 20058 26556 20198
rect 25872 20052 25924 20058
rect 25872 19994 25924 20000
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 25780 19916 25832 19922
rect 25780 19858 25832 19864
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25608 19718 25636 19790
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25320 19508 25372 19514
rect 25320 19450 25372 19456
rect 25504 19508 25556 19514
rect 25504 19450 25556 19456
rect 25240 19378 25360 19394
rect 25608 19378 25636 19654
rect 25240 19372 25372 19378
rect 25240 19366 25320 19372
rect 25320 19314 25372 19320
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 24676 19304 24728 19310
rect 24676 19246 24728 19252
rect 25332 18970 25360 19314
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23664 17604 23716 17610
rect 23664 17546 23716 17552
rect 25884 17338 25912 18566
rect 25872 17332 25924 17338
rect 25872 17274 25924 17280
rect 25228 17196 25280 17202
rect 25228 17138 25280 17144
rect 25412 17196 25464 17202
rect 25412 17138 25464 17144
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 25136 17128 25188 17134
rect 25136 17070 25188 17076
rect 23572 16788 23624 16794
rect 23572 16730 23624 16736
rect 23584 16658 23612 16730
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 23676 15502 23704 16594
rect 23756 16584 23808 16590
rect 23756 16526 23808 16532
rect 24768 16584 24820 16590
rect 24768 16526 24820 16532
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 23768 15502 23796 16526
rect 24780 16114 24808 16526
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 24768 16108 24820 16114
rect 24768 16050 24820 16056
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23952 15502 23980 15846
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23756 15496 23808 15502
rect 23756 15438 23808 15444
rect 23940 15496 23992 15502
rect 23940 15438 23992 15444
rect 23768 15162 23796 15438
rect 23756 15156 23808 15162
rect 23756 15098 23808 15104
rect 23480 14272 23532 14278
rect 23480 14214 23532 14220
rect 23952 13938 23980 15438
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 23940 13932 23992 13938
rect 23940 13874 23992 13880
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23388 13728 23440 13734
rect 23388 13670 23440 13676
rect 23676 13530 23704 13806
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23664 13524 23716 13530
rect 23664 13466 23716 13472
rect 23572 13320 23624 13326
rect 23572 13262 23624 13268
rect 23296 13184 23348 13190
rect 23296 13126 23348 13132
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 23204 12980 23256 12986
rect 23204 12922 23256 12928
rect 22836 12708 22888 12714
rect 22836 12650 22888 12656
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22560 11348 22612 11354
rect 22560 11290 22612 11296
rect 22664 11082 22692 12582
rect 22848 12442 22876 12650
rect 22836 12436 22888 12442
rect 22836 12378 22888 12384
rect 23216 12238 23244 12922
rect 23308 12442 23336 13126
rect 23388 12640 23440 12646
rect 23388 12582 23440 12588
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23400 12442 23428 12582
rect 23296 12436 23348 12442
rect 23296 12378 23348 12384
rect 23388 12436 23440 12442
rect 23388 12378 23440 12384
rect 22744 12232 22796 12238
rect 23204 12232 23256 12238
rect 22744 12174 22796 12180
rect 22834 12200 22890 12209
rect 22756 11558 22784 12174
rect 23204 12174 23256 12180
rect 22834 12135 22890 12144
rect 22848 12102 22876 12135
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22928 12096 22980 12102
rect 22928 12038 22980 12044
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22744 11552 22796 11558
rect 22744 11494 22796 11500
rect 22848 11286 22876 11630
rect 22940 11626 22968 12038
rect 23216 11898 23244 12174
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 22928 11620 22980 11626
rect 22928 11562 22980 11568
rect 23308 11558 23336 12378
rect 23388 12232 23440 12238
rect 23492 12220 23520 12582
rect 23440 12192 23520 12220
rect 23388 12174 23440 12180
rect 23584 12102 23612 13262
rect 23676 12850 23704 13466
rect 23952 13258 23980 13874
rect 23940 13252 23992 13258
rect 23940 13194 23992 13200
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 23676 12186 23704 12786
rect 23848 12300 23900 12306
rect 23848 12242 23900 12248
rect 23860 12186 23888 12242
rect 23676 12158 23888 12186
rect 23860 12102 23888 12158
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23848 12096 23900 12102
rect 23848 12038 23900 12044
rect 23940 12096 23992 12102
rect 23940 12038 23992 12044
rect 23584 11898 23612 12038
rect 23572 11892 23624 11898
rect 23624 11852 23704 11880
rect 23572 11834 23624 11840
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 22836 11280 22888 11286
rect 22756 11240 22836 11268
rect 22652 11076 22704 11082
rect 22652 11018 22704 11024
rect 22664 10742 22692 11018
rect 22652 10736 22704 10742
rect 22652 10678 22704 10684
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22284 10464 22336 10470
rect 22284 10406 22336 10412
rect 22572 10130 22600 10610
rect 22756 10538 22784 11240
rect 22836 11222 22888 11228
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 22744 10532 22796 10538
rect 22744 10474 22796 10480
rect 22848 10266 22876 11086
rect 23020 10668 23072 10674
rect 23020 10610 23072 10616
rect 23032 10266 23060 10610
rect 22836 10260 22888 10266
rect 22836 10202 22888 10208
rect 23020 10260 23072 10266
rect 23020 10202 23072 10208
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 22468 10056 22520 10062
rect 22468 9998 22520 10004
rect 22480 9654 22508 9998
rect 22848 9926 22876 10202
rect 22836 9920 22888 9926
rect 22836 9862 22888 9868
rect 22928 9920 22980 9926
rect 22928 9862 22980 9868
rect 22940 9722 22968 9862
rect 23032 9722 23060 10202
rect 22928 9716 22980 9722
rect 22928 9658 22980 9664
rect 23020 9716 23072 9722
rect 23020 9658 23072 9664
rect 23308 9654 23336 11494
rect 23676 11150 23704 11852
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23584 10674 23612 11018
rect 23572 10668 23624 10674
rect 23572 10610 23624 10616
rect 23584 10130 23612 10610
rect 23676 10606 23704 11086
rect 23860 10810 23888 12038
rect 23952 11830 23980 12038
rect 23940 11824 23992 11830
rect 23940 11766 23992 11772
rect 23952 11354 23980 11766
rect 23940 11348 23992 11354
rect 23940 11290 23992 11296
rect 24044 11150 24072 14962
rect 24136 14006 24164 16050
rect 24676 14272 24728 14278
rect 24676 14214 24728 14220
rect 24124 14000 24176 14006
rect 24124 13942 24176 13948
rect 24688 13938 24716 14214
rect 24964 14074 24992 16526
rect 25056 15026 25084 17070
rect 25148 16250 25176 17070
rect 25240 16794 25268 17138
rect 25228 16788 25280 16794
rect 25228 16730 25280 16736
rect 25424 16658 25452 17138
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25608 16658 25636 16934
rect 25412 16652 25464 16658
rect 25412 16594 25464 16600
rect 25596 16652 25648 16658
rect 25596 16594 25648 16600
rect 25136 16244 25188 16250
rect 25136 16186 25188 16192
rect 25424 15910 25452 16594
rect 25884 16590 25912 17070
rect 25964 16992 26016 16998
rect 25964 16934 26016 16940
rect 26240 16992 26292 16998
rect 26240 16934 26292 16940
rect 25872 16584 25924 16590
rect 25872 16526 25924 16532
rect 25976 16114 26004 16934
rect 26252 16794 26280 16934
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 25964 16108 26016 16114
rect 25964 16050 26016 16056
rect 25412 15904 25464 15910
rect 25412 15846 25464 15852
rect 25596 15428 25648 15434
rect 25596 15370 25648 15376
rect 25136 15088 25188 15094
rect 25136 15030 25188 15036
rect 25044 15020 25096 15026
rect 25044 14962 25096 14968
rect 25044 14612 25096 14618
rect 25044 14554 25096 14560
rect 24952 14068 25004 14074
rect 24952 14010 25004 14016
rect 25056 14006 25084 14554
rect 25148 14414 25176 15030
rect 25504 15020 25556 15026
rect 25504 14962 25556 14968
rect 25412 14884 25464 14890
rect 25412 14826 25464 14832
rect 25424 14618 25452 14826
rect 25412 14612 25464 14618
rect 25412 14554 25464 14560
rect 25516 14482 25544 14962
rect 25608 14890 25636 15370
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 26068 15026 26096 15302
rect 26160 15162 26188 16526
rect 26240 15360 26292 15366
rect 26240 15302 26292 15308
rect 26148 15156 26200 15162
rect 26148 15098 26200 15104
rect 26056 15020 26108 15026
rect 26056 14962 26108 14968
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 25596 14884 25648 14890
rect 25596 14826 25648 14832
rect 25504 14476 25556 14482
rect 25504 14418 25556 14424
rect 25608 14414 25636 14826
rect 25688 14816 25740 14822
rect 25688 14758 25740 14764
rect 25700 14550 25728 14758
rect 25688 14544 25740 14550
rect 25688 14486 25740 14492
rect 25136 14408 25188 14414
rect 25136 14350 25188 14356
rect 25596 14408 25648 14414
rect 25596 14350 25648 14356
rect 25044 14000 25096 14006
rect 25044 13942 25096 13948
rect 24676 13932 24728 13938
rect 24676 13874 24728 13880
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24504 13462 24532 13806
rect 24492 13456 24544 13462
rect 24492 13398 24544 13404
rect 24504 12850 24532 13398
rect 25056 12850 25084 13942
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 25044 12844 25096 12850
rect 25044 12786 25096 12792
rect 25056 12434 25084 12786
rect 25148 12782 25176 14350
rect 25228 14272 25280 14278
rect 25228 14214 25280 14220
rect 25240 13734 25268 14214
rect 25700 14074 25728 14486
rect 26160 14482 26188 14894
rect 26252 14890 26280 15302
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26344 14906 26372 14962
rect 26240 14884 26292 14890
rect 26344 14878 26464 14906
rect 26240 14826 26292 14832
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26148 14476 26200 14482
rect 26148 14418 26200 14424
rect 26056 14408 26108 14414
rect 26344 14362 26372 14758
rect 26436 14414 26464 14878
rect 26108 14356 26372 14362
rect 26056 14350 26372 14356
rect 26424 14408 26476 14414
rect 26424 14350 26476 14356
rect 26068 14334 26372 14350
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25240 12986 25268 13670
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25136 12776 25188 12782
rect 25136 12718 25188 12724
rect 25240 12442 25268 12922
rect 25872 12776 25924 12782
rect 25872 12718 25924 12724
rect 25228 12436 25280 12442
rect 25056 12406 25176 12434
rect 24216 12164 24268 12170
rect 24216 12106 24268 12112
rect 24228 11354 24256 12106
rect 24768 11892 24820 11898
rect 24768 11834 24820 11840
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 24676 11280 24728 11286
rect 24676 11222 24728 11228
rect 24032 11144 24084 11150
rect 24032 11086 24084 11092
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24492 11144 24544 11150
rect 24492 11086 24544 11092
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23676 10062 23704 10542
rect 24044 10266 24072 11086
rect 24412 10742 24440 11086
rect 24504 10742 24532 11086
rect 24688 11082 24716 11222
rect 24780 11150 24808 11834
rect 24768 11144 24820 11150
rect 24768 11086 24820 11092
rect 24676 11076 24728 11082
rect 24676 11018 24728 11024
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24492 10736 24544 10742
rect 24492 10678 24544 10684
rect 24216 10600 24268 10606
rect 24216 10542 24268 10548
rect 24228 10266 24256 10542
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24216 10260 24268 10266
rect 24216 10202 24268 10208
rect 24044 10146 24072 10202
rect 23952 10118 24072 10146
rect 24412 10146 24440 10678
rect 24688 10674 24716 11018
rect 24676 10668 24728 10674
rect 24676 10610 24728 10616
rect 25044 10668 25096 10674
rect 25044 10610 25096 10616
rect 25056 10470 25084 10610
rect 25044 10464 25096 10470
rect 25044 10406 25096 10412
rect 24412 10118 24532 10146
rect 23664 10056 23716 10062
rect 23664 9998 23716 10004
rect 23952 9994 23980 10118
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24124 10056 24176 10062
rect 24124 9998 24176 10004
rect 23940 9988 23992 9994
rect 23940 9930 23992 9936
rect 22468 9648 22520 9654
rect 22468 9590 22520 9596
rect 23296 9648 23348 9654
rect 23296 9590 23348 9596
rect 23952 9586 23980 9930
rect 24044 9722 24072 9998
rect 24136 9722 24164 9998
rect 24504 9994 24532 10118
rect 25044 10056 25096 10062
rect 25044 9998 25096 10004
rect 24492 9988 24544 9994
rect 24492 9930 24544 9936
rect 24308 9920 24360 9926
rect 24308 9862 24360 9868
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24044 9586 24072 9658
rect 24320 9654 24348 9862
rect 24308 9648 24360 9654
rect 24308 9590 24360 9596
rect 22192 9580 22244 9586
rect 22192 9522 22244 9528
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23032 9178 23060 9522
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23020 9172 23072 9178
rect 23020 9114 23072 9120
rect 10048 9104 10100 9110
rect 10048 9046 10100 9052
rect 23768 8974 23796 9318
rect 23952 9178 23980 9522
rect 23940 9172 23992 9178
rect 23940 9114 23992 9120
rect 25056 8974 25084 9998
rect 25148 9994 25176 12406
rect 25228 12378 25280 12384
rect 25884 12374 25912 12718
rect 26056 12640 26108 12646
rect 26056 12582 26108 12588
rect 25872 12368 25924 12374
rect 25872 12310 25924 12316
rect 26068 12238 26096 12582
rect 26252 12434 26280 14334
rect 26252 12406 26372 12434
rect 25688 12232 25740 12238
rect 26056 12232 26108 12238
rect 25688 12174 25740 12180
rect 25976 12192 26056 12220
rect 25320 12164 25372 12170
rect 25320 12106 25372 12112
rect 25332 11694 25360 12106
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25332 11354 25360 11630
rect 25700 11558 25728 12174
rect 25976 11762 26004 12192
rect 26056 12174 26108 12180
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25688 11552 25740 11558
rect 25688 11494 25740 11500
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25516 10810 25544 11086
rect 25504 10804 25556 10810
rect 25504 10746 25556 10752
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25792 10713 25820 10746
rect 25778 10704 25834 10713
rect 25976 10674 26004 11698
rect 25778 10639 25834 10648
rect 25964 10668 26016 10674
rect 25228 10600 25280 10606
rect 25228 10542 25280 10548
rect 25240 10266 25268 10542
rect 25228 10260 25280 10266
rect 25228 10202 25280 10208
rect 25792 10062 25820 10639
rect 25964 10610 26016 10616
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25976 9926 26004 10610
rect 26344 10538 26372 12406
rect 26516 11892 26568 11898
rect 26516 11834 26568 11840
rect 26528 10742 26556 11834
rect 26516 10736 26568 10742
rect 26516 10678 26568 10684
rect 26332 10532 26384 10538
rect 26332 10474 26384 10480
rect 26148 10260 26200 10266
rect 26148 10202 26200 10208
rect 26160 9994 26188 10202
rect 26148 9988 26200 9994
rect 26148 9930 26200 9936
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 23756 8968 23808 8974
rect 23756 8910 23808 8916
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25976 8906 26004 9862
rect 26620 9722 26648 24754
rect 27080 24274 27108 27066
rect 30024 26790 30052 27270
rect 28908 26784 28960 26790
rect 28908 26726 28960 26732
rect 29920 26784 29972 26790
rect 29920 26726 29972 26732
rect 30012 26784 30064 26790
rect 30012 26726 30064 26732
rect 28920 26382 28948 26726
rect 28908 26376 28960 26382
rect 28908 26318 28960 26324
rect 29932 25906 29960 26726
rect 30024 26586 30052 26726
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 30472 26308 30524 26314
rect 30472 26250 30524 26256
rect 30564 26308 30616 26314
rect 30564 26250 30616 26256
rect 30484 25922 30512 26250
rect 30576 26042 30604 26250
rect 30760 26246 30788 27390
rect 30840 27328 30892 27334
rect 30840 27270 30892 27276
rect 30852 27130 30880 27270
rect 30840 27124 30892 27130
rect 30840 27066 30892 27072
rect 30944 26926 30972 27814
rect 31036 27470 31064 27814
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 30932 26920 30984 26926
rect 30932 26862 30984 26868
rect 31036 26586 31064 27406
rect 31772 27402 31800 27814
rect 31208 27396 31260 27402
rect 31208 27338 31260 27344
rect 31760 27396 31812 27402
rect 31760 27338 31812 27344
rect 31220 26994 31248 27338
rect 31208 26988 31260 26994
rect 31208 26930 31260 26936
rect 31024 26580 31076 26586
rect 31024 26522 31076 26528
rect 32600 26382 32628 27814
rect 32968 27130 32996 27950
rect 32956 27124 33008 27130
rect 32956 27066 33008 27072
rect 33060 26790 33088 28426
rect 33152 27606 33180 36110
rect 34336 36100 34388 36106
rect 34336 36042 34388 36048
rect 34348 35737 34376 36042
rect 34334 35728 34390 35737
rect 34334 35663 34390 35672
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34520 33992 34572 33998
rect 34520 33934 34572 33940
rect 34428 31816 34480 31822
rect 34428 31758 34480 31764
rect 34060 31748 34112 31754
rect 34060 31690 34112 31696
rect 34072 31385 34100 31690
rect 34058 31376 34114 31385
rect 34058 31311 34114 31320
rect 34152 28552 34204 28558
rect 34152 28494 34204 28500
rect 33692 28144 33744 28150
rect 33692 28086 33744 28092
rect 33704 27674 33732 28086
rect 34164 27674 34192 28494
rect 34440 28218 34468 31758
rect 34532 28762 34560 33934
rect 34612 33924 34664 33930
rect 34612 33866 34664 33872
rect 34624 33561 34652 33866
rect 34610 33552 34666 33561
rect 34610 33487 34666 33496
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34612 29572 34664 29578
rect 34612 29514 34664 29520
rect 34624 29209 34652 29514
rect 34796 29504 34848 29510
rect 34796 29446 34848 29452
rect 34610 29200 34666 29209
rect 34610 29135 34666 29144
rect 34520 28756 34572 28762
rect 34520 28698 34572 28704
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34704 27872 34756 27878
rect 34704 27814 34756 27820
rect 33692 27668 33744 27674
rect 33692 27610 33744 27616
rect 34152 27668 34204 27674
rect 34152 27610 34204 27616
rect 33140 27600 33192 27606
rect 33140 27542 33192 27548
rect 34716 27538 34744 27814
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 33416 27464 33468 27470
rect 33416 27406 33468 27412
rect 34152 27464 34204 27470
rect 34152 27406 34204 27412
rect 33428 27130 33456 27406
rect 33416 27124 33468 27130
rect 33416 27066 33468 27072
rect 33692 26988 33744 26994
rect 33692 26930 33744 26936
rect 33048 26784 33100 26790
rect 33048 26726 33100 26732
rect 32588 26376 32640 26382
rect 32588 26318 32640 26324
rect 33048 26308 33100 26314
rect 33048 26250 33100 26256
rect 30748 26240 30800 26246
rect 30748 26182 30800 26188
rect 31576 26240 31628 26246
rect 31576 26182 31628 26188
rect 32128 26240 32180 26246
rect 32128 26182 32180 26188
rect 30564 26036 30616 26042
rect 30564 25978 30616 25984
rect 30656 25968 30708 25974
rect 30484 25916 30656 25922
rect 30484 25910 30708 25916
rect 29920 25900 29972 25906
rect 29920 25842 29972 25848
rect 30484 25894 30696 25910
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 30104 25696 30156 25702
rect 30104 25638 30156 25644
rect 27344 24608 27396 24614
rect 27344 24550 27396 24556
rect 27356 24410 27384 24550
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 27068 24268 27120 24274
rect 27068 24210 27120 24216
rect 26884 23860 26936 23866
rect 26884 23802 26936 23808
rect 26700 23656 26752 23662
rect 26700 23598 26752 23604
rect 26712 23322 26740 23598
rect 26700 23316 26752 23322
rect 26700 23258 26752 23264
rect 26896 23118 26924 23802
rect 27724 23730 27752 25638
rect 27804 25220 27856 25226
rect 27804 25162 27856 25168
rect 27816 24410 27844 25162
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 30116 24274 30144 25638
rect 30484 24954 30512 25894
rect 31588 25702 31616 26182
rect 32140 25838 32168 26182
rect 33060 26042 33088 26250
rect 33704 26042 33732 26930
rect 33048 26036 33100 26042
rect 33048 25978 33100 25984
rect 33692 26036 33744 26042
rect 33692 25978 33744 25984
rect 34164 25906 34192 27406
rect 34702 27024 34758 27033
rect 34702 26959 34704 26968
rect 34756 26959 34758 26968
rect 34704 26930 34756 26936
rect 34808 26586 34836 29446
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 34336 26308 34388 26314
rect 34336 26250 34388 26256
rect 34348 26042 34376 26250
rect 34336 26036 34388 26042
rect 34336 25978 34388 25984
rect 34152 25900 34204 25906
rect 34152 25842 34204 25848
rect 32128 25832 32180 25838
rect 32128 25774 32180 25780
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 31576 25696 31628 25702
rect 31576 25638 31628 25644
rect 30932 25356 30984 25362
rect 30932 25298 30984 25304
rect 30840 25288 30892 25294
rect 30840 25230 30892 25236
rect 30472 24948 30524 24954
rect 30472 24890 30524 24896
rect 30852 24614 30880 25230
rect 30944 24954 30972 25298
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 31588 24750 31616 25638
rect 32140 25158 32168 25774
rect 32416 25498 32444 25774
rect 32404 25492 32456 25498
rect 32404 25434 32456 25440
rect 34060 25220 34112 25226
rect 34060 25162 34112 25168
rect 32128 25152 32180 25158
rect 32128 25094 32180 25100
rect 32404 25152 32456 25158
rect 32404 25094 32456 25100
rect 31576 24744 31628 24750
rect 31576 24686 31628 24692
rect 31588 24614 31616 24686
rect 32416 24614 32444 25094
rect 34072 24857 34100 25162
rect 34058 24848 34114 24857
rect 33784 24812 33836 24818
rect 34058 24783 34114 24792
rect 33784 24754 33836 24760
rect 32680 24744 32732 24750
rect 32680 24686 32732 24692
rect 30656 24608 30708 24614
rect 30656 24550 30708 24556
rect 30840 24608 30892 24614
rect 30840 24550 30892 24556
rect 31576 24608 31628 24614
rect 31576 24550 31628 24556
rect 31668 24608 31720 24614
rect 31668 24550 31720 24556
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 30104 24268 30156 24274
rect 30104 24210 30156 24216
rect 29552 24064 29604 24070
rect 29552 24006 29604 24012
rect 29564 23866 29592 24006
rect 29552 23860 29604 23866
rect 29552 23802 29604 23808
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27724 23322 27752 23666
rect 30116 23526 30144 24210
rect 30668 24206 30696 24550
rect 30656 24200 30708 24206
rect 30656 24142 30708 24148
rect 31588 24070 31616 24550
rect 31680 24138 31708 24550
rect 31668 24132 31720 24138
rect 31668 24074 31720 24080
rect 31576 24064 31628 24070
rect 31576 24006 31628 24012
rect 30104 23520 30156 23526
rect 30104 23462 30156 23468
rect 27712 23316 27764 23322
rect 27712 23258 27764 23264
rect 28356 23316 28408 23322
rect 28356 23258 28408 23264
rect 26884 23112 26936 23118
rect 26884 23054 26936 23060
rect 28368 21622 28396 23258
rect 28356 21616 28408 21622
rect 28356 21558 28408 21564
rect 27160 19984 27212 19990
rect 27160 19926 27212 19932
rect 27172 19854 27200 19926
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26804 18970 26832 19654
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 27172 18902 27200 19790
rect 27712 19712 27764 19718
rect 27712 19654 27764 19660
rect 27724 19446 27752 19654
rect 28368 19514 28396 21558
rect 30116 21554 30144 23462
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30300 21690 30328 21830
rect 31128 21690 31156 22034
rect 31588 21690 31616 24006
rect 31680 22098 31708 24074
rect 31668 22092 31720 22098
rect 31668 22034 31720 22040
rect 32312 22092 32364 22098
rect 32416 22080 32444 24550
rect 32692 24410 32720 24686
rect 33324 24608 33376 24614
rect 33324 24550 33376 24556
rect 32680 24404 32732 24410
rect 32680 24346 32732 24352
rect 33336 24342 33364 24550
rect 33796 24410 33824 24754
rect 34164 24614 34192 25842
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34348 24954 34376 25230
rect 34336 24948 34388 24954
rect 34336 24890 34388 24896
rect 34152 24608 34204 24614
rect 34152 24550 34204 24556
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33784 24404 33836 24410
rect 33784 24346 33836 24352
rect 33140 24336 33192 24342
rect 33140 24278 33192 24284
rect 33324 24336 33376 24342
rect 33324 24278 33376 24284
rect 32364 22052 32444 22080
rect 32312 22034 32364 22040
rect 32036 21956 32088 21962
rect 32036 21898 32088 21904
rect 30288 21684 30340 21690
rect 30288 21626 30340 21632
rect 31116 21684 31168 21690
rect 31116 21626 31168 21632
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 32048 21554 32076 21898
rect 30104 21548 30156 21554
rect 30104 21490 30156 21496
rect 31024 21548 31076 21554
rect 31024 21490 31076 21496
rect 32036 21548 32088 21554
rect 32036 21490 32088 21496
rect 30116 20058 30144 21490
rect 30104 20052 30156 20058
rect 30104 19994 30156 20000
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 28356 19508 28408 19514
rect 28356 19450 28408 19456
rect 27712 19440 27764 19446
rect 27712 19382 27764 19388
rect 28368 19378 28396 19450
rect 29748 19446 29776 19654
rect 29736 19440 29788 19446
rect 29736 19382 29788 19388
rect 28356 19372 28408 19378
rect 28356 19314 28408 19320
rect 27160 18896 27212 18902
rect 27160 18838 27212 18844
rect 28724 18760 28776 18766
rect 28724 18702 28776 18708
rect 29368 18760 29420 18766
rect 29368 18702 29420 18708
rect 27160 18692 27212 18698
rect 27160 18634 27212 18640
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 27172 18290 27200 18634
rect 27160 18284 27212 18290
rect 27160 18226 27212 18232
rect 27540 17882 27568 18634
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27724 17882 27752 18566
rect 27896 18284 27948 18290
rect 27896 18226 27948 18232
rect 27528 17876 27580 17882
rect 27528 17818 27580 17824
rect 27712 17876 27764 17882
rect 27712 17818 27764 17824
rect 27528 17672 27580 17678
rect 27528 17614 27580 17620
rect 27436 17604 27488 17610
rect 27436 17546 27488 17552
rect 26976 17536 27028 17542
rect 26976 17478 27028 17484
rect 26988 15706 27016 17478
rect 27448 17134 27476 17546
rect 27540 17202 27568 17614
rect 27908 17610 27936 18226
rect 28736 17746 28764 18702
rect 28908 18624 28960 18630
rect 28908 18566 28960 18572
rect 28816 17808 28868 17814
rect 28816 17750 28868 17756
rect 28724 17740 28776 17746
rect 28724 17682 28776 17688
rect 28184 17610 28580 17626
rect 27896 17604 27948 17610
rect 27896 17546 27948 17552
rect 28172 17604 28580 17610
rect 28224 17598 28580 17604
rect 28172 17546 28224 17552
rect 27620 17536 27672 17542
rect 27620 17478 27672 17484
rect 27804 17536 27856 17542
rect 27804 17478 27856 17484
rect 27632 17338 27660 17478
rect 27816 17338 27844 17478
rect 27620 17332 27672 17338
rect 27620 17274 27672 17280
rect 27804 17332 27856 17338
rect 27804 17274 27856 17280
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27816 16250 27844 17138
rect 27804 16244 27856 16250
rect 27804 16186 27856 16192
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 27080 15366 27108 16050
rect 27172 15502 27200 16050
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 27068 15360 27120 15366
rect 27068 15302 27120 15308
rect 27080 15026 27108 15302
rect 27068 15020 27120 15026
rect 27068 14962 27120 14968
rect 27172 14958 27200 15438
rect 27540 15434 27568 16050
rect 27908 15502 27936 17546
rect 28552 17542 28580 17598
rect 28448 17536 28500 17542
rect 28448 17478 28500 17484
rect 28540 17536 28592 17542
rect 28540 17478 28592 17484
rect 28460 17338 28488 17478
rect 28828 17338 28856 17750
rect 28920 17610 28948 18566
rect 28908 17604 28960 17610
rect 28908 17546 28960 17552
rect 29380 17338 29408 18702
rect 30116 18426 30144 19994
rect 30196 19712 30248 19718
rect 30196 19654 30248 19660
rect 30208 19514 30236 19654
rect 30196 19508 30248 19514
rect 30196 19450 30248 19456
rect 31036 19310 31064 21490
rect 32048 20058 32076 21490
rect 32416 21350 32444 22052
rect 33152 21350 33180 24278
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34336 23112 34388 23118
rect 34336 23054 34388 23060
rect 34348 22234 34376 23054
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34624 22681 34652 22986
rect 34610 22672 34666 22681
rect 34610 22607 34666 22616
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34336 22228 34388 22234
rect 34336 22170 34388 22176
rect 33324 21956 33376 21962
rect 33324 21898 33376 21904
rect 33336 21690 33364 21898
rect 33324 21684 33376 21690
rect 33324 21626 33376 21632
rect 32404 21344 32456 21350
rect 32404 21286 32456 21292
rect 32680 21344 32732 21350
rect 32680 21286 32732 21292
rect 33140 21344 33192 21350
rect 33140 21286 33192 21292
rect 32496 20392 32548 20398
rect 32496 20334 32548 20340
rect 32508 20058 32536 20334
rect 32692 20262 32720 21286
rect 32680 20256 32732 20262
rect 32732 20204 32812 20210
rect 32680 20198 32812 20204
rect 32692 20182 32812 20198
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 32496 20052 32548 20058
rect 32496 19994 32548 20000
rect 31116 19916 31168 19922
rect 31116 19858 31168 19864
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31128 19514 31156 19858
rect 31116 19508 31168 19514
rect 31116 19450 31168 19456
rect 31404 19446 31432 19858
rect 31484 19712 31536 19718
rect 31484 19654 31536 19660
rect 31392 19440 31444 19446
rect 31392 19382 31444 19388
rect 31024 19304 31076 19310
rect 31024 19246 31076 19252
rect 31404 18970 31432 19382
rect 31496 19174 31524 19654
rect 32220 19236 32272 19242
rect 32220 19178 32272 19184
rect 31484 19168 31536 19174
rect 31484 19110 31536 19116
rect 31392 18964 31444 18970
rect 31392 18906 31444 18912
rect 31496 18698 31524 19110
rect 32232 18766 32260 19178
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 31484 18692 31536 18698
rect 31484 18634 31536 18640
rect 30300 18426 30328 18634
rect 30104 18420 30156 18426
rect 30104 18362 30156 18368
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 28448 17332 28500 17338
rect 28448 17274 28500 17280
rect 28816 17332 28868 17338
rect 28816 17274 28868 17280
rect 29368 17332 29420 17338
rect 29368 17274 29420 17280
rect 28356 15904 28408 15910
rect 28356 15846 28408 15852
rect 28368 15570 28396 15846
rect 28080 15564 28132 15570
rect 28080 15506 28132 15512
rect 28356 15564 28408 15570
rect 28356 15506 28408 15512
rect 27896 15496 27948 15502
rect 27896 15438 27948 15444
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27160 14952 27212 14958
rect 27160 14894 27212 14900
rect 27172 14482 27200 14894
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27264 13530 27292 15370
rect 27988 15360 28040 15366
rect 27988 15302 28040 15308
rect 28000 15026 28028 15302
rect 28092 15162 28120 15506
rect 28356 15428 28408 15434
rect 28356 15370 28408 15376
rect 28724 15428 28776 15434
rect 28724 15370 28776 15376
rect 28368 15162 28396 15370
rect 28736 15162 28764 15370
rect 29380 15162 29408 17274
rect 30116 16794 30144 18362
rect 31496 17338 31524 18634
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31956 18426 31984 18566
rect 31944 18420 31996 18426
rect 31944 18362 31996 18368
rect 31484 17332 31536 17338
rect 31484 17274 31536 17280
rect 30380 17264 30432 17270
rect 30380 17206 30432 17212
rect 30392 16794 30420 17206
rect 31760 17196 31812 17202
rect 31760 17138 31812 17144
rect 31944 17196 31996 17202
rect 31944 17138 31996 17144
rect 30104 16788 30156 16794
rect 30104 16730 30156 16736
rect 30380 16788 30432 16794
rect 30380 16730 30432 16736
rect 30656 16720 30708 16726
rect 30656 16662 30708 16668
rect 30196 15360 30248 15366
rect 30196 15302 30248 15308
rect 28080 15156 28132 15162
rect 28080 15098 28132 15104
rect 28356 15156 28408 15162
rect 28356 15098 28408 15104
rect 28724 15156 28776 15162
rect 28724 15098 28776 15104
rect 29368 15156 29420 15162
rect 29368 15098 29420 15104
rect 27988 15020 28040 15026
rect 27988 14962 28040 14968
rect 28540 15020 28592 15026
rect 28540 14962 28592 14968
rect 27804 13932 27856 13938
rect 27804 13874 27856 13880
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 27816 13326 27844 13874
rect 28000 13870 28028 14962
rect 27988 13864 28040 13870
rect 27988 13806 28040 13812
rect 28552 13530 28580 14962
rect 29092 13728 29144 13734
rect 29092 13670 29144 13676
rect 28540 13524 28592 13530
rect 28540 13466 28592 13472
rect 29104 13394 29132 13670
rect 29380 13394 29408 15098
rect 30208 15094 30236 15302
rect 30196 15088 30248 15094
rect 30196 15030 30248 15036
rect 30668 14618 30696 16662
rect 31772 16590 31800 17138
rect 31760 16584 31812 16590
rect 31760 16526 31812 16532
rect 31392 16516 31444 16522
rect 31392 16458 31444 16464
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30944 14618 30972 15030
rect 30656 14612 30708 14618
rect 30656 14554 30708 14560
rect 30932 14612 30984 14618
rect 30932 14554 30984 14560
rect 29828 13864 29880 13870
rect 29828 13806 29880 13812
rect 29092 13388 29144 13394
rect 29092 13330 29144 13336
rect 29368 13388 29420 13394
rect 29368 13330 29420 13336
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 28264 13320 28316 13326
rect 28264 13262 28316 13268
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 29000 13320 29052 13326
rect 29000 13262 29052 13268
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27068 12980 27120 12986
rect 27068 12922 27120 12928
rect 26884 12912 26936 12918
rect 26884 12854 26936 12860
rect 26792 12776 26844 12782
rect 26792 12718 26844 12724
rect 26700 12640 26752 12646
rect 26700 12582 26752 12588
rect 26712 12102 26740 12582
rect 26804 12238 26832 12718
rect 26896 12238 26924 12854
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 27080 12102 27108 12922
rect 27264 12850 27292 13126
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27264 12646 27292 12786
rect 27252 12640 27304 12646
rect 27252 12582 27304 12588
rect 27448 12442 27476 13262
rect 27988 13252 28040 13258
rect 27988 13194 28040 13200
rect 27712 12912 27764 12918
rect 27540 12872 27712 12900
rect 27436 12436 27488 12442
rect 27436 12378 27488 12384
rect 27540 12238 27568 12872
rect 27712 12854 27764 12860
rect 27620 12708 27672 12714
rect 27620 12650 27672 12656
rect 27160 12232 27212 12238
rect 27158 12200 27160 12209
rect 27528 12232 27580 12238
rect 27212 12200 27214 12209
rect 27528 12174 27580 12180
rect 27158 12135 27214 12144
rect 26700 12096 26752 12102
rect 26700 12038 26752 12044
rect 27068 12096 27120 12102
rect 27068 12038 27120 12044
rect 27080 11898 27108 12038
rect 27068 11892 27120 11898
rect 27068 11834 27120 11840
rect 26700 11824 26752 11830
rect 26700 11766 26752 11772
rect 26712 11558 26740 11766
rect 27080 11762 27108 11834
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26712 11150 26740 11494
rect 26700 11144 26752 11150
rect 26700 11086 26752 11092
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 26608 9716 26660 9722
rect 26608 9658 26660 9664
rect 26252 8974 26280 9658
rect 27172 9654 27200 12135
rect 27632 11898 27660 12650
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27724 11898 27752 12038
rect 28000 11898 28028 13194
rect 28080 13184 28132 13190
rect 28080 13126 28132 13132
rect 28092 12782 28120 13126
rect 28276 12986 28304 13262
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28368 12782 28396 13262
rect 29012 12986 29040 13262
rect 29380 12986 29408 13330
rect 29000 12980 29052 12986
rect 29000 12922 29052 12928
rect 29368 12980 29420 12986
rect 29368 12922 29420 12928
rect 29736 12980 29788 12986
rect 29736 12922 29788 12928
rect 28080 12776 28132 12782
rect 28080 12718 28132 12724
rect 28356 12776 28408 12782
rect 28356 12718 28408 12724
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27712 11892 27764 11898
rect 27712 11834 27764 11840
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 27252 11552 27304 11558
rect 27252 11494 27304 11500
rect 27264 11150 27292 11494
rect 27724 11354 27752 11834
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27896 11688 27948 11694
rect 27802 11656 27858 11665
rect 27896 11630 27948 11636
rect 27802 11591 27804 11600
rect 27856 11591 27858 11600
rect 27804 11562 27856 11568
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27908 11286 27936 11630
rect 28092 11286 28120 11698
rect 28368 11354 28396 12718
rect 29748 12170 29776 12922
rect 29840 12306 29868 13806
rect 30668 12986 30696 14554
rect 30748 13252 30800 13258
rect 30748 13194 30800 13200
rect 30760 12986 30788 13194
rect 31404 13190 31432 16458
rect 31956 16454 31984 17138
rect 32232 16794 32260 18702
rect 32784 18086 32812 20182
rect 33152 19854 33180 21286
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 33324 20936 33376 20942
rect 33324 20878 33376 20884
rect 33336 20602 33364 20878
rect 34336 20868 34388 20874
rect 34336 20810 34388 20816
rect 33324 20596 33376 20602
rect 33324 20538 33376 20544
rect 33232 20528 33284 20534
rect 34348 20505 34376 20810
rect 33232 20470 33284 20476
rect 34334 20496 34390 20505
rect 33244 20058 33272 20470
rect 34334 20431 34390 20440
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 33140 19848 33192 19854
rect 33140 19790 33192 19796
rect 33600 19712 33652 19718
rect 33600 19654 33652 19660
rect 32772 18080 32824 18086
rect 32772 18022 32824 18028
rect 32220 16788 32272 16794
rect 32220 16730 32272 16736
rect 32680 16788 32732 16794
rect 32680 16730 32732 16736
rect 32692 16658 32720 16730
rect 32680 16652 32732 16658
rect 32680 16594 32732 16600
rect 31944 16448 31996 16454
rect 31944 16390 31996 16396
rect 31760 14816 31812 14822
rect 31760 14758 31812 14764
rect 31576 13932 31628 13938
rect 31576 13874 31628 13880
rect 31484 13864 31536 13870
rect 31484 13806 31536 13812
rect 31496 13530 31524 13806
rect 31588 13546 31616 13874
rect 31772 13734 31800 14758
rect 31956 14074 31984 16390
rect 32784 15910 32812 18022
rect 33612 17542 33640 19654
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34532 18426 34560 18702
rect 34612 18692 34664 18698
rect 34612 18634 34664 18640
rect 34520 18420 34572 18426
rect 34520 18362 34572 18368
rect 33784 18352 33836 18358
rect 34624 18329 34652 18634
rect 33784 18294 33836 18300
rect 34610 18320 34666 18329
rect 33796 17882 33824 18294
rect 34610 18255 34666 18264
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 33784 17876 33836 17882
rect 33784 17818 33836 17824
rect 33600 17536 33652 17542
rect 33600 17478 33652 17484
rect 33140 16720 33192 16726
rect 33140 16662 33192 16668
rect 33152 16182 33180 16662
rect 33140 16176 33192 16182
rect 33140 16118 33192 16124
rect 32772 15904 32824 15910
rect 32772 15846 32824 15852
rect 32784 14958 32812 15846
rect 33612 15502 33640 17478
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34520 16584 34572 16590
rect 34520 16526 34572 16532
rect 34532 16250 34560 16526
rect 34612 16516 34664 16522
rect 34612 16458 34664 16464
rect 34520 16244 34572 16250
rect 34520 16186 34572 16192
rect 33968 16176 34020 16182
rect 34624 16153 34652 16458
rect 33968 16118 34020 16124
rect 34610 16144 34666 16153
rect 33980 15706 34008 16118
rect 34610 16079 34666 16088
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 33968 15700 34020 15706
rect 33968 15642 34020 15648
rect 33600 15496 33652 15502
rect 33600 15438 33652 15444
rect 32772 14952 32824 14958
rect 32772 14894 32824 14900
rect 31944 14068 31996 14074
rect 31944 14010 31996 14016
rect 32784 13870 32812 14894
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 34152 14000 34204 14006
rect 34624 13977 34652 14282
rect 34152 13942 34204 13948
rect 34610 13968 34666 13977
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 32772 13864 32824 13870
rect 32772 13806 32824 13812
rect 31760 13728 31812 13734
rect 31760 13670 31812 13676
rect 31484 13524 31536 13530
rect 31588 13518 31800 13546
rect 32232 13530 32260 13806
rect 31484 13466 31536 13472
rect 31772 13462 31800 13518
rect 32220 13524 32272 13530
rect 32220 13466 32272 13472
rect 31760 13456 31812 13462
rect 31760 13398 31812 13404
rect 31668 13320 31720 13326
rect 31668 13262 31720 13268
rect 31392 13184 31444 13190
rect 31392 13126 31444 13132
rect 31404 12986 31432 13126
rect 30656 12980 30708 12986
rect 30656 12922 30708 12928
rect 30748 12980 30800 12986
rect 30748 12922 30800 12928
rect 31392 12980 31444 12986
rect 31392 12922 31444 12928
rect 30668 12434 30696 12922
rect 31680 12918 31708 13262
rect 31668 12912 31720 12918
rect 31668 12854 31720 12860
rect 31772 12850 31800 13398
rect 31944 13184 31996 13190
rect 31944 13126 31996 13132
rect 31956 12850 31984 13126
rect 31760 12844 31812 12850
rect 31760 12786 31812 12792
rect 31944 12844 31996 12850
rect 31944 12786 31996 12792
rect 30392 12406 30696 12434
rect 29828 12300 29880 12306
rect 29828 12242 29880 12248
rect 29736 12164 29788 12170
rect 29736 12106 29788 12112
rect 29748 11898 29776 12106
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 29012 11354 29040 11834
rect 30392 11762 30420 12406
rect 30932 12232 30984 12238
rect 30932 12174 30984 12180
rect 30944 11898 30972 12174
rect 31300 12096 31352 12102
rect 31300 12038 31352 12044
rect 30932 11892 30984 11898
rect 30932 11834 30984 11840
rect 31312 11830 31340 12038
rect 31300 11824 31352 11830
rect 31300 11766 31352 11772
rect 31576 11824 31628 11830
rect 31576 11766 31628 11772
rect 30380 11756 30432 11762
rect 30380 11698 30432 11704
rect 28356 11348 28408 11354
rect 28356 11290 28408 11296
rect 29000 11348 29052 11354
rect 29000 11290 29052 11296
rect 27896 11280 27948 11286
rect 27896 11222 27948 11228
rect 28080 11280 28132 11286
rect 28080 11222 28132 11228
rect 27252 11144 27304 11150
rect 27620 11144 27672 11150
rect 27252 11086 27304 11092
rect 27540 11104 27620 11132
rect 27540 10810 27568 11104
rect 27620 11086 27672 11092
rect 28908 11008 28960 11014
rect 28908 10950 28960 10956
rect 27528 10804 27580 10810
rect 27528 10746 27580 10752
rect 28920 10674 28948 10950
rect 29012 10810 29040 11290
rect 30392 11082 30420 11698
rect 31484 11688 31536 11694
rect 31484 11630 31536 11636
rect 30472 11552 30524 11558
rect 30472 11494 30524 11500
rect 30484 11354 30512 11494
rect 31496 11354 31524 11630
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 31484 11348 31536 11354
rect 31484 11290 31536 11296
rect 30380 11076 30432 11082
rect 30380 11018 30432 11024
rect 31116 11076 31168 11082
rect 31116 11018 31168 11024
rect 29000 10804 29052 10810
rect 29000 10746 29052 10752
rect 29368 10804 29420 10810
rect 29368 10746 29420 10752
rect 28908 10668 28960 10674
rect 28908 10610 28960 10616
rect 27252 10600 27304 10606
rect 27252 10542 27304 10548
rect 27264 10062 27292 10542
rect 27528 10464 27580 10470
rect 27528 10406 27580 10412
rect 27252 10056 27304 10062
rect 27252 9998 27304 10004
rect 27160 9648 27212 9654
rect 27160 9590 27212 9596
rect 27540 9586 27568 10406
rect 28920 10266 28948 10610
rect 28908 10260 28960 10266
rect 28908 10202 28960 10208
rect 28080 10124 28132 10130
rect 28080 10066 28132 10072
rect 28092 9722 28120 10066
rect 29380 10062 29408 10746
rect 30104 10464 30156 10470
rect 30104 10406 30156 10412
rect 29368 10056 29420 10062
rect 29368 9998 29420 10004
rect 28540 9920 28592 9926
rect 28540 9862 28592 9868
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 28080 9716 28132 9722
rect 28080 9658 28132 9664
rect 28552 9654 28580 9862
rect 29288 9654 29316 9862
rect 28540 9648 28592 9654
rect 28540 9590 28592 9596
rect 29276 9648 29328 9654
rect 29276 9590 29328 9596
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 29380 9518 29408 9998
rect 30116 9994 30144 10406
rect 31128 10062 31156 11018
rect 31496 10674 31524 11290
rect 31588 11150 31616 11766
rect 31772 11354 31800 12786
rect 31956 11898 31984 12786
rect 32680 12708 32732 12714
rect 32680 12650 32732 12656
rect 32692 12442 32720 12650
rect 32680 12436 32732 12442
rect 32680 12378 32732 12384
rect 32784 12238 32812 13806
rect 34164 13530 34192 13942
rect 34610 13903 34666 13912
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34152 13524 34204 13530
rect 34152 13466 34204 13472
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 34716 12646 34744 13126
rect 34704 12640 34756 12646
rect 34704 12582 34756 12588
rect 34716 12238 34744 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 32772 12232 32824 12238
rect 32772 12174 32824 12180
rect 34704 12232 34756 12238
rect 34704 12174 34756 12180
rect 31944 11892 31996 11898
rect 31944 11834 31996 11840
rect 31852 11552 31904 11558
rect 31852 11494 31904 11500
rect 31864 11354 31892 11494
rect 31760 11348 31812 11354
rect 31760 11290 31812 11296
rect 31852 11348 31904 11354
rect 31852 11290 31904 11296
rect 31576 11144 31628 11150
rect 31576 11086 31628 11092
rect 31760 11144 31812 11150
rect 31760 11086 31812 11092
rect 31588 10674 31616 11086
rect 31772 10674 31800 11086
rect 31956 10810 31984 11834
rect 32784 11150 32812 12174
rect 34520 12096 34572 12102
rect 34520 12038 34572 12044
rect 34532 11898 34560 12038
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 34612 11212 34664 11218
rect 34612 11154 34664 11160
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 32784 10810 32812 11086
rect 31944 10804 31996 10810
rect 31944 10746 31996 10752
rect 32772 10804 32824 10810
rect 32772 10746 32824 10752
rect 31484 10668 31536 10674
rect 31484 10610 31536 10616
rect 31576 10668 31628 10674
rect 31576 10610 31628 10616
rect 31760 10668 31812 10674
rect 31760 10610 31812 10616
rect 31300 10532 31352 10538
rect 31300 10474 31352 10480
rect 31312 10266 31340 10474
rect 31392 10464 31444 10470
rect 31392 10406 31444 10412
rect 31404 10266 31432 10406
rect 31956 10266 31984 10746
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 31300 10260 31352 10266
rect 31300 10202 31352 10208
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31944 10260 31996 10266
rect 31944 10202 31996 10208
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 30104 9988 30156 9994
rect 30104 9930 30156 9936
rect 31128 9518 31156 9998
rect 31312 9586 31340 10202
rect 32232 10062 32260 10610
rect 32784 10062 32812 10746
rect 34060 10464 34112 10470
rect 34060 10406 34112 10412
rect 34072 10062 34100 10406
rect 32220 10056 32272 10062
rect 32772 10056 32824 10062
rect 32220 9998 32272 10004
rect 32692 10004 32772 10010
rect 32692 9998 32824 10004
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 32692 9982 32812 9998
rect 32220 9920 32272 9926
rect 32220 9862 32272 9868
rect 31300 9580 31352 9586
rect 31300 9522 31352 9528
rect 32232 9518 32260 9862
rect 29368 9512 29420 9518
rect 29368 9454 29420 9460
rect 31116 9512 31168 9518
rect 31116 9454 31168 9460
rect 32220 9512 32272 9518
rect 32220 9454 32272 9460
rect 32588 9376 32640 9382
rect 32588 9318 32640 9324
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 25964 8900 26016 8906
rect 25964 8842 26016 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 26252 8566 26280 8910
rect 32600 8634 32628 9318
rect 32588 8628 32640 8634
rect 32588 8570 32640 8576
rect 32692 8566 32720 9982
rect 32772 9920 32824 9926
rect 32772 9862 32824 9868
rect 32784 9586 32812 9862
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32956 9376 33008 9382
rect 32956 9318 33008 9324
rect 32968 9178 32996 9318
rect 32956 9172 33008 9178
rect 32956 9114 33008 9120
rect 34072 8974 34100 9998
rect 34520 9920 34572 9926
rect 34520 9862 34572 9868
rect 34532 9586 34560 9862
rect 34520 9580 34572 9586
rect 34520 9522 34572 9528
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 33048 8832 33100 8838
rect 33048 8774 33100 8780
rect 33508 8832 33560 8838
rect 33508 8774 33560 8780
rect 26240 8560 26292 8566
rect 26240 8502 26292 8508
rect 32680 8560 32732 8566
rect 32680 8502 32732 8508
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 27816 2650 27844 8434
rect 32692 8090 32720 8502
rect 32680 8084 32732 8090
rect 32680 8026 32732 8032
rect 33060 7954 33088 8774
rect 33520 8566 33548 8774
rect 34072 8634 34100 8910
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 33508 8560 33560 8566
rect 33508 8502 33560 8508
rect 34244 8356 34296 8362
rect 34244 8298 34296 8304
rect 33048 7948 33100 7954
rect 33048 7890 33100 7896
rect 34256 6914 34284 8298
rect 34428 8288 34480 8294
rect 34428 8230 34480 8236
rect 34440 7886 34468 8230
rect 34428 7880 34480 7886
rect 34428 7822 34480 7828
rect 34520 7744 34572 7750
rect 34520 7686 34572 7692
rect 34256 6886 34376 6914
rect 34348 5710 34376 6886
rect 34336 5704 34388 5710
rect 34336 5646 34388 5652
rect 34060 5636 34112 5642
rect 34060 5578 34112 5584
rect 34072 5273 34100 5578
rect 34058 5264 34114 5273
rect 34058 5199 34114 5208
rect 34532 3534 34560 7686
rect 34624 7410 34652 11154
rect 34716 11150 34744 12174
rect 34794 11792 34850 11801
rect 34794 11727 34796 11736
rect 34848 11727 34850 11736
rect 34796 11698 34848 11704
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34704 11144 34756 11150
rect 34704 11086 34756 11092
rect 34716 10470 34744 11086
rect 34704 10464 34756 10470
rect 34704 10406 34756 10412
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34794 9616 34850 9625
rect 34794 9551 34796 9560
rect 34848 9551 34850 9560
rect 34796 9522 34848 9528
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34794 7440 34850 7449
rect 34612 7404 34664 7410
rect 34794 7375 34796 7384
rect 34612 7346 34664 7352
rect 34848 7375 34850 7384
rect 34796 7346 34848 7352
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34520 3528 34572 3534
rect 34520 3470 34572 3476
rect 34612 3460 34664 3466
rect 34612 3402 34664 3408
rect 34624 3097 34652 3402
rect 34610 3088 34666 3097
rect 34610 3023 34666 3032
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 952 2009 980 2382
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 9140 1306 9168 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 27356 1306 27384 2382
rect 9048 1278 9168 1306
rect 27264 1278 27384 1306
rect 9048 800 9076 1278
rect 27264 800 27292 1278
rect 9034 0 9090 800
rect 27250 0 27306 800
<< via2 >>
rect 938 36760 994 36816
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 938 34584 994 34640
rect 938 32408 994 32464
rect 1398 30232 1454 30288
rect 938 28056 994 28112
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 938 25900 994 25936
rect 938 25880 940 25900
rect 940 25880 992 25900
rect 992 25880 994 25900
rect 938 23704 994 23760
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 938 21528 994 21584
rect 938 19352 994 19408
rect 938 17176 994 17232
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 1398 15136 1454 15192
rect 938 12844 994 12880
rect 938 12824 940 12844
rect 940 12824 992 12844
rect 992 12824 994 12844
rect 1398 10920 1454 10976
rect 938 8472 994 8528
rect 938 6296 994 6352
rect 938 4120 994 4176
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 14186 24148 14188 24168
rect 14188 24148 14240 24168
rect 14240 24148 14242 24168
rect 11978 21684 12034 21720
rect 11978 21664 11980 21684
rect 11980 21664 12032 21684
rect 12032 21664 12034 21684
rect 12622 23976 12678 24032
rect 14186 24112 14242 24148
rect 12346 19624 12402 19680
rect 15198 24112 15254 24168
rect 13174 18028 13176 18048
rect 13176 18028 13228 18048
rect 13228 18028 13230 18048
rect 13174 17992 13230 18028
rect 15014 19624 15070 19680
rect 14186 16108 14242 16144
rect 14186 16088 14188 16108
rect 14188 16088 14240 16108
rect 14240 16088 14242 16108
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 17406 23976 17462 24032
rect 16302 21664 16358 21720
rect 16578 19660 16580 19680
rect 16580 19660 16632 19680
rect 16632 19660 16634 19680
rect 16578 19624 16634 19660
rect 16578 19508 16634 19544
rect 16578 19488 16580 19508
rect 16580 19488 16632 19508
rect 16632 19488 16634 19508
rect 15014 12280 15070 12336
rect 15658 12300 15714 12336
rect 15658 12280 15660 12300
rect 15660 12280 15712 12300
rect 15712 12280 15714 12300
rect 15934 12180 15936 12200
rect 15936 12180 15988 12200
rect 15988 12180 15990 12200
rect 15934 12144 15990 12180
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20626 23704 20682 23760
rect 17958 19508 18014 19544
rect 17958 19488 17960 19508
rect 17960 19488 18012 19508
rect 18012 19488 18014 19508
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19338 17992 19394 18048
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 18878 16124 18880 16144
rect 18880 16124 18932 16144
rect 18932 16124 18934 16144
rect 18878 16088 18934 16124
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 17222 12180 17224 12200
rect 17224 12180 17276 12200
rect 17276 12180 17278 12200
rect 17222 12144 17278 12180
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 22650 23740 22652 23760
rect 22652 23740 22704 23760
rect 22704 23740 22706 23760
rect 22650 23704 22706 23740
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19982 10684 19984 10704
rect 19984 10684 20036 10704
rect 20036 10684 20038 10704
rect 19982 10648 20038 10684
rect 21362 11620 21418 11656
rect 21362 11600 21364 11620
rect 21364 11600 21416 11620
rect 21416 11600 21418 11620
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 22834 12144 22890 12200
rect 25778 10648 25834 10704
rect 34334 35672 34390 35728
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34058 31320 34114 31376
rect 34610 33496 34666 33552
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34610 29144 34666 29200
rect 34702 26988 34758 27024
rect 34702 26968 34704 26988
rect 34704 26968 34756 26988
rect 34756 26968 34758 26988
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34058 24792 34114 24848
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34610 22616 34666 22672
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 27158 12180 27160 12200
rect 27160 12180 27212 12200
rect 27212 12180 27214 12200
rect 27158 12144 27214 12180
rect 27802 11620 27858 11656
rect 27802 11600 27804 11620
rect 27804 11600 27856 11620
rect 27856 11600 27858 11620
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34334 20440 34390 20496
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34610 18264 34666 18320
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34610 16088 34666 16144
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34610 13912 34666 13968
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34058 5208 34114 5264
rect 34794 11756 34850 11792
rect 34794 11736 34796 11756
rect 34796 11736 34848 11756
rect 34848 11736 34850 11756
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34794 9580 34850 9616
rect 34794 9560 34796 9580
rect 34796 9560 34848 9580
rect 34848 9560 34850 9580
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34794 7404 34850 7440
rect 34794 7384 34796 7404
rect 34796 7384 34848 7404
rect 34848 7384 34850 7404
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34610 3032 34666 3088
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 938 1944 994 2000
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 34329 35730 34395 35733
rect 35600 35730 36400 35760
rect 34329 35728 36400 35730
rect 34329 35672 34334 35728
rect 34390 35672 36400 35728
rect 34329 35670 36400 35672
rect 34329 35667 34395 35670
rect 35600 35640 36400 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 0 34642 800 34672
rect 933 34642 999 34645
rect 0 34640 999 34642
rect 0 34584 938 34640
rect 994 34584 999 34640
rect 0 34582 999 34584
rect 0 34552 800 34582
rect 933 34579 999 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 34605 33554 34671 33557
rect 35600 33554 36400 33584
rect 34605 33552 36400 33554
rect 34605 33496 34610 33552
rect 34666 33496 36400 33552
rect 34605 33494 36400 33496
rect 34605 33491 34671 33494
rect 35600 33464 36400 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 0 32466 800 32496
rect 933 32466 999 32469
rect 0 32464 999 32466
rect 0 32408 938 32464
rect 994 32408 999 32464
rect 0 32406 999 32408
rect 0 32376 800 32406
rect 933 32403 999 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 34053 31378 34119 31381
rect 35600 31378 36400 31408
rect 34053 31376 36400 31378
rect 34053 31320 34058 31376
rect 34114 31320 36400 31376
rect 34053 31318 36400 31320
rect 34053 31315 34119 31318
rect 35600 31288 36400 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 30290 800 30320
rect 1393 30290 1459 30293
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 800 30230
rect 1393 30227 1459 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 34605 29202 34671 29205
rect 35600 29202 36400 29232
rect 34605 29200 36400 29202
rect 34605 29144 34610 29200
rect 34666 29144 36400 29200
rect 34605 29142 36400 29144
rect 34605 29139 34671 29142
rect 35600 29112 36400 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 0 28114 800 28144
rect 933 28114 999 28117
rect 0 28112 999 28114
rect 0 28056 938 28112
rect 994 28056 999 28112
rect 0 28054 999 28056
rect 0 28024 800 28054
rect 933 28051 999 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 34697 27026 34763 27029
rect 35600 27026 36400 27056
rect 34697 27024 36400 27026
rect 34697 26968 34702 27024
rect 34758 26968 36400 27024
rect 34697 26966 36400 26968
rect 34697 26963 34763 26966
rect 35600 26936 36400 26966
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25938 800 25968
rect 933 25938 999 25941
rect 0 25936 999 25938
rect 0 25880 938 25936
rect 994 25880 999 25936
rect 0 25878 999 25880
rect 0 25848 800 25878
rect 933 25875 999 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 34053 24850 34119 24853
rect 35600 24850 36400 24880
rect 34053 24848 36400 24850
rect 34053 24792 34058 24848
rect 34114 24792 36400 24848
rect 34053 24790 36400 24792
rect 34053 24787 34119 24790
rect 35600 24760 36400 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 14181 24170 14247 24173
rect 15193 24170 15259 24173
rect 14181 24168 15259 24170
rect 14181 24112 14186 24168
rect 14242 24112 15198 24168
rect 15254 24112 15259 24168
rect 14181 24110 15259 24112
rect 14181 24107 14247 24110
rect 15193 24107 15259 24110
rect 12617 24034 12683 24037
rect 17401 24034 17467 24037
rect 12617 24032 17467 24034
rect 12617 23976 12622 24032
rect 12678 23976 17406 24032
rect 17462 23976 17467 24032
rect 12617 23974 17467 23976
rect 12617 23971 12683 23974
rect 17401 23971 17467 23974
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 20621 23762 20687 23765
rect 22645 23762 22711 23765
rect 20621 23760 22711 23762
rect 20621 23704 20626 23760
rect 20682 23704 22650 23760
rect 22706 23704 22711 23760
rect 20621 23702 22711 23704
rect 20621 23699 20687 23702
rect 22645 23699 22711 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 34605 22674 34671 22677
rect 35600 22674 36400 22704
rect 34605 22672 36400 22674
rect 34605 22616 34610 22672
rect 34666 22616 36400 22672
rect 34605 22614 36400 22616
rect 34605 22611 34671 22614
rect 35600 22584 36400 22614
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 11973 21722 12039 21725
rect 16297 21722 16363 21725
rect 11973 21720 16363 21722
rect 11973 21664 11978 21720
rect 12034 21664 16302 21720
rect 16358 21664 16363 21720
rect 11973 21662 16363 21664
rect 11973 21659 12039 21662
rect 16297 21659 16363 21662
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 34329 20498 34395 20501
rect 35600 20498 36400 20528
rect 34329 20496 36400 20498
rect 34329 20440 34334 20496
rect 34390 20440 36400 20496
rect 34329 20438 36400 20440
rect 34329 20435 34395 20438
rect 35600 20408 36400 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 12341 19682 12407 19685
rect 15009 19682 15075 19685
rect 16573 19682 16639 19685
rect 12341 19680 16639 19682
rect 12341 19624 12346 19680
rect 12402 19624 15014 19680
rect 15070 19624 16578 19680
rect 16634 19624 16639 19680
rect 12341 19622 16639 19624
rect 12341 19619 12407 19622
rect 15009 19619 15075 19622
rect 16573 19619 16639 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 16573 19546 16639 19549
rect 17953 19546 18019 19549
rect 16573 19544 18019 19546
rect 16573 19488 16578 19544
rect 16634 19488 17958 19544
rect 18014 19488 18019 19544
rect 16573 19486 18019 19488
rect 16573 19483 16639 19486
rect 17953 19483 18019 19486
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 34605 18322 34671 18325
rect 35600 18322 36400 18352
rect 34605 18320 36400 18322
rect 34605 18264 34610 18320
rect 34666 18264 36400 18320
rect 34605 18262 36400 18264
rect 34605 18259 34671 18262
rect 35600 18232 36400 18262
rect 13169 18050 13235 18053
rect 19333 18050 19399 18053
rect 13169 18048 19399 18050
rect 13169 17992 13174 18048
rect 13230 17992 19338 18048
rect 19394 17992 19399 18048
rect 13169 17990 19399 17992
rect 13169 17987 13235 17990
rect 19333 17987 19399 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 0 17234 800 17264
rect 933 17234 999 17237
rect 0 17232 999 17234
rect 0 17176 938 17232
rect 994 17176 999 17232
rect 0 17174 999 17176
rect 0 17144 800 17174
rect 933 17171 999 17174
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 14181 16146 14247 16149
rect 18873 16146 18939 16149
rect 14181 16144 18939 16146
rect 14181 16088 14186 16144
rect 14242 16088 18878 16144
rect 18934 16088 18939 16144
rect 14181 16086 18939 16088
rect 14181 16083 14247 16086
rect 18873 16083 18939 16086
rect 34605 16146 34671 16149
rect 35600 16146 36400 16176
rect 34605 16144 36400 16146
rect 34605 16088 34610 16144
rect 34666 16088 36400 16144
rect 34605 16086 36400 16088
rect 34605 16083 34671 16086
rect 35600 16056 36400 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 1393 15194 1459 15197
rect 798 15192 1459 15194
rect 798 15136 1398 15192
rect 1454 15136 1459 15192
rect 798 15134 1459 15136
rect 798 15088 858 15134
rect 1393 15131 1459 15134
rect 0 14998 858 15088
rect 0 14968 800 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 34605 13970 34671 13973
rect 35600 13970 36400 14000
rect 34605 13968 36400 13970
rect 34605 13912 34610 13968
rect 34666 13912 36400 13968
rect 34605 13910 36400 13912
rect 34605 13907 34671 13910
rect 35600 13880 36400 13910
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 15009 12338 15075 12341
rect 15653 12338 15719 12341
rect 15009 12336 15719 12338
rect 15009 12280 15014 12336
rect 15070 12280 15658 12336
rect 15714 12280 15719 12336
rect 15009 12278 15719 12280
rect 15009 12275 15075 12278
rect 15653 12275 15719 12278
rect 15929 12202 15995 12205
rect 17217 12202 17283 12205
rect 15929 12200 17283 12202
rect 15929 12144 15934 12200
rect 15990 12144 17222 12200
rect 17278 12144 17283 12200
rect 15929 12142 17283 12144
rect 15929 12139 15995 12142
rect 17217 12139 17283 12142
rect 22829 12202 22895 12205
rect 27153 12202 27219 12205
rect 22829 12200 27219 12202
rect 22829 12144 22834 12200
rect 22890 12144 27158 12200
rect 27214 12144 27219 12200
rect 22829 12142 27219 12144
rect 22829 12139 22895 12142
rect 27153 12139 27219 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 34789 11794 34855 11797
rect 35600 11794 36400 11824
rect 34789 11792 36400 11794
rect 34789 11736 34794 11792
rect 34850 11736 36400 11792
rect 34789 11734 36400 11736
rect 34789 11731 34855 11734
rect 35600 11704 36400 11734
rect 21357 11658 21423 11661
rect 27797 11658 27863 11661
rect 21357 11656 27863 11658
rect 21357 11600 21362 11656
rect 21418 11600 27802 11656
rect 27858 11600 27863 11656
rect 21357 11598 27863 11600
rect 21357 11595 21423 11598
rect 27797 11595 27863 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 1393 10978 1459 10981
rect 798 10976 1459 10978
rect 798 10920 1398 10976
rect 1454 10920 1459 10976
rect 798 10918 1459 10920
rect 798 10736 858 10918
rect 1393 10915 1459 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 0 10646 858 10736
rect 19977 10706 20043 10709
rect 25773 10706 25839 10709
rect 19977 10704 25839 10706
rect 19977 10648 19982 10704
rect 20038 10648 25778 10704
rect 25834 10648 25839 10704
rect 19977 10646 25839 10648
rect 0 10616 800 10646
rect 19977 10643 20043 10646
rect 25773 10643 25839 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 34789 9618 34855 9621
rect 35600 9618 36400 9648
rect 34789 9616 36400 9618
rect 34789 9560 34794 9616
rect 34850 9560 36400 9616
rect 34789 9558 36400 9560
rect 34789 9555 34855 9558
rect 35600 9528 36400 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 34789 7442 34855 7445
rect 35600 7442 36400 7472
rect 34789 7440 36400 7442
rect 34789 7384 34794 7440
rect 34850 7384 36400 7440
rect 34789 7382 36400 7384
rect 34789 7379 34855 7382
rect 35600 7352 36400 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 34053 5266 34119 5269
rect 35600 5266 36400 5296
rect 34053 5264 36400 5266
rect 34053 5208 34058 5264
rect 34114 5208 36400 5264
rect 34053 5206 36400 5208
rect 34053 5203 34119 5206
rect 35600 5176 36400 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 34605 3090 34671 3093
rect 35600 3090 36400 3120
rect 34605 3088 36400 3090
rect 34605 3032 34610 3088
rect 34666 3032 36400 3088
rect 34605 3030 36400 3032
rect 34605 3027 34671 3030
rect 35600 3000 36400 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
<< via3 >>
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 36480 4528 36496
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 35936 19888 36496
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 36480 35248 36496
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__or4_1  _0543_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0544_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0545_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5704 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0546_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0547_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 7084 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0548_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0549_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0550_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4600 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0551_
timestamp 1688980957
transform 1 0 4600 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0552_
timestamp 1688980957
transform 1 0 3956 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0553_
timestamp 1688980957
transform 1 0 3956 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0554_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0555_
timestamp 1688980957
transform 1 0 3680 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0556_
timestamp 1688980957
transform -1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0557_
timestamp 1688980957
transform 1 0 4784 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0558_
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0559_
timestamp 1688980957
transform 1 0 4600 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0560_
timestamp 1688980957
transform -1 0 5796 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0561_
timestamp 1688980957
transform -1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _0562_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4048 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0563_
timestamp 1688980957
transform 1 0 4600 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0564_
timestamp 1688980957
transform -1 0 5428 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0565_
timestamp 1688980957
transform 1 0 5796 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0566_
timestamp 1688980957
transform -1 0 6624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0567_
timestamp 1688980957
transform 1 0 4692 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0568_
timestamp 1688980957
transform 1 0 5152 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0569_
timestamp 1688980957
transform -1 0 5152 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0570_
timestamp 1688980957
transform 1 0 5152 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0571_
timestamp 1688980957
transform -1 0 5888 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0572_
timestamp 1688980957
transform 1 0 4784 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0573_
timestamp 1688980957
transform 1 0 4232 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0574_
timestamp 1688980957
transform 1 0 3772 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _0575_
timestamp 1688980957
transform -1 0 5704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0576_
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0577_
timestamp 1688980957
transform -1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0578_
timestamp 1688980957
transform 1 0 5612 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0579_
timestamp 1688980957
transform -1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0580_
timestamp 1688980957
transform -1 0 7268 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0581_
timestamp 1688980957
transform 1 0 31280 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0582_
timestamp 1688980957
transform 1 0 31556 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0583_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31924 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0584_
timestamp 1688980957
transform 1 0 31648 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0585_
timestamp 1688980957
transform -1 0 32108 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0586_
timestamp 1688980957
transform -1 0 30912 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0587_
timestamp 1688980957
transform 1 0 30452 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0588_
timestamp 1688980957
transform 1 0 5152 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0589_
timestamp 1688980957
transform 1 0 6072 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0590_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29716 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0591_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0592_
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0593_
timestamp 1688980957
transform -1 0 31188 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0594_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29900 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0595_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30820 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0596_
timestamp 1688980957
transform 1 0 30912 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0597_
timestamp 1688980957
transform 1 0 31464 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0598_
timestamp 1688980957
transform 1 0 30820 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0599_
timestamp 1688980957
transform 1 0 30912 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0600_
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0601_
timestamp 1688980957
transform -1 0 31648 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0602_
timestamp 1688980957
transform 1 0 30728 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0603_
timestamp 1688980957
transform -1 0 31372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0604_
timestamp 1688980957
transform 1 0 31004 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0605_
timestamp 1688980957
transform -1 0 31464 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0606_
timestamp 1688980957
transform 1 0 31004 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0607_
timestamp 1688980957
transform 1 0 32016 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0608_
timestamp 1688980957
transform 1 0 31372 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0609_
timestamp 1688980957
transform 1 0 32384 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0610_
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0611_
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0612_
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0613_
timestamp 1688980957
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0614_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0615_
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0616_
timestamp 1688980957
transform 1 0 31372 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0617_
timestamp 1688980957
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0618_
timestamp 1688980957
transform 1 0 31832 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0619_
timestamp 1688980957
transform 1 0 32016 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0620_
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0621_
timestamp 1688980957
transform -1 0 33028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0622_
timestamp 1688980957
transform -1 0 33120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0623_
timestamp 1688980957
transform 1 0 9016 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _0624_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _0625_
timestamp 1688980957
transform 1 0 10212 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0626_
timestamp 1688980957
transform 1 0 18400 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _0627_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8372 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _0628_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  _0629_
timestamp 1688980957
transform 1 0 10580 0 1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _0630_
timestamp 1688980957
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_1  _0631_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17296 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0632_
timestamp 1688980957
transform 1 0 15824 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0633_
timestamp 1688980957
transform -1 0 17756 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0634_
timestamp 1688980957
transform 1 0 16468 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0635_
timestamp 1688980957
transform -1 0 11776 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0636_
timestamp 1688980957
transform 1 0 11040 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0637_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0638_
timestamp 1688980957
transform -1 0 12696 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0639_
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0640_
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0641_
timestamp 1688980957
transform -1 0 19136 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0642_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0643_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19044 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0644_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13340 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0645_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13892 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0646_
timestamp 1688980957
transform -1 0 15732 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0647_
timestamp 1688980957
transform -1 0 15364 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0648_
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0649_
timestamp 1688980957
transform -1 0 15824 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0650_
timestamp 1688980957
transform 1 0 14628 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0651_
timestamp 1688980957
transform 1 0 15272 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0652_
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0653_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0654_
timestamp 1688980957
transform -1 0 14904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0655_
timestamp 1688980957
transform 1 0 12696 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0656_
timestamp 1688980957
transform 1 0 13432 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0657_
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0658_
timestamp 1688980957
transform 1 0 16744 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0659_
timestamp 1688980957
transform -1 0 17664 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0660_
timestamp 1688980957
transform 1 0 18216 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_1  _0661_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18308 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _0662_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0663_
timestamp 1688980957
transform -1 0 16376 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0664_
timestamp 1688980957
transform 1 0 14996 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0665_
timestamp 1688980957
transform -1 0 15364 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0666_
timestamp 1688980957
transform 1 0 15364 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _0667_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0668_
timestamp 1688980957
transform 1 0 18400 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0669_
timestamp 1688980957
transform 1 0 18308 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0670_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17940 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0671_
timestamp 1688980957
transform -1 0 20148 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0672_
timestamp 1688980957
transform 1 0 16744 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0673_
timestamp 1688980957
transform 1 0 17848 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0674_
timestamp 1688980957
transform -1 0 20240 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0675_
timestamp 1688980957
transform 1 0 19412 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0676_
timestamp 1688980957
transform -1 0 20608 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _0677_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20240 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0678_
timestamp 1688980957
transform 1 0 18952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0679_
timestamp 1688980957
transform -1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0680_
timestamp 1688980957
transform -1 0 21620 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0681_
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _0682_
timestamp 1688980957
transform 1 0 10764 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0683_
timestamp 1688980957
transform -1 0 18308 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _0684_
timestamp 1688980957
transform 1 0 10120 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0685_
timestamp 1688980957
transform 1 0 19044 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _0686_
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0687_
timestamp 1688980957
transform 1 0 16008 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_4  _0688_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_4  _0689_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0690_
timestamp 1688980957
transform 1 0 11592 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0691_
timestamp 1688980957
transform 1 0 11960 0 1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0692_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0693_
timestamp 1688980957
transform 1 0 10948 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0694_
timestamp 1688980957
transform 1 0 11408 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _0695_
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0696_
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0697_
timestamp 1688980957
transform -1 0 12788 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0698_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0699_
timestamp 1688980957
transform -1 0 18584 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0700_
timestamp 1688980957
transform 1 0 18400 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_2  _0701_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _0702_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0703_
timestamp 1688980957
transform -1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0704_
timestamp 1688980957
transform 1 0 14076 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0705_
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0706_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _0707_
timestamp 1688980957
transform 1 0 15732 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0708_
timestamp 1688980957
transform 1 0 13524 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0709_
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0710_
timestamp 1688980957
transform 1 0 17848 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0711_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0712_
timestamp 1688980957
transform -1 0 19596 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0713_
timestamp 1688980957
transform -1 0 19872 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0714_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0715_
timestamp 1688980957
transform -1 0 15272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0716_
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nor3_1  _0717_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14996 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0718_
timestamp 1688980957
transform -1 0 15732 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _0719_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0720_
timestamp 1688980957
transform -1 0 15180 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0721_
timestamp 1688980957
transform 1 0 18400 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0722_
timestamp 1688980957
transform 1 0 19412 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0723_
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0724_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _0725_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17480 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0726_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14352 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0727_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14352 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1688980957
transform -1 0 16376 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0729_
timestamp 1688980957
transform -1 0 20608 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0730_
timestamp 1688980957
transform -1 0 19044 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0731_
timestamp 1688980957
transform -1 0 17020 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0732_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0733_
timestamp 1688980957
transform -1 0 15824 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0734_
timestamp 1688980957
transform -1 0 16560 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0735_
timestamp 1688980957
transform -1 0 16560 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0736_
timestamp 1688980957
transform -1 0 17204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0737_
timestamp 1688980957
transform 1 0 16560 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31oi_1  _0738_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _0739_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17388 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0740_
timestamp 1688980957
transform -1 0 19504 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0741_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_2  _0742_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1688980957
transform 1 0 21252 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0744_
timestamp 1688980957
transform 1 0 9016 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _0745_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13800 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0746_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _0747_
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_1  _0748_
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_2  _0749_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0750_
timestamp 1688980957
transform -1 0 9660 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0751_
timestamp 1688980957
transform 1 0 9844 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0752_
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _0753_
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _0754_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15180 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0755_
timestamp 1688980957
transform -1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0756_
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0757_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_1  _0758_
timestamp 1688980957
transform -1 0 15732 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0759_
timestamp 1688980957
transform -1 0 14628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0760_
timestamp 1688980957
transform 1 0 15548 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0761_
timestamp 1688980957
transform -1 0 14260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0762_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14720 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__clkinvlp_2  _0763_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0764_
timestamp 1688980957
transform -1 0 11316 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0765_
timestamp 1688980957
transform -1 0 13984 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0766_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  _0767_
timestamp 1688980957
transform -1 0 17480 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0768_
timestamp 1688980957
transform 1 0 17204 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0769_
timestamp 1688980957
transform -1 0 12328 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0770_
timestamp 1688980957
transform 1 0 12144 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0771_
timestamp 1688980957
transform -1 0 13984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0772_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0773_
timestamp 1688980957
transform -1 0 11960 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _0774_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13616 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o311a_1  _0775_
timestamp 1688980957
transform -1 0 14352 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0776_
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0777_
timestamp 1688980957
transform -1 0 12328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0778_
timestamp 1688980957
transform -1 0 10212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0779_
timestamp 1688980957
transform 1 0 9568 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0780_
timestamp 1688980957
transform 1 0 10304 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _0781_
timestamp 1688980957
transform -1 0 12052 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _0782_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13432 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _0783_
timestamp 1688980957
transform 1 0 17848 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0784_
timestamp 1688980957
transform 1 0 18676 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _0785_
timestamp 1688980957
transform 1 0 22632 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0786_
timestamp 1688980957
transform 1 0 23276 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _0787_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0788_
timestamp 1688980957
transform -1 0 23828 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0789_
timestamp 1688980957
transform -1 0 22908 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1688980957
transform -1 0 23184 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0791_
timestamp 1688980957
transform 1 0 21988 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0792_
timestamp 1688980957
transform 1 0 22448 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0793_
timestamp 1688980957
transform 1 0 22356 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0794_
timestamp 1688980957
transform 1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0795_
timestamp 1688980957
transform 1 0 22632 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _0796_
timestamp 1688980957
transform -1 0 23092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0797_
timestamp 1688980957
transform 1 0 12328 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0798_
timestamp 1688980957
transform -1 0 13340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _0799_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0800_
timestamp 1688980957
transform 1 0 11776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _0801_
timestamp 1688980957
transform 1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _0802_
timestamp 1688980957
transform -1 0 13248 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_1  _0803_
timestamp 1688980957
transform -1 0 13248 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0804_
timestamp 1688980957
transform 1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0805_
timestamp 1688980957
transform 1 0 19688 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _0806_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _0807_
timestamp 1688980957
transform -1 0 21344 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _0808_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20792 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0809_
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0810_
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _0811_
timestamp 1688980957
transform 1 0 20792 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _0812_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20792 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0813_
timestamp 1688980957
transform -1 0 20056 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1688980957
transform -1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0815_
timestamp 1688980957
transform 1 0 15272 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _0816_
timestamp 1688980957
transform -1 0 16192 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _0817_
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0818_
timestamp 1688980957
transform 1 0 12880 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0819_
timestamp 1688980957
transform 1 0 12788 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0820_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a41o_1  _0821_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0823_
timestamp 1688980957
transform -1 0 21344 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a211oi_1  _0824_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0825_
timestamp 1688980957
transform -1 0 17572 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0826_
timestamp 1688980957
transform 1 0 16376 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0827_
timestamp 1688980957
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0828_
timestamp 1688980957
transform -1 0 16100 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _0829_
timestamp 1688980957
transform -1 0 15640 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _0830_
timestamp 1688980957
transform 1 0 16008 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0831_
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0832_
timestamp 1688980957
transform 1 0 17204 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0833_
timestamp 1688980957
transform -1 0 20884 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0834_
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0835_
timestamp 1688980957
transform -1 0 17940 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0836_
timestamp 1688980957
transform 1 0 17204 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _0837_
timestamp 1688980957
transform -1 0 18768 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0838_
timestamp 1688980957
transform 1 0 15272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0839_
timestamp 1688980957
transform 1 0 15548 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0840_
timestamp 1688980957
transform 1 0 15272 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0841_
timestamp 1688980957
transform 1 0 11960 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0842_
timestamp 1688980957
transform 1 0 11684 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0843_
timestamp 1688980957
transform -1 0 12604 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _0844_
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a41o_1  _0845_
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _0846_
timestamp 1688980957
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _0847_
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0848_
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a41o_1  _0849_
timestamp 1688980957
transform 1 0 10488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1688980957
transform -1 0 12052 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0851_
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0852_
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _0853_
timestamp 1688980957
transform 1 0 15640 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0854_
timestamp 1688980957
transform 1 0 16468 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _0855_
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0856_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21252 0 1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_1  _0857_
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0858_
timestamp 1688980957
transform 1 0 21896 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0859_
timestamp 1688980957
transform 1 0 22080 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _0860_
timestamp 1688980957
transform 1 0 21160 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0861_
timestamp 1688980957
transform 1 0 23000 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0862_
timestamp 1688980957
transform 1 0 22172 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _0863_
timestamp 1688980957
transform -1 0 24288 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a311oi_4  _0864_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_2  _0865_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25392 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _0866_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0867_
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0868_
timestamp 1688980957
transform -1 0 19688 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0869_
timestamp 1688980957
transform 1 0 18400 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0870_
timestamp 1688980957
transform 1 0 23368 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0871_
timestamp 1688980957
transform 1 0 23828 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0872_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _0873_
timestamp 1688980957
transform -1 0 27968 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_2  _0874_
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0875_
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0876_
timestamp 1688980957
transform -1 0 22356 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0877_
timestamp 1688980957
transform -1 0 22448 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o2111ai_4  _0878_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__and3_1  _0879_
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0880_
timestamp 1688980957
transform -1 0 24932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0881_
timestamp 1688980957
transform 1 0 25576 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1688980957
transform -1 0 23276 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0883_
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0884_
timestamp 1688980957
transform 1 0 24932 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0885_
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0886_
timestamp 1688980957
transform 1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0887_
timestamp 1688980957
transform 1 0 23736 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0888_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_1  _0889_
timestamp 1688980957
transform 1 0 24840 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0890_
timestamp 1688980957
transform -1 0 25944 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0891_
timestamp 1688980957
transform 1 0 24472 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0892_
timestamp 1688980957
transform 1 0 25300 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a41oi_4  _0893_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27600 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _0894_
timestamp 1688980957
transform 1 0 27968 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0895_
timestamp 1688980957
transform 1 0 22632 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0896_
timestamp 1688980957
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0897_
timestamp 1688980957
transform -1 0 26404 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0898_
timestamp 1688980957
transform 1 0 25944 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _0899_
timestamp 1688980957
transform 1 0 26680 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0900_
timestamp 1688980957
transform -1 0 27140 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor3b_1  _0901_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27508 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _0902_
timestamp 1688980957
transform -1 0 24196 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _0903_
timestamp 1688980957
transform 1 0 22816 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1688980957
transform 1 0 27324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _0905_
timestamp 1688980957
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _0906_
timestamp 1688980957
transform -1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _0907_
timestamp 1688980957
transform 1 0 27692 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0908_
timestamp 1688980957
transform 1 0 23736 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0909_
timestamp 1688980957
transform 1 0 27232 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0910_
timestamp 1688980957
transform 1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0911_
timestamp 1688980957
transform 1 0 20608 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _0912_
timestamp 1688980957
transform 1 0 27232 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0913_
timestamp 1688980957
transform 1 0 27600 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0914_
timestamp 1688980957
transform -1 0 27600 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0915_
timestamp 1688980957
transform -1 0 28612 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0916_
timestamp 1688980957
transform -1 0 28796 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _0917_
timestamp 1688980957
transform 1 0 23092 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0918_
timestamp 1688980957
transform -1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0919_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0920_
timestamp 1688980957
transform 1 0 27600 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0921_
timestamp 1688980957
transform -1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a221oi_4  _0922_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27324 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_1  _0923_
timestamp 1688980957
transform -1 0 27876 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0925_
timestamp 1688980957
transform -1 0 26680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0926_
timestamp 1688980957
transform 1 0 23920 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _0927_
timestamp 1688980957
transform -1 0 25576 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0928_
timestamp 1688980957
transform 1 0 24748 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _0929_
timestamp 1688980957
transform -1 0 25668 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0930_
timestamp 1688980957
transform 1 0 25668 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0931_
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0932_
timestamp 1688980957
transform 1 0 20240 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0933_
timestamp 1688980957
transform 1 0 21068 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_1  _0934_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0935_
timestamp 1688980957
transform 1 0 27324 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0936_
timestamp 1688980957
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _0937_
timestamp 1688980957
transform 1 0 18584 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0938_
timestamp 1688980957
transform -1 0 19504 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0939_
timestamp 1688980957
transform 1 0 19504 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0940_
timestamp 1688980957
transform -1 0 19320 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_2  _0941_
timestamp 1688980957
transform -1 0 24840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _0942_
timestamp 1688980957
transform 1 0 25668 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0943_
timestamp 1688980957
transform -1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _0944_
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _0945_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _0946_
timestamp 1688980957
transform 1 0 20424 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0947_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _0948_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26312 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _0949_
timestamp 1688980957
transform -1 0 25760 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0950_
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0951_
timestamp 1688980957
transform -1 0 19136 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0952_
timestamp 1688980957
transform -1 0 20976 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0953_
timestamp 1688980957
transform -1 0 20976 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0954_
timestamp 1688980957
transform 1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _0955_
timestamp 1688980957
transform 1 0 17480 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0956_
timestamp 1688980957
transform 1 0 16744 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0957_
timestamp 1688980957
transform 1 0 17572 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0958_
timestamp 1688980957
transform 1 0 17020 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0959_
timestamp 1688980957
transform 1 0 16928 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0960_
timestamp 1688980957
transform 1 0 16744 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_2  _0961_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0962_
timestamp 1688980957
transform 1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _0963_
timestamp 1688980957
transform -1 0 18216 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _0964_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18584 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _0965_
timestamp 1688980957
transform 1 0 20240 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0966_
timestamp 1688980957
transform -1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0967_
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0968_
timestamp 1688980957
transform 1 0 20148 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0969_
timestamp 1688980957
transform -1 0 21252 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0970_
timestamp 1688980957
transform -1 0 21068 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_2  _0971_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21436 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0972_
timestamp 1688980957
transform 1 0 22356 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0973_
timestamp 1688980957
transform 1 0 21896 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _0974_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _0975_
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0976_
timestamp 1688980957
transform 1 0 22356 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0977_
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _0978_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22448 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _0979_
timestamp 1688980957
transform 1 0 23368 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0980_
timestamp 1688980957
transform 1 0 22356 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _0981_
timestamp 1688980957
transform -1 0 23644 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0982_
timestamp 1688980957
transform 1 0 23460 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0983_
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0984_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0985_
timestamp 1688980957
transform -1 0 12788 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0986_
timestamp 1688980957
transform 1 0 12788 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0987_
timestamp 1688980957
transform -1 0 14720 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0988_
timestamp 1688980957
transform -1 0 14904 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0989_
timestamp 1688980957
transform 1 0 14628 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0990_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14628 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0992_
timestamp 1688980957
transform 1 0 22356 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0993_
timestamp 1688980957
transform 1 0 23092 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__o2111a_1  _0994_
timestamp 1688980957
transform 1 0 24932 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__a311o_1  _0995_
timestamp 1688980957
transform 1 0 24564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _0996_
timestamp 1688980957
transform -1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_2  _0997_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24932 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o2111ai_4  _0998_
timestamp 1688980957
transform 1 0 24840 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__o2111a_1  _0999_
timestamp 1688980957
transform -1 0 24656 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_2  _1000_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23368 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1001_
timestamp 1688980957
transform -1 0 24564 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1002_
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1003_
timestamp 1688980957
transform 1 0 16744 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1004_
timestamp 1688980957
transform 1 0 23184 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1688980957
transform -1 0 23552 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1006_
timestamp 1688980957
transform -1 0 23828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _1007_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24932 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1008_
timestamp 1688980957
transform 1 0 23368 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1009_
timestamp 1688980957
transform 1 0 19320 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1010_
timestamp 1688980957
transform -1 0 19044 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1011_
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _1012_
timestamp 1688980957
transform 1 0 22264 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1013_
timestamp 1688980957
transform 1 0 20792 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _1014_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1015_
timestamp 1688980957
transform 1 0 22080 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1016_
timestamp 1688980957
transform -1 0 20792 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1017_
timestamp 1688980957
transform 1 0 20424 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1018_
timestamp 1688980957
transform -1 0 20608 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o221ai_1  _1019_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1020_
timestamp 1688980957
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1021_
timestamp 1688980957
transform 1 0 22264 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _1022_
timestamp 1688980957
transform -1 0 22264 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1023_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1024_
timestamp 1688980957
transform 1 0 20976 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1025_
timestamp 1688980957
transform 1 0 22356 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1026_
timestamp 1688980957
transform 1 0 23828 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1027_
timestamp 1688980957
transform 1 0 24656 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1028_
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1029_
timestamp 1688980957
transform -1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1030_
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1031_
timestamp 1688980957
transform 1 0 25208 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1032_
timestamp 1688980957
transform -1 0 24840 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1033_
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1034_
timestamp 1688980957
transform 1 0 26772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1035_
timestamp 1688980957
transform -1 0 26772 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1036_
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1037_
timestamp 1688980957
transform -1 0 26496 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1038_
timestamp 1688980957
transform 1 0 25208 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1039_
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1040_
timestamp 1688980957
transform 1 0 28244 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _1041_
timestamp 1688980957
transform 1 0 28152 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1042_
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1043_
timestamp 1688980957
transform -1 0 27140 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1044_
timestamp 1688980957
transform 1 0 26036 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1045_
timestamp 1688980957
transform 1 0 27140 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1046_
timestamp 1688980957
transform 1 0 27324 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1047_
timestamp 1688980957
transform 1 0 27968 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1048_
timestamp 1688980957
transform -1 0 20700 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1688980957
transform -1 0 20976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1050_
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1051_
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1052_
timestamp 1688980957
transform 1 0 20240 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1053_
timestamp 1688980957
transform 1 0 20700 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1054_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1055_
timestamp 1688980957
transform -1 0 21436 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1056_
timestamp 1688980957
transform 1 0 28612 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1057_
timestamp 1688980957
transform 1 0 27416 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1058_
timestamp 1688980957
transform 1 0 27968 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1059_
timestamp 1688980957
transform -1 0 27876 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1060_
timestamp 1688980957
transform -1 0 28888 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1061_
timestamp 1688980957
transform 1 0 28060 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1062_
timestamp 1688980957
transform 1 0 28612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1063_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1064_
timestamp 1688980957
transform -1 0 30820 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  _1065_
timestamp 1688980957
transform -1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  _1066_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9292 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1688980957
transform 1 0 27140 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1068_
timestamp 1688980957
transform -1 0 29072 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1069_
timestamp 1688980957
transform 1 0 25852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1070_
timestamp 1688980957
transform -1 0 29992 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1071_
timestamp 1688980957
transform 1 0 27508 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1072_
timestamp 1688980957
transform -1 0 29900 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1073_
timestamp 1688980957
transform -1 0 30636 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1074_
timestamp 1688980957
transform -1 0 29808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1075_
timestamp 1688980957
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1077_
timestamp 1688980957
transform 1 0 30820 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1078_
timestamp 1688980957
transform 1 0 30636 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1079_
timestamp 1688980957
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1688980957
transform -1 0 30820 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1081_
timestamp 1688980957
transform 1 0 29992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1082_
timestamp 1688980957
transform -1 0 31096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1083_
timestamp 1688980957
transform 1 0 9476 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1084_
timestamp 1688980957
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1085_
timestamp 1688980957
transform 1 0 9384 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1086_
timestamp 1688980957
transform 1 0 26404 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1087_
timestamp 1688980957
transform 1 0 9844 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1088_
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1089_
timestamp 1688980957
transform -1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1688980957
transform -1 0 7544 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1091_
timestamp 1688980957
transform -1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1092_
timestamp 1688980957
transform -1 0 8832 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1688980957
transform -1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1688980957
transform 1 0 7268 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1095_
timestamp 1688980957
transform 1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1096_
timestamp 1688980957
transform -1 0 8464 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1097_
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1098_
timestamp 1688980957
transform 1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1099_
timestamp 1688980957
transform -1 0 9752 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1100_
timestamp 1688980957
transform -1 0 34592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1101_
timestamp 1688980957
transform 1 0 33396 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1103_
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1104_
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1105_
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1106_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1688980957
transform 1 0 33856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1688980957
transform 1 0 33672 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1109_
timestamp 1688980957
transform 1 0 33212 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1110_
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1111_
timestamp 1688980957
transform 1 0 33396 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1112_
timestamp 1688980957
transform -1 0 34224 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1113_
timestamp 1688980957
transform -1 0 34500 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1114_
timestamp 1688980957
transform 1 0 33580 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1115_
timestamp 1688980957
transform -1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1116_
timestamp 1688980957
transform -1 0 33488 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1117_
timestamp 1688980957
transform -1 0 4048 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1688980957
transform -1 0 3496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1119_
timestamp 1688980957
transform -1 0 2576 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1688980957
transform -1 0 3496 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1121_
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1123_
timestamp 1688980957
transform 1 0 4048 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1688980957
transform -1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1125_
timestamp 1688980957
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1126_
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1127_
timestamp 1688980957
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1128_
timestamp 1688980957
transform -1 0 3496 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1688980957
transform 1 0 2208 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1130_
timestamp 1688980957
transform -1 0 4140 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1688980957
transform 1 0 4600 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1132_
timestamp 1688980957
transform -1 0 2024 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1133_
timestamp 1688980957
transform -1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _1134_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1135_
timestamp 1688980957
transform 1 0 27048 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1136_
timestamp 1688980957
transform 1 0 24932 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1137_
timestamp 1688980957
transform 1 0 27876 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1138_
timestamp 1688980957
transform 1 0 26496 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1139_
timestamp 1688980957
transform 1 0 27784 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1140_
timestamp 1688980957
transform 1 0 28520 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1141_
timestamp 1688980957
transform 1 0 28428 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1142_
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1143_
timestamp 1688980957
transform 1 0 29348 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1144_
timestamp 1688980957
transform 1 0 29992 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1145_
timestamp 1688980957
transform 1 0 29716 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1146_
timestamp 1688980957
transform 1 0 28520 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1147_
timestamp 1688980957
transform 1 0 28704 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1148_
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1149_
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1150_ unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1151_
timestamp 1688980957
transform 1 0 6532 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1152_
timestamp 1688980957
transform 1 0 8372 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1153_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1154_
timestamp 1688980957
transform 1 0 6164 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1155_
timestamp 1688980957
transform 1 0 7176 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1156_
timestamp 1688980957
transform 1 0 6164 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1157_
timestamp 1688980957
transform 1 0 6992 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1158_
timestamp 1688980957
transform 1 0 6716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1159_
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1160_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1161_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1162_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1163_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1164_
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1165_
timestamp 1688980957
transform 1 0 7636 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1166_
timestamp 1688980957
transform 1 0 32752 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1167_
timestamp 1688980957
transform 1 0 32476 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1168_
timestamp 1688980957
transform 1 0 32752 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1169_
timestamp 1688980957
transform 1 0 32752 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1170_
timestamp 1688980957
transform 1 0 32752 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1171_
timestamp 1688980957
transform 1 0 33120 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1172_
timestamp 1688980957
transform 1 0 32936 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1173_
timestamp 1688980957
transform 1 0 32752 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1174_
timestamp 1688980957
transform 1 0 32200 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1175_
timestamp 1688980957
transform 1 0 32292 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1176_
timestamp 1688980957
transform 1 0 32384 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1177_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1178_
timestamp 1688980957
transform 1 0 32752 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1179_
timestamp 1688980957
transform 1 0 32660 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1180_
timestamp 1688980957
transform 1 0 32752 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1181_
timestamp 1688980957
transform 1 0 31372 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1182_
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1183_
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1184_
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1185_
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1186_
timestamp 1688980957
transform 1 0 2300 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1187_
timestamp 1688980957
transform 1 0 1840 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1188_
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1189_
timestamp 1688980957
transform 1 0 1564 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1190_
timestamp 1688980957
transform 1 0 1840 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1191_
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1192_
timestamp 1688980957
transform 1 0 1840 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1193_
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1194_
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1195_
timestamp 1688980957
transform 1 0 2024 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1196_
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1197_
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1198_
timestamp 1688980957
transform 1 0 1564 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B1 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__A
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__B1
timestamp 1688980957
transform -1 0 3496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__C1
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__B1
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1688980957
transform 1 0 4416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__B1
timestamp 1688980957
transform 1 0 4876 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1688980957
transform 1 0 4508 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__B1
timestamp 1688980957
transform 1 0 4232 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1688980957
transform 1 0 6072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__C1
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__B1
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A
timestamp 1688980957
transform -1 0 6900 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A
timestamp 1688980957
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B1
timestamp 1688980957
transform 1 0 29992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__B1
timestamp 1688980957
transform 1 0 30636 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1688980957
transform 1 0 31280 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1688980957
transform 1 0 31280 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__B1
timestamp 1688980957
transform 1 0 31464 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1688980957
transform 1 0 31832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A
timestamp 1688980957
transform 1 0 31556 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B1
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 1688980957
transform 1 0 32476 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1688980957
transform -1 0 33028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__B1
timestamp 1688980957
transform 1 0 32292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1688980957
transform 1 0 31556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B1
timestamp 1688980957
transform 1 0 31188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__B1
timestamp 1688980957
transform 1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B
timestamp 1688980957
transform 1 0 32476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__B
timestamp 1688980957
transform 1 0 18216 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__B
timestamp 1688980957
transform 1 0 16008 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__C
timestamp 1688980957
transform 1 0 16100 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__D
timestamp 1688980957
transform 1 0 17480 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A
timestamp 1688980957
transform 1 0 15640 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__B
timestamp 1688980957
transform -1 0 15640 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__C
timestamp 1688980957
transform 1 0 15272 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__D
timestamp 1688980957
transform -1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1688980957
transform 1 0 16928 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__C
timestamp 1688980957
transform 1 0 17296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__D
timestamp 1688980957
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1688980957
transform -1 0 10764 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__B
timestamp 1688980957
transform 1 0 11132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1688980957
transform 1 0 10396 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B
timestamp 1688980957
transform 1 0 10212 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__B
timestamp 1688980957
transform 1 0 11960 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__B
timestamp 1688980957
transform 1 0 11960 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B
timestamp 1688980957
transform 1 0 19320 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1688980957
transform 1 0 19872 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1688980957
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1688980957
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1688980957
transform -1 0 14720 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A
timestamp 1688980957
transform 1 0 14444 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B
timestamp 1688980957
transform 1 0 14076 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A
timestamp 1688980957
transform 1 0 14720 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__B
timestamp 1688980957
transform -1 0 15180 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A
timestamp 1688980957
transform 1 0 12788 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__B
timestamp 1688980957
transform 1 0 12420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A1
timestamp 1688980957
transform 1 0 13524 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__B2
timestamp 1688980957
transform -1 0 14536 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__B1
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__C1
timestamp 1688980957
transform 1 0 17572 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B
timestamp 1688980957
transform 1 0 17848 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1688980957
transform 1 0 18124 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1688980957
transform 1 0 17572 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1688980957
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A
timestamp 1688980957
transform 1 0 20424 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B
timestamp 1688980957
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1688980957
transform -1 0 16008 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B
timestamp 1688980957
transform 1 0 15640 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A1
timestamp 1688980957
transform 1 0 16284 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A2
timestamp 1688980957
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1688980957
transform 1 0 11776 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1688980957
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1688980957
transform -1 0 11408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B
timestamp 1688980957
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1688980957
transform -1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__B
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1688980957
transform 1 0 10764 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B
timestamp 1688980957
transform 1 0 10396 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1688980957
transform -1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B
timestamp 1688980957
transform -1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__C
timestamp 1688980957
transform -1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__D
timestamp 1688980957
transform -1 0 10580 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1688980957
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__C
timestamp 1688980957
transform 1 0 11592 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__D
timestamp 1688980957
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1688980957
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1688980957
transform 1 0 18216 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 1688980957
transform 1 0 17848 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1688980957
transform 1 0 14536 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1688980957
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1688980957
transform 1 0 13248 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1688980957
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A
timestamp 1688980957
transform -1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B
timestamp 1688980957
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A
timestamp 1688980957
transform -1 0 17848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A1
timestamp 1688980957
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A2
timestamp 1688980957
transform 1 0 16928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B1
timestamp 1688980957
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B2
timestamp 1688980957
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A
timestamp 1688980957
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B
timestamp 1688980957
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__C
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__D
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp 1688980957
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__C
timestamp 1688980957
transform -1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__D
timestamp 1688980957
transform 1 0 18768 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1688980957
transform 1 0 18860 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1688980957
transform -1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B
timestamp 1688980957
transform 1 0 19596 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A1
timestamp 1688980957
transform -1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1688980957
transform 1 0 20056 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 1688980957
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1688980957
transform 1 0 13432 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1688980957
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1688980957
transform 1 0 13064 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1688980957
transform 1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1688980957
transform 1 0 14628 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__C1
timestamp 1688980957
transform -1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1688980957
transform 1 0 9292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B
timestamp 1688980957
transform -1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 1688980957
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B1
timestamp 1688980957
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__C1
timestamp 1688980957
transform -1 0 14444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1
timestamp 1688980957
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1688980957
transform 1 0 16284 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B
timestamp 1688980957
transform 1 0 15456 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B
timestamp 1688980957
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1688980957
transform 1 0 15364 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1688980957
transform 1 0 14444 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__B
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__C_N
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B
timestamp 1688980957
transform 1 0 10212 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B
timestamp 1688980957
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1688980957
transform 1 0 13524 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B
timestamp 1688980957
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2
timestamp 1688980957
transform 1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A
timestamp 1688980957
transform -1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B
timestamp 1688980957
transform 1 0 11132 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1
timestamp 1688980957
transform 1 0 12420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A2
timestamp 1688980957
transform 1 0 12052 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A
timestamp 1688980957
transform 1 0 9752 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B
timestamp 1688980957
transform 1 0 9568 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1688980957
transform 1 0 9568 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__B
timestamp 1688980957
transform -1 0 8832 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__C
timestamp 1688980957
transform -1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__D
timestamp 1688980957
transform -1 0 9568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A2
timestamp 1688980957
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1688980957
transform -1 0 23368 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__B
timestamp 1688980957
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1688980957
transform 1 0 23460 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1688980957
transform 1 0 22448 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B
timestamp 1688980957
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B
timestamp 1688980957
transform 1 0 23368 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1688980957
transform 1 0 22172 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B
timestamp 1688980957
transform 1 0 21988 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A
timestamp 1688980957
transform -1 0 23368 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1688980957
transform 1 0 10672 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B
timestamp 1688980957
transform 1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1688980957
transform 1 0 12696 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A_N
timestamp 1688980957
transform 1 0 9844 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1688980957
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A1
timestamp 1688980957
transform 1 0 13524 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A1
timestamp 1688980957
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B
timestamp 1688980957
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A_N
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B
timestamp 1688980957
transform 1 0 21252 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A1
timestamp 1688980957
transform 1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A2
timestamp 1688980957
transform 1 0 20148 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__B1_N
timestamp 1688980957
transform -1 0 21712 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A_N
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B
timestamp 1688980957
transform 1 0 17940 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__C
timestamp 1688980957
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1688980957
transform 1 0 19780 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__C1
timestamp 1688980957
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B
timestamp 1688980957
transform -1 0 15088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B
timestamp 1688980957
transform 1 0 15088 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1688980957
transform -1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__B
timestamp 1688980957
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A1
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B1
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A1
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1688980957
transform 1 0 11316 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A
timestamp 1688980957
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__C
timestamp 1688980957
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__D
timestamp 1688980957
transform 1 0 10488 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1688980957
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1688980957
transform 1 0 21988 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__B
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__C
timestamp 1688980957
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__D
timestamp 1688980957
transform 1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1688980957
transform 1 0 23092 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__C
timestamp 1688980957
transform 1 0 21620 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__D
timestamp 1688980957
transform 1 0 22724 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1688980957
transform 1 0 21620 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B
timestamp 1688980957
transform 1 0 21528 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__B
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A
timestamp 1688980957
transform -1 0 22908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__C1
timestamp 1688980957
transform 1 0 23552 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__D1
timestamp 1688980957
transform 1 0 23828 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A1
timestamp 1688980957
transform 1 0 25024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A2
timestamp 1688980957
transform -1 0 25576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1688980957
transform 1 0 23552 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__B
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__C
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__D
timestamp 1688980957
transform 1 0 23184 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1688980957
transform 1 0 18032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B
timestamp 1688980957
transform -1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1688980957
transform 1 0 19872 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B
timestamp 1688980957
transform 1 0 18400 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A
timestamp 1688980957
transform -1 0 23552 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B
timestamp 1688980957
transform -1 0 23184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1688980957
transform -1 0 24564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1688980957
transform -1 0 24196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A
timestamp 1688980957
transform 1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B
timestamp 1688980957
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1688980957
transform -1 0 22172 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B
timestamp 1688980957
transform 1 0 23460 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1688980957
transform 1 0 21896 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A1
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A3
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1688980957
transform -1 0 25576 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__B
timestamp 1688980957
transform -1 0 24932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1688980957
transform -1 0 23276 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__B
timestamp 1688980957
transform 1 0 24196 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1688980957
transform 1 0 23276 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__B
timestamp 1688980957
transform 1 0 23092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1688980957
transform 1 0 23644 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A1
timestamp 1688980957
transform -1 0 24472 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A
timestamp 1688980957
transform -1 0 25760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B
timestamp 1688980957
transform -1 0 25208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__C
timestamp 1688980957
transform -1 0 24748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__D
timestamp 1688980957
transform 1 0 24656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A1
timestamp 1688980957
transform 1 0 23920 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1688980957
transform 1 0 24012 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1688980957
transform 1 0 21252 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1688980957
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1688980957
transform -1 0 24748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B
timestamp 1688980957
transform 1 0 23552 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__B
timestamp 1688980957
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A2
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A3
timestamp 1688980957
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A4
timestamp 1688980957
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1688980957
transform 1 0 16560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__B
timestamp 1688980957
transform 1 0 16192 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B1
timestamp 1688980957
transform 1 0 17480 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__C1
timestamp 1688980957
transform -1 0 17480 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A1
timestamp 1688980957
transform 1 0 13156 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__B
timestamp 1688980957
transform 1 0 12972 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__B2
timestamp 1688980957
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A1_N
timestamp 1688980957
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A2_N
timestamp 1688980957
transform 1 0 13432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1688980957
transform -1 0 23552 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1688980957
transform 1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1688980957
transform 1 0 22172 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B
timestamp 1688980957
transform 1 0 21988 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A1
timestamp 1688980957
transform -1 0 18676 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A2
timestamp 1688980957
transform -1 0 18308 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1688980957
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__B
timestamp 1688980957
transform 1 0 20056 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A
timestamp 1688980957
transform 1 0 21252 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1688980957
transform 1 0 21160 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1688980957
transform 1 0 20700 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__C
timestamp 1688980957
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1
timestamp 1688980957
transform 1 0 22172 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A1
timestamp 1688980957
transform 1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1688980957
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A
timestamp 1688980957
transform -1 0 27140 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A
timestamp 1688980957
transform 1 0 29256 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A
timestamp 1688980957
transform 1 0 25668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1688980957
transform 1 0 30176 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A
timestamp 1688980957
transform 1 0 27324 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A
timestamp 1688980957
transform 1 0 30084 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A
timestamp 1688980957
transform 1 0 30820 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1688980957
transform 1 0 29992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1688980957
transform 1 0 29992 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A
timestamp 1688980957
transform 1 0 30728 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1688980957
transform 1 0 30452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A
timestamp 1688980957
transform 1 0 28980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A
timestamp 1688980957
transform 1 0 30360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1688980957
transform 1 0 29808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1688980957
transform -1 0 31464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__A
timestamp 1688980957
transform 1 0 9936 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__A
timestamp 1688980957
transform -1 0 8832 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A
timestamp 1688980957
transform 1 0 9752 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A
timestamp 1688980957
transform 1 0 28428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__A
timestamp 1688980957
transform 1 0 10304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__A
timestamp 1688980957
transform -1 0 6900 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__A
timestamp 1688980957
transform 1 0 9292 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__A
timestamp 1688980957
transform 1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1688980957
transform -1 0 9016 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__A
timestamp 1688980957
transform 1 0 8556 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__A
timestamp 1688980957
transform 1 0 7728 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1688980957
transform 1 0 7728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__A
timestamp 1688980957
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__A
timestamp 1688980957
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A
timestamp 1688980957
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A
timestamp 1688980957
transform 1 0 9936 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__A
timestamp 1688980957
transform -1 0 34960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__A
timestamp 1688980957
transform 1 0 33856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__A
timestamp 1688980957
transform 1 0 34500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1688980957
transform 1 0 34132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__A
timestamp 1688980957
transform 1 0 34500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__A
timestamp 1688980957
transform 1 0 33856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A
timestamp 1688980957
transform -1 0 29164 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1688980957
transform 1 0 33672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1688980957
transform 1 0 33488 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1688980957
transform 1 0 33028 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1688980957
transform 1 0 33028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A
timestamp 1688980957
transform 1 0 33212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A
timestamp 1688980957
transform -1 0 34868 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1688980957
transform 1 0 34408 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1688980957
transform 1 0 32660 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1688980957
transform -1 0 34868 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A
timestamp 1688980957
transform 1 0 33028 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__A
timestamp 1688980957
transform 1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1688980957
transform 1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1688980957
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A
timestamp 1688980957
transform 1 0 2668 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1688980957
transform 1 0 4508 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__A
timestamp 1688980957
transform 1 0 4048 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1688980957
transform 1 0 4232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1688980957
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1688980957
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__A
timestamp 1688980957
transform 1 0 2668 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1688980957
transform 1 0 4324 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1688980957
transform 1 0 5060 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1688980957
transform 1 0 2024 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__A
timestamp 1688980957
transform 1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__CLK
timestamp 1688980957
transform 1 0 26680 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__CLK
timestamp 1688980957
transform 1 0 26864 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__CLK
timestamp 1688980957
transform 1 0 24748 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__CLK
timestamp 1688980957
transform 1 0 27692 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__CLK
timestamp 1688980957
transform 1 0 26312 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__CLK
timestamp 1688980957
transform 1 0 27600 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__CLK
timestamp 1688980957
transform 1 0 28336 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__CLK
timestamp 1688980957
transform 1 0 28244 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__CLK
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__CLK
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1688980957
transform 1 0 29808 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1688980957
transform 1 0 29532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1688980957
transform 1 0 28336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__CLK
timestamp 1688980957
transform 1 0 28520 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1688980957
transform 1 0 29348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1688980957
transform 1 0 29256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1688980957
transform 1 0 8372 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__CLK
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1688980957
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__CLK
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__CLK
timestamp 1688980957
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__CLK
timestamp 1688980957
transform 1 0 8464 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__CLK
timestamp 1688980957
transform 1 0 7820 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__CLK
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1688980957
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__CLK
timestamp 1688980957
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1688980957
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__CLK
timestamp 1688980957
transform 1 0 9476 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__CLK
timestamp 1688980957
transform 1 0 32568 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__CLK
timestamp 1688980957
transform 1 0 32568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__CLK
timestamp 1688980957
transform 1 0 32936 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__CLK
timestamp 1688980957
transform 1 0 32568 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1688980957
transform 1 0 32936 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__CLK
timestamp 1688980957
transform 1 0 32752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__CLK
timestamp 1688980957
transform 1 0 32568 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1688980957
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1688980957
transform 1 0 31832 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1688980957
transform 1 0 31924 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1688980957
transform 1 0 32568 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__CLK
timestamp 1688980957
transform 1 0 32476 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1688980957
transform 1 0 32568 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1688980957
transform 1 0 31648 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1688980957
transform 1 0 4508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__CLK
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__CLK
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1688980957
transform 1 0 4140 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1688980957
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1688980957
transform 1 0 5796 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1688980957
transform 1 0 3680 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1688980957
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1688980957
transform 1 0 4048 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1688980957
transform 1 0 3404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1688980957
transform 1 0 3956 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1688980957
transform 1 0 5796 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1688980957
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_281 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_288
timestamp 1688980957
transform 1 0 27600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_300
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_367
timestamp 1688980957
transform 1 0 34868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_367
timestamp 1688980957
transform 1 0 34868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_367
timestamp 1688980957
transform 1 0 34868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_367
timestamp 1688980957
transform 1 0 34868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 1688980957
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1688980957
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_341
timestamp 1688980957
transform 1 0 32476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_364
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_237
timestamp 1688980957
transform 1 0 22908 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_240
timestamp 1688980957
transform 1 0 23184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_244
timestamp 1688980957
transform 1 0 23552 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_295
timestamp 1688980957
transform 1 0 28244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_299
timestamp 1688980957
transform 1 0 28612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_348
timestamp 1688980957
transform 1 0 33120 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_354
timestamp 1688980957
transform 1 0 33672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_358
timestamp 1688980957
transform 1 0 34040 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_20
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_24
timestamp 1688980957
transform 1 0 3312 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_36
timestamp 1688980957
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_48
timestamp 1688980957
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_185
timestamp 1688980957
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_188
timestamp 1688980957
transform 1 0 18400 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_200
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_212
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_229
timestamp 1688980957
transform 1 0 22172 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_233
timestamp 1688980957
transform 1 0 22540 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_241
timestamp 1688980957
transform 1 0 23276 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_247
timestamp 1688980957
transform 1 0 23828 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_251
timestamp 1688980957
transform 1 0 24196 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_255
timestamp 1688980957
transform 1 0 24564 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_259
timestamp 1688980957
transform 1 0 24932 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_271
timestamp 1688980957
transform 1 0 26036 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_288
timestamp 1688980957
transform 1 0 27600 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_318
timestamp 1688980957
transform 1 0 30360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_330
timestamp 1688980957
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_347
timestamp 1688980957
transform 1 0 33028 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_351
timestamp 1688980957
transform 1 0 33396 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_33
timestamp 1688980957
transform 1 0 4140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_45
timestamp 1688980957
transform 1 0 5244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_57
timestamp 1688980957
transform 1 0 6348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_69
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_183
timestamp 1688980957
transform 1 0 17940 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_186
timestamp 1688980957
transform 1 0 18216 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_202
timestamp 1688980957
transform 1 0 19688 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_206
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_216
timestamp 1688980957
transform 1 0 20976 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_220
timestamp 1688980957
transform 1 0 21344 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_224
timestamp 1688980957
transform 1 0 21712 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_228
timestamp 1688980957
transform 1 0 22080 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_234
timestamp 1688980957
transform 1 0 22632 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_238
timestamp 1688980957
transform 1 0 23000 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_242
timestamp 1688980957
transform 1 0 23368 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_246
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_258
timestamp 1688980957
transform 1 0 24840 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_262
timestamp 1688980957
transform 1 0 25208 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_266
timestamp 1688980957
transform 1 0 25576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_299
timestamp 1688980957
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_339
timestamp 1688980957
transform 1 0 32292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_343
timestamp 1688980957
transform 1 0 32660 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_117
timestamp 1688980957
transform 1 0 11868 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_129
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_141
timestamp 1688980957
transform 1 0 14076 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_153
timestamp 1688980957
transform 1 0 15180 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1688980957
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_187
timestamp 1688980957
transform 1 0 18308 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_216
timestamp 1688980957
transform 1 0 20976 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_231
timestamp 1688980957
transform 1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_241
timestamp 1688980957
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_245
timestamp 1688980957
transform 1 0 23644 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_253
timestamp 1688980957
transform 1 0 24380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 1688980957
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_287
timestamp 1688980957
transform 1 0 27508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_299
timestamp 1688980957
transform 1 0 28612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_309
timestamp 1688980957
transform 1 0 29532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_325
timestamp 1688980957
transform 1 0 31004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_341
timestamp 1688980957
transform 1 0 32476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_344
timestamp 1688980957
transform 1 0 32752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_348
timestamp 1688980957
transform 1 0 33120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_356
timestamp 1688980957
transform 1 0 33856 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_365
timestamp 1688980957
transform 1 0 34684 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 1688980957
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 1688980957
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1688980957
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_93
timestamp 1688980957
transform 1 0 9660 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_129
timestamp 1688980957
transform 1 0 12972 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1688980957
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_187
timestamp 1688980957
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_191
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_205
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_208
timestamp 1688980957
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_217
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_225
timestamp 1688980957
transform 1 0 21804 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_231
timestamp 1688980957
transform 1 0 22356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_235
timestamp 1688980957
transform 1 0 22724 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_274
timestamp 1688980957
transform 1 0 26312 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_283
timestamp 1688980957
transform 1 0 27140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_291
timestamp 1688980957
transform 1 0 27876 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_300
timestamp 1688980957
transform 1 0 28704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_317
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_320
timestamp 1688980957
transform 1 0 30544 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_341
timestamp 1688980957
transform 1 0 32476 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_35
timestamp 1688980957
transform 1 0 4324 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_94
timestamp 1688980957
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_107
timestamp 1688980957
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_131
timestamp 1688980957
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_140
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_152
timestamp 1688980957
transform 1 0 15088 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_160
timestamp 1688980957
transform 1 0 15824 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_178
timestamp 1688980957
transform 1 0 17480 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_182
timestamp 1688980957
transform 1 0 17848 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_199
timestamp 1688980957
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_203
timestamp 1688980957
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_207
timestamp 1688980957
transform 1 0 20148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_211
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_215
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_238
timestamp 1688980957
transform 1 0 23000 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_242
timestamp 1688980957
transform 1 0 23368 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_246
timestamp 1688980957
transform 1 0 23736 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_250
timestamp 1688980957
transform 1 0 24104 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_254
timestamp 1688980957
transform 1 0 24472 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_258
timestamp 1688980957
transform 1 0 24840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_262
timestamp 1688980957
transform 1 0 25208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_266
timestamp 1688980957
transform 1 0 25576 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_297
timestamp 1688980957
transform 1 0 28428 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_326
timestamp 1688980957
transform 1 0 31096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_330
timestamp 1688980957
transform 1 0 31464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_341
timestamp 1688980957
transform 1 0 32476 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1688980957
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_32
timestamp 1688980957
transform 1 0 4048 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_36
timestamp 1688980957
transform 1 0 4416 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_48
timestamp 1688980957
transform 1 0 5520 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_59
timestamp 1688980957
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_63
timestamp 1688980957
transform 1 0 6900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_75
timestamp 1688980957
transform 1 0 8004 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_79
timestamp 1688980957
transform 1 0 8372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_114
timestamp 1688980957
transform 1 0 11592 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_147
timestamp 1688980957
transform 1 0 14628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_163
timestamp 1688980957
transform 1 0 16100 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_179
timestamp 1688980957
transform 1 0 17572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_183
timestamp 1688980957
transform 1 0 17940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_204
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_227
timestamp 1688980957
transform 1 0 21988 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_231
timestamp 1688980957
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_257
timestamp 1688980957
transform 1 0 24748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_264
timestamp 1688980957
transform 1 0 25392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_275
timestamp 1688980957
transform 1 0 26404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_288
timestamp 1688980957
transform 1 0 27600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_300
timestamp 1688980957
transform 1 0 28704 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_329
timestamp 1688980957
transform 1 0 31372 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_341
timestamp 1688980957
transform 1 0 32476 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_6
timestamp 1688980957
transform 1 0 1656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_12
timestamp 1688980957
transform 1 0 2208 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_16
timestamp 1688980957
transform 1 0 2576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_20
timestamp 1688980957
transform 1 0 2944 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_28
timestamp 1688980957
transform 1 0 3680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_62
timestamp 1688980957
transform 1 0 6808 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_85
timestamp 1688980957
transform 1 0 8924 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_92
timestamp 1688980957
transform 1 0 9568 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_96
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_106
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_132
timestamp 1688980957
transform 1 0 13248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_154
timestamp 1688980957
transform 1 0 15272 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_160
timestamp 1688980957
transform 1 0 15824 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_174
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_178
timestamp 1688980957
transform 1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_201
timestamp 1688980957
transform 1 0 19596 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_209
timestamp 1688980957
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_213
timestamp 1688980957
transform 1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_232
timestamp 1688980957
transform 1 0 22448 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_236
timestamp 1688980957
transform 1 0 22816 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_245
timestamp 1688980957
transform 1 0 23644 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_277
timestamp 1688980957
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_300
timestamp 1688980957
transform 1 0 28704 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_308
timestamp 1688980957
transform 1 0 29440 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_311
timestamp 1688980957
transform 1 0 29716 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_324
timestamp 1688980957
transform 1 0 30912 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_330
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_344
timestamp 1688980957
transform 1 0 32752 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_356
timestamp 1688980957
transform 1 0 33856 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_362
timestamp 1688980957
transform 1 0 34408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_365
timestamp 1688980957
transform 1 0 34684 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_23
timestamp 1688980957
transform 1 0 3220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_57
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_69
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_81
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_114
timestamp 1688980957
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_127
timestamp 1688980957
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_131
timestamp 1688980957
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_145
timestamp 1688980957
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_152
timestamp 1688980957
transform 1 0 15088 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_160
timestamp 1688980957
transform 1 0 15824 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_175
timestamp 1688980957
transform 1 0 17204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_180
timestamp 1688980957
transform 1 0 17664 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_184
timestamp 1688980957
transform 1 0 18032 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 1688980957
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_205
timestamp 1688980957
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_213
timestamp 1688980957
transform 1 0 20700 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_217
timestamp 1688980957
transform 1 0 21068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_231
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_235
timestamp 1688980957
transform 1 0 22724 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_239
timestamp 1688980957
transform 1 0 23092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_243
timestamp 1688980957
transform 1 0 23460 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_247
timestamp 1688980957
transform 1 0 23828 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_283
timestamp 1688980957
transform 1 0 27140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_291
timestamp 1688980957
transform 1 0 27876 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_299
timestamp 1688980957
transform 1 0 28612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_331
timestamp 1688980957
transform 1 0 31556 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_337
timestamp 1688980957
transform 1 0 32108 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_341
timestamp 1688980957
transform 1 0 32476 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_353
timestamp 1688980957
transform 1 0 33580 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_361
timestamp 1688980957
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_11
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_19
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_80
timestamp 1688980957
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_84
timestamp 1688980957
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_88
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_106
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1688980957
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_126
timestamp 1688980957
transform 1 0 12696 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_134
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_146
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_151
timestamp 1688980957
transform 1 0 14996 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_174
timestamp 1688980957
transform 1 0 17112 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_178
timestamp 1688980957
transform 1 0 17480 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_185
timestamp 1688980957
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_189
timestamp 1688980957
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_220
timestamp 1688980957
transform 1 0 21344 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_233
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_241
timestamp 1688980957
transform 1 0 23276 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_245
timestamp 1688980957
transform 1 0 23644 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_251
timestamp 1688980957
transform 1 0 24196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_259
timestamp 1688980957
transform 1 0 24932 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_268
timestamp 1688980957
transform 1 0 25760 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_301
timestamp 1688980957
transform 1 0 28796 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_313
timestamp 1688980957
transform 1 0 29900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_325
timestamp 1688980957
transform 1 0 31004 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_344
timestamp 1688980957
transform 1 0 32752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_7
timestamp 1688980957
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_32
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_36
timestamp 1688980957
transform 1 0 4416 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_40
timestamp 1688980957
transform 1 0 4784 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_52
timestamp 1688980957
transform 1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_75
timestamp 1688980957
transform 1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_79
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_96
timestamp 1688980957
transform 1 0 9936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_100
timestamp 1688980957
transform 1 0 10304 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_103
timestamp 1688980957
transform 1 0 10580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_149
timestamp 1688980957
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_159
timestamp 1688980957
transform 1 0 15732 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_166
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_173
timestamp 1688980957
transform 1 0 17020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_178
timestamp 1688980957
transform 1 0 17480 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_190
timestamp 1688980957
transform 1 0 18584 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_204
timestamp 1688980957
transform 1 0 19872 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_218
timestamp 1688980957
transform 1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_257
timestamp 1688980957
transform 1 0 24748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_288
timestamp 1688980957
transform 1 0 27600 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_300
timestamp 1688980957
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_326
timestamp 1688980957
transform 1 0 31096 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_338
timestamp 1688980957
transform 1 0 32200 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_346
timestamp 1688980957
transform 1 0 32936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_23
timestamp 1688980957
transform 1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_30
timestamp 1688980957
transform 1 0 3864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_34
timestamp 1688980957
transform 1 0 4232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_45
timestamp 1688980957
transform 1 0 5244 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_63
timestamp 1688980957
transform 1 0 6900 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_84
timestamp 1688980957
transform 1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_98
timestamp 1688980957
transform 1 0 10120 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_106
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_118
timestamp 1688980957
transform 1 0 11960 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_122
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_135
timestamp 1688980957
transform 1 0 13524 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_147
timestamp 1688980957
transform 1 0 14628 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_156
timestamp 1688980957
transform 1 0 15456 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_162
timestamp 1688980957
transform 1 0 16008 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_200
timestamp 1688980957
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_204
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_208
timestamp 1688980957
transform 1 0 20240 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_212
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_216
timestamp 1688980957
transform 1 0 20976 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_220
timestamp 1688980957
transform 1 0 21344 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_229
timestamp 1688980957
transform 1 0 22172 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_239
timestamp 1688980957
transform 1 0 23092 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_243
timestamp 1688980957
transform 1 0 23460 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_247
timestamp 1688980957
transform 1 0 23828 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_259
timestamp 1688980957
transform 1 0 24932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_278
timestamp 1688980957
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_287
timestamp 1688980957
transform 1 0 27508 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_301
timestamp 1688980957
transform 1 0 28796 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_309
timestamp 1688980957
transform 1 0 29532 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_334
timestamp 1688980957
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_367
timestamp 1688980957
transform 1 0 34868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_6
timestamp 1688980957
transform 1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_32
timestamp 1688980957
transform 1 0 4048 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_43
timestamp 1688980957
transform 1 0 5060 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_55
timestamp 1688980957
transform 1 0 6164 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_70
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_74
timestamp 1688980957
transform 1 0 7912 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_79
timestamp 1688980957
transform 1 0 8372 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_103
timestamp 1688980957
transform 1 0 10580 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_112
timestamp 1688980957
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_116
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_120
timestamp 1688980957
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_124
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_132
timestamp 1688980957
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_136
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_193
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_204
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_225
timestamp 1688980957
transform 1 0 21804 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_229
timestamp 1688980957
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_232
timestamp 1688980957
transform 1 0 22448 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_237
timestamp 1688980957
transform 1 0 22908 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_241
timestamp 1688980957
transform 1 0 23276 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_249
timestamp 1688980957
transform 1 0 24012 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_266
timestamp 1688980957
transform 1 0 25576 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_273
timestamp 1688980957
transform 1 0 26220 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_306
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_323
timestamp 1688980957
transform 1 0 30820 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_335
timestamp 1688980957
transform 1 0 31924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_347
timestamp 1688980957
transform 1 0 33028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_353
timestamp 1688980957
transform 1 0 33580 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_359
timestamp 1688980957
transform 1 0 34132 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_25
timestamp 1688980957
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_29
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_37
timestamp 1688980957
transform 1 0 4508 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_49
timestamp 1688980957
transform 1 0 5612 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_60
timestamp 1688980957
transform 1 0 6624 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_72
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_84
timestamp 1688980957
transform 1 0 8832 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_92
timestamp 1688980957
transform 1 0 9568 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_97
timestamp 1688980957
transform 1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_101
timestamp 1688980957
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_127
timestamp 1688980957
transform 1 0 12788 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_131
timestamp 1688980957
transform 1 0 13156 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_134
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_144
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_148
timestamp 1688980957
transform 1 0 14720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_156
timestamp 1688980957
transform 1 0 15456 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_160
timestamp 1688980957
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_164
timestamp 1688980957
transform 1 0 16192 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_184
timestamp 1688980957
transform 1 0 18032 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_191
timestamp 1688980957
transform 1 0 18676 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_200
timestamp 1688980957
transform 1 0 19504 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_204
timestamp 1688980957
transform 1 0 19872 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_208
timestamp 1688980957
transform 1 0 20240 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_220
timestamp 1688980957
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_240
timestamp 1688980957
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_244
timestamp 1688980957
transform 1 0 23552 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_248
timestamp 1688980957
transform 1 0 23920 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_256
timestamp 1688980957
transform 1 0 24656 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_263
timestamp 1688980957
transform 1 0 25300 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_275
timestamp 1688980957
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_291
timestamp 1688980957
transform 1 0 27876 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_297
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_309
timestamp 1688980957
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_321
timestamp 1688980957
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 1688980957
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_343
timestamp 1688980957
transform 1 0 32660 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_366
timestamp 1688980957
transform 1 0 34776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_45
timestamp 1688980957
transform 1 0 5244 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_75
timestamp 1688980957
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_96
timestamp 1688980957
transform 1 0 9936 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_104
timestamp 1688980957
transform 1 0 10672 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_113
timestamp 1688980957
transform 1 0 11500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_116
timestamp 1688980957
transform 1 0 11776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_120
timestamp 1688980957
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_124
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_128
timestamp 1688980957
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_154
timestamp 1688980957
transform 1 0 15272 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_158
timestamp 1688980957
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_168
timestamp 1688980957
transform 1 0 16560 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_185
timestamp 1688980957
transform 1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_205
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_212
timestamp 1688980957
transform 1 0 20608 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_217
timestamp 1688980957
transform 1 0 21068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_229
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_234
timestamp 1688980957
transform 1 0 22632 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_242
timestamp 1688980957
transform 1 0 23368 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_246
timestamp 1688980957
transform 1 0 23736 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_257
timestamp 1688980957
transform 1 0 24748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_266
timestamp 1688980957
transform 1 0 25576 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_274
timestamp 1688980957
transform 1 0 26312 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_286
timestamp 1688980957
transform 1 0 27416 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_298
timestamp 1688980957
transform 1 0 28520 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_320
timestamp 1688980957
transform 1 0 30544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_324
timestamp 1688980957
transform 1 0 30912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_332
timestamp 1688980957
transform 1 0 31648 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_343
timestamp 1688980957
transform 1 0 32660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_347
timestamp 1688980957
transform 1 0 33028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_23
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_35
timestamp 1688980957
transform 1 0 4324 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_47
timestamp 1688980957
transform 1 0 5428 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_101
timestamp 1688980957
transform 1 0 10396 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_107
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_122
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_157
timestamp 1688980957
transform 1 0 15548 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_194
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_206
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_215
timestamp 1688980957
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_222
timestamp 1688980957
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_244
timestamp 1688980957
transform 1 0 23552 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_252
timestamp 1688980957
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_274
timestamp 1688980957
transform 1 0 26312 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_291
timestamp 1688980957
transform 1 0 27876 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_302
timestamp 1688980957
transform 1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_327
timestamp 1688980957
transform 1 0 31188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_6
timestamp 1688980957
transform 1 0 1656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_18
timestamp 1688980957
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1688980957
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_36
timestamp 1688980957
transform 1 0 4416 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_51
timestamp 1688980957
transform 1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_59
timestamp 1688980957
transform 1 0 6532 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_63
timestamp 1688980957
transform 1 0 6900 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_75
timestamp 1688980957
transform 1 0 8004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_91
timestamp 1688980957
transform 1 0 9476 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_101
timestamp 1688980957
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_105
timestamp 1688980957
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_115
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_120
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_145
timestamp 1688980957
transform 1 0 14444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_149
timestamp 1688980957
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_180
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_192
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_230
timestamp 1688980957
transform 1 0 22264 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_247
timestamp 1688980957
transform 1 0 23828 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_266
timestamp 1688980957
transform 1 0 25576 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_278
timestamp 1688980957
transform 1 0 26680 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_284
timestamp 1688980957
transform 1 0 27232 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_302
timestamp 1688980957
transform 1 0 28888 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_351
timestamp 1688980957
transform 1 0 33396 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_26
timestamp 1688980957
transform 1 0 3496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_30
timestamp 1688980957
transform 1 0 3864 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_34
timestamp 1688980957
transform 1 0 4232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_46
timestamp 1688980957
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1688980957
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_87
timestamp 1688980957
transform 1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_91
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_100
timestamp 1688980957
transform 1 0 10304 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_132
timestamp 1688980957
transform 1 0 13248 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_173
timestamp 1688980957
transform 1 0 17020 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_185
timestamp 1688980957
transform 1 0 18124 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_189
timestamp 1688980957
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_204
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_216
timestamp 1688980957
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_231
timestamp 1688980957
transform 1 0 22356 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_238
timestamp 1688980957
transform 1 0 23000 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_242
timestamp 1688980957
transform 1 0 23368 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_254
timestamp 1688980957
transform 1 0 24472 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_266
timestamp 1688980957
transform 1 0 25576 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_278
timestamp 1688980957
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_313
timestamp 1688980957
transform 1 0 29900 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_319
timestamp 1688980957
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_331
timestamp 1688980957
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_341
timestamp 1688980957
transform 1 0 32476 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_364
timestamp 1688980957
transform 1 0 34592 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_115
timestamp 1688980957
transform 1 0 11684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_125
timestamp 1688980957
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_129
timestamp 1688980957
transform 1 0 12972 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_132
timestamp 1688980957
transform 1 0 13248 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_136
timestamp 1688980957
transform 1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_145
timestamp 1688980957
transform 1 0 14444 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_151
timestamp 1688980957
transform 1 0 14996 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_169
timestamp 1688980957
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_172
timestamp 1688980957
transform 1 0 16928 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_176
timestamp 1688980957
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_180
timestamp 1688980957
transform 1 0 17664 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_210
timestamp 1688980957
transform 1 0 20424 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_222
timestamp 1688980957
transform 1 0 21528 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_226
timestamp 1688980957
transform 1 0 21896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_229
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_247
timestamp 1688980957
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_271
timestamp 1688980957
transform 1 0 26036 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_303
timestamp 1688980957
transform 1 0 28980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_339
timestamp 1688980957
transform 1 0 32292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_347
timestamp 1688980957
transform 1 0 33028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_89
timestamp 1688980957
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_100
timestamp 1688980957
transform 1 0 10304 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_104
timestamp 1688980957
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_108
timestamp 1688980957
transform 1 0 11040 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_129
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_133
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_140
timestamp 1688980957
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_144
timestamp 1688980957
transform 1 0 14352 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_164
timestamp 1688980957
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_186
timestamp 1688980957
transform 1 0 18216 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_198
timestamp 1688980957
transform 1 0 19320 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_238
timestamp 1688980957
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_242
timestamp 1688980957
transform 1 0 23368 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_254
timestamp 1688980957
transform 1 0 24472 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_262
timestamp 1688980957
transform 1 0 25208 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_267
timestamp 1688980957
transform 1 0 25668 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_323
timestamp 1688980957
transform 1 0 30820 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_330
timestamp 1688980957
transform 1 0 31464 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_367
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_6
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_18
timestamp 1688980957
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_70
timestamp 1688980957
transform 1 0 7544 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_74
timestamp 1688980957
transform 1 0 7912 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 1688980957
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_113
timestamp 1688980957
transform 1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_120
timestamp 1688980957
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_124
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_127
timestamp 1688980957
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_145
timestamp 1688980957
transform 1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_151
timestamp 1688980957
transform 1 0 14996 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_157
timestamp 1688980957
transform 1 0 15548 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_163
timestamp 1688980957
transform 1 0 16100 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_166
timestamp 1688980957
transform 1 0 16376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_175
timestamp 1688980957
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_179
timestamp 1688980957
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_191
timestamp 1688980957
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_220
timestamp 1688980957
transform 1 0 21344 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_225
timestamp 1688980957
transform 1 0 21804 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_229
timestamp 1688980957
transform 1 0 22172 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_274
timestamp 1688980957
transform 1 0 26312 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_290
timestamp 1688980957
transform 1 0 27784 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_302
timestamp 1688980957
transform 1 0 28888 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_312
timestamp 1688980957
transform 1 0 29808 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_316
timestamp 1688980957
transform 1 0 30176 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_324
timestamp 1688980957
transform 1 0 30912 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_337
timestamp 1688980957
transform 1 0 32108 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_352
timestamp 1688980957
transform 1 0 33488 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_77
timestamp 1688980957
transform 1 0 8188 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_90
timestamp 1688980957
transform 1 0 9384 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_101
timestamp 1688980957
transform 1 0 10396 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1688980957
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_116
timestamp 1688980957
transform 1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_121
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_144
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_148
timestamp 1688980957
transform 1 0 14720 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_180
timestamp 1688980957
transform 1 0 17664 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_189
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_204
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_208
timestamp 1688980957
transform 1 0 20240 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_231
timestamp 1688980957
transform 1 0 22356 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_235
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_240
timestamp 1688980957
transform 1 0 23184 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_244
timestamp 1688980957
transform 1 0 23552 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_252
timestamp 1688980957
transform 1 0 24288 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_263
timestamp 1688980957
transform 1 0 25300 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_333
timestamp 1688980957
transform 1 0 31740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_358
timestamp 1688980957
transform 1 0 34040 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_366
timestamp 1688980957
transform 1 0 34776 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_26
timestamp 1688980957
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_33
timestamp 1688980957
transform 1 0 4140 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_36
timestamp 1688980957
transform 1 0 4416 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_52
timestamp 1688980957
transform 1 0 5888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_56
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_64
timestamp 1688980957
transform 1 0 6992 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_70
timestamp 1688980957
transform 1 0 7544 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_74
timestamp 1688980957
transform 1 0 7912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_80
timestamp 1688980957
transform 1 0 8464 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_89
timestamp 1688980957
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_122
timestamp 1688980957
transform 1 0 12328 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_134
timestamp 1688980957
transform 1 0 13432 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_159
timestamp 1688980957
transform 1 0 15732 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_163
timestamp 1688980957
transform 1 0 16100 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_178
timestamp 1688980957
transform 1 0 17480 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_183
timestamp 1688980957
transform 1 0 17940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_241
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_276
timestamp 1688980957
transform 1 0 26496 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_288
timestamp 1688980957
transform 1 0 27600 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_300
timestamp 1688980957
transform 1 0 28704 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_11
timestamp 1688980957
transform 1 0 2116 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_33
timestamp 1688980957
transform 1 0 4140 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_77
timestamp 1688980957
transform 1 0 8188 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_90
timestamp 1688980957
transform 1 0 9384 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_99
timestamp 1688980957
transform 1 0 10212 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_104
timestamp 1688980957
transform 1 0 10672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_108
timestamp 1688980957
transform 1 0 11040 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_119
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_143
timestamp 1688980957
transform 1 0 14260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_147
timestamp 1688980957
transform 1 0 14628 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_151
timestamp 1688980957
transform 1 0 14996 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_154
timestamp 1688980957
transform 1 0 15272 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_158
timestamp 1688980957
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1688980957
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_179
timestamp 1688980957
transform 1 0 17572 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_192
timestamp 1688980957
transform 1 0 18768 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_204
timestamp 1688980957
transform 1 0 19872 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_216
timestamp 1688980957
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_238
timestamp 1688980957
transform 1 0 23000 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_245
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_257
timestamp 1688980957
transform 1 0 24748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_269
timestamp 1688980957
transform 1 0 25852 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_321
timestamp 1688980957
transform 1 0 30636 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_325
timestamp 1688980957
transform 1 0 31004 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_341
timestamp 1688980957
transform 1 0 32476 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_352
timestamp 1688980957
transform 1 0 33488 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_364
timestamp 1688980957
transform 1 0 34592 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_6
timestamp 1688980957
transform 1 0 1656 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_14
timestamp 1688980957
transform 1 0 2392 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_22
timestamp 1688980957
transform 1 0 3128 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_35
timestamp 1688980957
transform 1 0 4324 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_43
timestamp 1688980957
transform 1 0 5060 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_55
timestamp 1688980957
transform 1 0 6164 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_67
timestamp 1688980957
transform 1 0 7268 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_75
timestamp 1688980957
transform 1 0 8004 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_79
timestamp 1688980957
transform 1 0 8372 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_91
timestamp 1688980957
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_94
timestamp 1688980957
transform 1 0 9752 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_106
timestamp 1688980957
transform 1 0 10856 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_114
timestamp 1688980957
transform 1 0 11592 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_118
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_132
timestamp 1688980957
transform 1 0 13248 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_136
timestamp 1688980957
transform 1 0 13616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_148
timestamp 1688980957
transform 1 0 14720 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_160
timestamp 1688980957
transform 1 0 15824 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_191
timestamp 1688980957
transform 1 0 18676 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_210
timestamp 1688980957
transform 1 0 20424 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_222
timestamp 1688980957
transform 1 0 21528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_248
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_258
timestamp 1688980957
transform 1 0 24840 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_270
timestamp 1688980957
transform 1 0 25944 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_282
timestamp 1688980957
transform 1 0 27048 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_294
timestamp 1688980957
transform 1 0 28152 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_337
timestamp 1688980957
transform 1 0 32108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_359
timestamp 1688980957
transform 1 0 34132 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_7
timestamp 1688980957
transform 1 0 1748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_28
timestamp 1688980957
transform 1 0 3680 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_36
timestamp 1688980957
transform 1 0 4416 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_40
timestamp 1688980957
transform 1 0 4784 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_47
timestamp 1688980957
transform 1 0 5428 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_80
timestamp 1688980957
transform 1 0 8464 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_92
timestamp 1688980957
transform 1 0 9568 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_98
timestamp 1688980957
transform 1 0 10120 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_102
timestamp 1688980957
transform 1 0 10488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_107
timestamp 1688980957
transform 1 0 10948 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_117
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_127
timestamp 1688980957
transform 1 0 12788 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_139
timestamp 1688980957
transform 1 0 13892 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_147
timestamp 1688980957
transform 1 0 14628 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_152
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_175
timestamp 1688980957
transform 1 0 17204 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_190
timestamp 1688980957
transform 1 0 18584 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_202
timestamp 1688980957
transform 1 0 19688 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_214
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_222
timestamp 1688980957
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_236
timestamp 1688980957
transform 1 0 22816 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_244
timestamp 1688980957
transform 1 0 23552 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_256
timestamp 1688980957
transform 1 0 24656 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_268
timestamp 1688980957
transform 1 0 25760 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_367
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_11
timestamp 1688980957
transform 1 0 2116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_19
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_25
timestamp 1688980957
transform 1 0 3404 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_38
timestamp 1688980957
transform 1 0 4600 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_56
timestamp 1688980957
transform 1 0 6256 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_60
timestamp 1688980957
transform 1 0 6624 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_105
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_123
timestamp 1688980957
transform 1 0 12420 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_127
timestamp 1688980957
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_131
timestamp 1688980957
transform 1 0 13156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_136
timestamp 1688980957
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_150
timestamp 1688980957
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_156
timestamp 1688980957
transform 1 0 15456 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_160
timestamp 1688980957
transform 1 0 15824 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_172
timestamp 1688980957
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_178
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_184
timestamp 1688980957
transform 1 0 18032 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_203
timestamp 1688980957
transform 1 0 19780 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_222
timestamp 1688980957
transform 1 0 21528 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_230
timestamp 1688980957
transform 1 0 22264 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_238
timestamp 1688980957
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_282
timestamp 1688980957
transform 1 0 27048 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_290
timestamp 1688980957
transform 1 0 27784 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_302
timestamp 1688980957
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_23
timestamp 1688980957
transform 1 0 3220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_31
timestamp 1688980957
transform 1 0 3956 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_34
timestamp 1688980957
transform 1 0 4232 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_60
timestamp 1688980957
transform 1 0 6624 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_72
timestamp 1688980957
transform 1 0 7728 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_82
timestamp 1688980957
transform 1 0 8648 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_92
timestamp 1688980957
transform 1 0 9568 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_96
timestamp 1688980957
transform 1 0 9936 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_119
timestamp 1688980957
transform 1 0 12052 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_159
timestamp 1688980957
transform 1 0 15732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_163
timestamp 1688980957
transform 1 0 16100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_174
timestamp 1688980957
transform 1 0 17112 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_178
timestamp 1688980957
transform 1 0 17480 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_182
timestamp 1688980957
transform 1 0 17848 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_212
timestamp 1688980957
transform 1 0 20608 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_230
timestamp 1688980957
transform 1 0 22264 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_248
timestamp 1688980957
transform 1 0 23920 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_260
timestamp 1688980957
transform 1 0 25024 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_268
timestamp 1688980957
transform 1 0 25760 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_272
timestamp 1688980957
transform 1 0 26128 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_288
timestamp 1688980957
transform 1 0 27600 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_313
timestamp 1688980957
transform 1 0 29900 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_367
timestamp 1688980957
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_32
timestamp 1688980957
transform 1 0 4048 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_40
timestamp 1688980957
transform 1 0 4784 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_51
timestamp 1688980957
transform 1 0 5796 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_63
timestamp 1688980957
transform 1 0 6900 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_75
timestamp 1688980957
transform 1 0 8004 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_88
timestamp 1688980957
transform 1 0 9200 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_99
timestamp 1688980957
transform 1 0 10212 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_114
timestamp 1688980957
transform 1 0 11592 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_120
timestamp 1688980957
transform 1 0 12144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_125
timestamp 1688980957
transform 1 0 12604 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_129
timestamp 1688980957
transform 1 0 12972 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_158
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_181
timestamp 1688980957
transform 1 0 17756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_192
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_202
timestamp 1688980957
transform 1 0 19688 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_206
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_217
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_229
timestamp 1688980957
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_241
timestamp 1688980957
transform 1 0 23276 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_249
timestamp 1688980957
transform 1 0 24012 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_290
timestamp 1688980957
transform 1 0 27784 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_302
timestamp 1688980957
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_332
timestamp 1688980957
transform 1 0 31648 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_336
timestamp 1688980957
transform 1 0 32016 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_348
timestamp 1688980957
transform 1 0 33120 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_354
timestamp 1688980957
transform 1 0 33672 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_362
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_6
timestamp 1688980957
transform 1 0 1656 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_18
timestamp 1688980957
transform 1 0 2760 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_26
timestamp 1688980957
transform 1 0 3496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_45
timestamp 1688980957
transform 1 0 5244 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_116
timestamp 1688980957
transform 1 0 11776 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_126
timestamp 1688980957
transform 1 0 12696 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_130
timestamp 1688980957
transform 1 0 13064 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_135
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_139
timestamp 1688980957
transform 1 0 13892 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_143
timestamp 1688980957
transform 1 0 14260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_160
timestamp 1688980957
transform 1 0 15824 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_164
timestamp 1688980957
transform 1 0 16192 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_176
timestamp 1688980957
transform 1 0 17296 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_180
timestamp 1688980957
transform 1 0 17664 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_196
timestamp 1688980957
transform 1 0 19136 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_200
timestamp 1688980957
transform 1 0 19504 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_212
timestamp 1688980957
transform 1 0 20608 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_258
timestamp 1688980957
transform 1 0 24840 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_264
timestamp 1688980957
transform 1 0 25392 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_276
timestamp 1688980957
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_301
timestamp 1688980957
transform 1 0 28796 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_328
timestamp 1688980957
transform 1 0 31280 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_332
timestamp 1688980957
transform 1 0 31648 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_360
timestamp 1688980957
transform 1 0 34224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_364
timestamp 1688980957
transform 1 0 34592 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_9
timestamp 1688980957
transform 1 0 1932 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_12
timestamp 1688980957
transform 1 0 2208 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_24
timestamp 1688980957
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_33
timestamp 1688980957
transform 1 0 4140 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_50
timestamp 1688980957
transform 1 0 5704 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_62
timestamp 1688980957
transform 1 0 6808 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_74
timestamp 1688980957
transform 1 0 7912 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_78
timestamp 1688980957
transform 1 0 8280 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 1688980957
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_101
timestamp 1688980957
transform 1 0 10396 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_131
timestamp 1688980957
transform 1 0 13156 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_146
timestamp 1688980957
transform 1 0 14536 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_150
timestamp 1688980957
transform 1 0 14904 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_154
timestamp 1688980957
transform 1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_158
timestamp 1688980957
transform 1 0 15640 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_162
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_169
timestamp 1688980957
transform 1 0 16652 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_179
timestamp 1688980957
transform 1 0 17572 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_191
timestamp 1688980957
transform 1 0 18676 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_216
timestamp 1688980957
transform 1 0 20976 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_238
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_244
timestamp 1688980957
transform 1 0 23552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_260
timestamp 1688980957
transform 1 0 25024 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_269
timestamp 1688980957
transform 1 0 25852 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_273
timestamp 1688980957
transform 1 0 26220 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_296
timestamp 1688980957
transform 1 0 28336 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_328
timestamp 1688980957
transform 1 0 31280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_334
timestamp 1688980957
transform 1 0 31832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_337
timestamp 1688980957
transform 1 0 32108 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_6
timestamp 1688980957
transform 1 0 1656 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_33
timestamp 1688980957
transform 1 0 4140 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_37
timestamp 1688980957
transform 1 0 4508 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_41
timestamp 1688980957
transform 1 0 4876 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_45
timestamp 1688980957
transform 1 0 5244 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_49
timestamp 1688980957
transform 1 0 5612 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_89
timestamp 1688980957
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_94
timestamp 1688980957
transform 1 0 9752 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_98
timestamp 1688980957
transform 1 0 10120 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_110
timestamp 1688980957
transform 1 0 11224 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_133
timestamp 1688980957
transform 1 0 13340 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_141
timestamp 1688980957
transform 1 0 14076 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_145
timestamp 1688980957
transform 1 0 14444 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_148
timestamp 1688980957
transform 1 0 14720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_153
timestamp 1688980957
transform 1 0 15180 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_175
timestamp 1688980957
transform 1 0 17204 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_187
timestamp 1688980957
transform 1 0 18308 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_199
timestamp 1688980957
transform 1 0 19412 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_222
timestamp 1688980957
transform 1 0 21528 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_231
timestamp 1688980957
transform 1 0 22356 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_243
timestamp 1688980957
transform 1 0 23460 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_255
timestamp 1688980957
transform 1 0 24564 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_267
timestamp 1688980957
transform 1 0 25668 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_314
timestamp 1688980957
transform 1 0 29992 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_318
timestamp 1688980957
transform 1 0 30360 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_322
timestamp 1688980957
transform 1 0 30728 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_333
timestamp 1688980957
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_363
timestamp 1688980957
transform 1 0 34500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_367
timestamp 1688980957
transform 1 0 34868 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_49
timestamp 1688980957
transform 1 0 5612 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_61
timestamp 1688980957
transform 1 0 6716 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_108
timestamp 1688980957
transform 1 0 11040 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_112
timestamp 1688980957
transform 1 0 11408 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_124
timestamp 1688980957
transform 1 0 12512 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_157
timestamp 1688980957
transform 1 0 15548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_169
timestamp 1688980957
transform 1 0 16652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_173
timestamp 1688980957
transform 1 0 17020 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_191
timestamp 1688980957
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_205
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_212
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_236
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_248
timestamp 1688980957
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_263
timestamp 1688980957
transform 1 0 25300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_275
timestamp 1688980957
transform 1 0 26404 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_279
timestamp 1688980957
transform 1 0 26772 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_302
timestamp 1688980957
transform 1 0 28888 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_317
timestamp 1688980957
transform 1 0 30268 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_324
timestamp 1688980957
transform 1 0 30912 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_330
timestamp 1688980957
transform 1 0 31464 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_23
timestamp 1688980957
transform 1 0 3220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_28
timestamp 1688980957
transform 1 0 3680 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_35
timestamp 1688980957
transform 1 0 4324 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_145
timestamp 1688980957
transform 1 0 14444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_166
timestamp 1688980957
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_195
timestamp 1688980957
transform 1 0 19044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_202
timestamp 1688980957
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_213
timestamp 1688980957
transform 1 0 20700 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_234
timestamp 1688980957
transform 1 0 22632 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_240
timestamp 1688980957
transform 1 0 23184 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_259
timestamp 1688980957
transform 1 0 24932 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_272
timestamp 1688980957
transform 1 0 26128 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_304
timestamp 1688980957
transform 1 0 29072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_308
timestamp 1688980957
transform 1 0 29440 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_312
timestamp 1688980957
transform 1 0 29808 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_320
timestamp 1688980957
transform 1 0 30544 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_331
timestamp 1688980957
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_345
timestamp 1688980957
transform 1 0 32844 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_49
timestamp 1688980957
transform 1 0 5612 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_159
timestamp 1688980957
transform 1 0 15732 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_171
timestamp 1688980957
transform 1 0 16836 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_180
timestamp 1688980957
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_184
timestamp 1688980957
transform 1 0 18032 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_187
timestamp 1688980957
transform 1 0 18308 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_191
timestamp 1688980957
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_201
timestamp 1688980957
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_208
timestamp 1688980957
transform 1 0 20240 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_220
timestamp 1688980957
transform 1 0 21344 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_232
timestamp 1688980957
transform 1 0 22448 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_240
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_246
timestamp 1688980957
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_279
timestamp 1688980957
transform 1 0 26772 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_286
timestamp 1688980957
transform 1 0 27416 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_298
timestamp 1688980957
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_306
timestamp 1688980957
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_327
timestamp 1688980957
transform 1 0 31188 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_352
timestamp 1688980957
transform 1 0 33488 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_356
timestamp 1688980957
transform 1 0 33856 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_361
timestamp 1688980957
transform 1 0 34316 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_218
timestamp 1688980957
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_238
timestamp 1688980957
transform 1 0 23000 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_250
timestamp 1688980957
transform 1 0 24104 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_262
timestamp 1688980957
transform 1 0 25208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_274
timestamp 1688980957
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_313
timestamp 1688980957
transform 1 0 29900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_316
timestamp 1688980957
transform 1 0 30176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_320
timestamp 1688980957
transform 1 0 30544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_326
timestamp 1688980957
transform 1 0 31096 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_330
timestamp 1688980957
transform 1 0 31464 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_334
timestamp 1688980957
transform 1 0 31832 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_363
timestamp 1688980957
transform 1 0 34500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_367
timestamp 1688980957
transform 1 0 34868 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_6
timestamp 1688980957
transform 1 0 1656 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_18
timestamp 1688980957
transform 1 0 2760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_207
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_215
timestamp 1688980957
transform 1 0 20884 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_223
timestamp 1688980957
transform 1 0 21620 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_235
timestamp 1688980957
transform 1 0 22724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_247
timestamp 1688980957
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_341
timestamp 1688980957
transform 1 0 32476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_367
timestamp 1688980957
transform 1 0 34868 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_367
timestamp 1688980957
transform 1 0 34868 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_6
timestamp 1688980957
transform 1 0 1656 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_18
timestamp 1688980957
transform 1 0 2760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_367
timestamp 1688980957
transform 1 0 34868 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_367
timestamp 1688980957
transform 1 0 34868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_6
timestamp 1688980957
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_18
timestamp 1688980957
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_26
timestamp 1688980957
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_367
timestamp 1688980957
transform 1 0 34868 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_367
timestamp 1688980957
transform 1 0 34868 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_6
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_18
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_367
timestamp 1688980957
transform 1 0 34868 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_6
timestamp 1688980957
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1688980957
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_69
timestamp 1688980957
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_81
timestamp 1688980957
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_113
timestamp 1688980957
transform 1 0 11500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_125
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_169
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_181
timestamp 1688980957
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_237
timestamp 1688980957
transform 1 0 22908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_249
timestamp 1688980957
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_281
timestamp 1688980957
transform 1 0 26956 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_293
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_305
timestamp 1688980957
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_337
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 1656 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 1656 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 1656 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input17 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 27324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap36
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output20
timestamp 1688980957
transform -1 0 34592 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 1688980957
transform -1 0 34592 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 1688980957
transform 1 0 33488 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 1688980957
transform -1 0 34592 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 1688980957
transform -1 0 34592 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 1688980957
transform -1 0 34592 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 1688980957
transform 1 0 33120 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 1688980957
transform -1 0 34592 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 1688980957
transform -1 0 34960 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 1688980957
transform -1 0 34960 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 1688980957
transform -1 0 34960 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 1688980957
transform -1 0 34592 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 1688980957
transform -1 0 34592 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 1688980957
transform -1 0 34592 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output35
timestamp 1688980957
transform -1 0 34592 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 35236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 35236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 35236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 35236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 35236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 35236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 35236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 35236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 35236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 35236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 35236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 35236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 35236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 35236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 35236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 35236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 35236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 35236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 35236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 35236 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 35236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 35236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 35236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 35236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 35236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 35236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 35236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 35236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 35236 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 35236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 35236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 35236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 35236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 35236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 35236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 35236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 35236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 35236 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 35236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 35236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 35236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 35236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 35236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 35236 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 35236 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 35236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 35236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 35236 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126 unic-cass/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 11408 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 21712 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 32016 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 a[0]
port 0 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 a[1]
port 1 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 a[2]
port 2 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 a[3]
port 3 nsew signal input
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 a[4]
port 4 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 a[5]
port 5 nsew signal input
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 a[6]
port 6 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 a[7]
port 7 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 b[0]
port 8 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 b[1]
port 9 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 b[2]
port 10 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 b[3]
port 11 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 b[4]
port 12 nsew signal input
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 b[5]
port 13 nsew signal input
flabel metal3 s 0 32376 800 32496 0 FreeSans 480 0 0 0 b[6]
port 14 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 b[7]
port 15 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 control
port 17 nsew signal input
flabel metal3 s 35600 3000 36400 3120 0 FreeSans 480 0 0 0 p[0]
port 18 nsew signal tristate
flabel metal3 s 35600 24760 36400 24880 0 FreeSans 480 0 0 0 p[10]
port 19 nsew signal tristate
flabel metal3 s 35600 26936 36400 27056 0 FreeSans 480 0 0 0 p[11]
port 20 nsew signal tristate
flabel metal3 s 35600 29112 36400 29232 0 FreeSans 480 0 0 0 p[12]
port 21 nsew signal tristate
flabel metal3 s 35600 31288 36400 31408 0 FreeSans 480 0 0 0 p[13]
port 22 nsew signal tristate
flabel metal3 s 35600 33464 36400 33584 0 FreeSans 480 0 0 0 p[14]
port 23 nsew signal tristate
flabel metal3 s 35600 35640 36400 35760 0 FreeSans 480 0 0 0 p[15]
port 24 nsew signal tristate
flabel metal3 s 35600 5176 36400 5296 0 FreeSans 480 0 0 0 p[1]
port 25 nsew signal tristate
flabel metal3 s 35600 7352 36400 7472 0 FreeSans 480 0 0 0 p[2]
port 26 nsew signal tristate
flabel metal3 s 35600 9528 36400 9648 0 FreeSans 480 0 0 0 p[3]
port 27 nsew signal tristate
flabel metal3 s 35600 11704 36400 11824 0 FreeSans 480 0 0 0 p[4]
port 28 nsew signal tristate
flabel metal3 s 35600 13880 36400 14000 0 FreeSans 480 0 0 0 p[5]
port 29 nsew signal tristate
flabel metal3 s 35600 16056 36400 16176 0 FreeSans 480 0 0 0 p[6]
port 30 nsew signal tristate
flabel metal3 s 35600 18232 36400 18352 0 FreeSans 480 0 0 0 p[7]
port 31 nsew signal tristate
flabel metal3 s 35600 20408 36400 20528 0 FreeSans 480 0 0 0 p[8]
port 32 nsew signal tristate
flabel metal3 s 35600 22584 36400 22704 0 FreeSans 480 0 0 0 p[9]
port 33 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 rst
port 34 nsew signal input
flabel metal4 s 4208 2128 4528 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 34928 2128 35248 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 19568 2128 19888 36496 0 FreeSans 1920 90 0 0 vssd1
port 36 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36400 38800
<< end >>
