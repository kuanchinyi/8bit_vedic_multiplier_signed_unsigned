magic
tech sky130A
magscale 1 2
timestamp 1729948588
<< viali >>
rect 1409 36125 1443 36159
rect 33333 36125 33367 36159
rect 34345 36057 34379 36091
rect 1593 35989 1627 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 34069 34017 34103 34051
rect 34529 33949 34563 33983
rect 1409 32861 1443 32895
rect 1593 32725 1627 32759
rect 34069 31841 34103 31875
rect 34529 31773 34563 31807
rect 1409 30685 1443 30719
rect 32873 30685 32907 30719
rect 32781 30617 32815 30651
rect 1593 30549 1627 30583
rect 32965 30549 32999 30583
rect 30941 30209 30975 30243
rect 32137 30209 32171 30243
rect 34345 30209 34379 30243
rect 28549 30141 28583 30175
rect 28825 30141 28859 30175
rect 30297 30141 30331 30175
rect 31033 30141 31067 30175
rect 32413 30141 32447 30175
rect 31309 30073 31343 30107
rect 33885 30073 33919 30107
rect 28457 30005 28491 30039
rect 31861 30005 31895 30039
rect 34253 30005 34287 30039
rect 34621 30005 34655 30039
rect 26525 29801 26559 29835
rect 29285 29801 29319 29835
rect 34529 29801 34563 29835
rect 25421 29733 25455 29767
rect 25145 29665 25179 29699
rect 27813 29665 27847 29699
rect 29561 29665 29595 29699
rect 31309 29665 31343 29699
rect 32229 29665 32263 29699
rect 24041 29597 24075 29631
rect 24225 29597 24259 29631
rect 25053 29597 25087 29631
rect 26157 29597 26191 29631
rect 26249 29597 26283 29631
rect 26341 29597 26375 29631
rect 27905 29597 27939 29631
rect 29193 29597 29227 29631
rect 32137 29597 32171 29631
rect 32781 29597 32815 29631
rect 29837 29529 29871 29563
rect 33057 29529 33091 29563
rect 24225 29461 24259 29495
rect 28273 29461 28307 29495
rect 29101 29461 29135 29495
rect 32505 29461 32539 29495
rect 23305 29257 23339 29291
rect 25145 29257 25179 29291
rect 29469 29257 29503 29291
rect 30389 29257 30423 29291
rect 32597 29257 32631 29291
rect 32965 29257 32999 29291
rect 34897 29257 34931 29291
rect 23949 29189 23983 29223
rect 23213 29121 23247 29155
rect 23489 29121 23523 29155
rect 23581 29121 23615 29155
rect 23765 29121 23799 29155
rect 24225 29121 24259 29155
rect 24409 29121 24443 29155
rect 24685 29121 24719 29155
rect 24869 29121 24903 29155
rect 24961 29121 24995 29155
rect 25145 29121 25179 29155
rect 25513 29121 25547 29155
rect 25697 29121 25731 29155
rect 30297 29121 30331 29155
rect 33149 29121 33183 29155
rect 24593 29053 24627 29087
rect 24869 28985 24903 29019
rect 25605 28985 25639 29019
rect 23489 28917 23523 28951
rect 30205 28917 30239 28951
rect 33406 28917 33440 28951
rect 24041 28713 24075 28747
rect 28365 28713 28399 28747
rect 31401 28713 31435 28747
rect 32505 28713 32539 28747
rect 34805 28713 34839 28747
rect 24777 28645 24811 28679
rect 25927 28645 25961 28679
rect 31677 28645 31711 28679
rect 32781 28645 32815 28679
rect 25329 28577 25363 28611
rect 25789 28577 25823 28611
rect 26893 28577 26927 28611
rect 26985 28577 27019 28611
rect 27629 28577 27663 28611
rect 29377 28577 29411 28611
rect 29561 28577 29595 28611
rect 31309 28577 31343 28611
rect 32321 28577 32355 28611
rect 34069 28577 34103 28611
rect 1409 28509 1443 28543
rect 23765 28509 23799 28543
rect 23857 28509 23891 28543
rect 24133 28509 24167 28543
rect 24409 28509 24443 28543
rect 24593 28509 24627 28543
rect 25513 28509 25547 28543
rect 25605 28509 25639 28543
rect 26065 28509 26099 28543
rect 27353 28509 27387 28543
rect 27721 28509 27755 28543
rect 27905 28509 27939 28543
rect 27997 28509 28031 28543
rect 28181 28509 28215 28543
rect 28273 28509 28307 28543
rect 28641 28509 28675 28543
rect 31585 28509 31619 28543
rect 31769 28509 31803 28543
rect 31861 28509 31895 28543
rect 32229 28509 32263 28543
rect 32689 28509 32723 28543
rect 32873 28509 32907 28543
rect 34529 28509 34563 28543
rect 34713 28509 34747 28543
rect 24501 28441 24535 28475
rect 24777 28441 24811 28475
rect 25697 28441 25731 28475
rect 27261 28441 27295 28475
rect 28365 28441 28399 28475
rect 28549 28441 28583 28475
rect 29837 28441 29871 28475
rect 1593 28373 1627 28407
rect 23581 28373 23615 28407
rect 25237 28373 25271 28407
rect 27169 28373 27203 28407
rect 27721 28169 27755 28203
rect 27905 28169 27939 28203
rect 30297 28169 30331 28203
rect 32413 28169 32447 28203
rect 27537 28033 27571 28067
rect 27721 28033 27755 28067
rect 27813 28033 27847 28067
rect 27997 28033 28031 28067
rect 30205 28033 30239 28067
rect 32137 28033 32171 28067
rect 32413 27965 32447 27999
rect 30113 27829 30147 27863
rect 32229 27829 32263 27863
rect 34253 27829 34287 27863
rect 34529 27829 34563 27863
rect 19809 27625 19843 27659
rect 24593 27625 24627 27659
rect 24777 27625 24811 27659
rect 26249 27625 26283 27659
rect 26341 27625 26375 27659
rect 31769 27625 31803 27659
rect 34529 27625 34563 27659
rect 22661 27557 22695 27591
rect 20269 27489 20303 27523
rect 22385 27489 22419 27523
rect 25237 27489 25271 27523
rect 28089 27489 28123 27523
rect 28365 27489 28399 27523
rect 28641 27489 28675 27523
rect 32137 27489 32171 27523
rect 32781 27489 32815 27523
rect 19257 27421 19291 27455
rect 19349 27421 19383 27455
rect 19533 27421 19567 27455
rect 19625 27421 19659 27455
rect 19993 27421 20027 27455
rect 20085 27421 20119 27455
rect 20177 27421 20211 27455
rect 22293 27421 22327 27455
rect 24869 27421 24903 27455
rect 25053 27421 25087 27455
rect 25697 27421 25731 27455
rect 25789 27421 25823 27455
rect 25973 27421 26007 27455
rect 26065 27421 26099 27455
rect 26617 27421 26651 27455
rect 27997 27421 28031 27455
rect 28733 27421 28767 27455
rect 31401 27421 31435 27455
rect 32045 27421 32079 27455
rect 34713 27421 34747 27455
rect 24409 27353 24443 27387
rect 26341 27353 26375 27387
rect 31585 27353 31619 27387
rect 33057 27353 33091 27387
rect 34805 27353 34839 27387
rect 20453 27285 20487 27319
rect 24609 27285 24643 27319
rect 26525 27285 26559 27319
rect 29101 27285 29135 27319
rect 32413 27285 32447 27319
rect 17601 27081 17635 27115
rect 19441 27081 19475 27115
rect 20177 27081 20211 27115
rect 20637 27081 20671 27115
rect 24501 27081 24535 27115
rect 25789 27081 25823 27115
rect 26709 27081 26743 27115
rect 27077 27081 27111 27115
rect 29561 27081 29595 27115
rect 31401 27081 31435 27115
rect 32229 27081 32263 27115
rect 32597 27081 32631 27115
rect 25513 27013 25547 27047
rect 29929 27013 29963 27047
rect 31585 27013 31619 27047
rect 13369 26945 13403 26979
rect 17417 26945 17451 26979
rect 17601 26945 17635 26979
rect 17693 26945 17727 26979
rect 17877 26945 17911 26979
rect 18797 26945 18831 26979
rect 18976 26945 19010 26979
rect 19073 26945 19107 26979
rect 19165 26945 19199 26979
rect 19533 26945 19567 26979
rect 19717 26945 19751 26979
rect 19809 26945 19843 26979
rect 19901 26945 19935 26979
rect 20545 26945 20579 26979
rect 21281 26945 21315 26979
rect 21373 26945 21407 26979
rect 23213 26945 23247 26979
rect 24409 26945 24443 26979
rect 24593 26945 24627 26979
rect 24685 26945 24719 26979
rect 24869 26945 24903 26979
rect 25329 26945 25363 26979
rect 25973 26945 26007 26979
rect 26065 26945 26099 26979
rect 26157 26945 26191 26979
rect 26341 26945 26375 26979
rect 26433 26945 26467 26979
rect 26525 26945 26559 26979
rect 26801 26945 26835 26979
rect 26985 26945 27019 26979
rect 27169 26945 27203 26979
rect 31493 26945 31527 26979
rect 32137 26945 32171 26979
rect 32321 26945 32355 26979
rect 34713 26945 34747 26979
rect 13185 26877 13219 26911
rect 22385 26877 22419 26911
rect 25697 26877 25731 26911
rect 29653 26877 29687 26911
rect 34437 26877 34471 26911
rect 17877 26809 17911 26843
rect 26525 26809 26559 26843
rect 13553 26741 13587 26775
rect 15393 26741 15427 26775
rect 16037 26741 16071 26775
rect 23489 26741 23523 26775
rect 23857 26741 23891 26775
rect 25053 26741 25087 26775
rect 13093 26537 13127 26571
rect 13369 26537 13403 26571
rect 15393 26537 15427 26571
rect 19993 26537 20027 26571
rect 22201 26537 22235 26571
rect 22477 26537 22511 26571
rect 23857 26537 23891 26571
rect 26249 26537 26283 26571
rect 32597 26537 32631 26571
rect 34529 26537 34563 26571
rect 15577 26469 15611 26503
rect 19073 26469 19107 26503
rect 19625 26469 19659 26503
rect 23213 26469 23247 26503
rect 15945 26401 15979 26435
rect 18245 26401 18279 26435
rect 19533 26401 19567 26435
rect 21097 26401 21131 26435
rect 22845 26401 22879 26435
rect 23397 26401 23431 26435
rect 32781 26401 32815 26435
rect 1409 26333 1443 26367
rect 13001 26333 13035 26367
rect 13277 26333 13311 26367
rect 13553 26333 13587 26367
rect 13645 26333 13679 26367
rect 13829 26333 13863 26367
rect 13921 26333 13955 26367
rect 14565 26333 14599 26367
rect 14749 26333 14783 26367
rect 15485 26333 15519 26367
rect 15761 26333 15795 26367
rect 16037 26333 16071 26367
rect 16221 26333 16255 26367
rect 16497 26333 16531 26367
rect 16681 26333 16715 26367
rect 17233 26333 17267 26367
rect 17417 26333 17451 26367
rect 18429 26333 18463 26367
rect 18613 26333 18647 26367
rect 18705 26333 18739 26367
rect 18797 26333 18831 26367
rect 19257 26333 19291 26367
rect 19441 26333 19475 26367
rect 19717 26333 19751 26367
rect 22109 26333 22143 26367
rect 22293 26333 22327 26367
rect 22385 26333 22419 26367
rect 22569 26333 22603 26367
rect 23029 26333 23063 26367
rect 23489 26333 23523 26367
rect 23581 26333 23615 26367
rect 23673 26333 23707 26367
rect 25717 26333 25751 26367
rect 25881 26333 25915 26367
rect 26065 26333 26099 26367
rect 34713 26333 34747 26367
rect 21465 26265 21499 26299
rect 24133 26265 24167 26299
rect 25973 26265 26007 26299
rect 33057 26265 33091 26299
rect 34805 26265 34839 26299
rect 1593 26197 1627 26231
rect 9505 26197 9539 26231
rect 12725 26197 12759 26231
rect 17049 26197 17083 26231
rect 20729 26197 20763 26231
rect 21741 26197 21775 26231
rect 31309 26197 31343 26231
rect 12725 25993 12759 26027
rect 16221 25993 16255 26027
rect 16681 25993 16715 26027
rect 18061 25993 18095 26027
rect 19441 25993 19475 26027
rect 21189 25993 21223 26027
rect 27261 25993 27295 26027
rect 29101 25993 29135 26027
rect 31585 25993 31619 26027
rect 32689 25993 32723 26027
rect 11253 25925 11287 25959
rect 12357 25925 12391 25959
rect 12449 25925 12483 25959
rect 12909 25925 12943 25959
rect 15669 25925 15703 25959
rect 15869 25925 15903 25959
rect 17509 25925 17543 25959
rect 19349 25925 19383 25959
rect 29469 25925 29503 25959
rect 29837 25925 29871 25959
rect 8677 25857 8711 25891
rect 10425 25857 10459 25891
rect 11069 25857 11103 25891
rect 11529 25857 11563 25891
rect 11621 25857 11655 25891
rect 11805 25857 11839 25891
rect 12239 25857 12273 25891
rect 12541 25857 12575 25891
rect 12817 25857 12851 25891
rect 13001 25857 13035 25891
rect 13461 25857 13495 25891
rect 13550 25863 13584 25897
rect 13645 25857 13679 25891
rect 13829 25857 13863 25891
rect 13921 25857 13955 25891
rect 14105 25857 14139 25891
rect 14841 25857 14875 25891
rect 15025 25857 15059 25891
rect 15577 25857 15611 25891
rect 16129 25857 16163 25891
rect 16313 25857 16347 25891
rect 16865 25857 16899 25891
rect 17049 25857 17083 25891
rect 17141 25857 17175 25891
rect 18061 25857 18095 25891
rect 18889 25857 18923 25891
rect 18981 25857 19015 25891
rect 19165 25857 19199 25891
rect 19625 25857 19659 25891
rect 21403 25857 21437 25891
rect 21557 25857 21591 25891
rect 27537 25857 27571 25891
rect 27813 25857 27847 25891
rect 28733 25857 28767 25891
rect 31953 25857 31987 25891
rect 32321 25857 32355 25891
rect 10885 25789 10919 25823
rect 11989 25789 12023 25823
rect 12081 25789 12115 25823
rect 15117 25789 15151 25823
rect 18153 25789 18187 25823
rect 18337 25789 18371 25823
rect 19257 25789 19291 25823
rect 19809 25789 19843 25823
rect 27261 25789 27295 25823
rect 27721 25789 27755 25823
rect 28181 25789 28215 25823
rect 28641 25789 28675 25823
rect 29561 25789 29595 25823
rect 31309 25789 31343 25823
rect 31861 25789 31895 25823
rect 32229 25789 32263 25823
rect 9413 25721 9447 25755
rect 14473 25721 14507 25755
rect 16957 25721 16991 25755
rect 23765 25721 23799 25755
rect 27445 25721 27479 25755
rect 8953 25653 8987 25687
rect 9689 25653 9723 25687
rect 10793 25653 10827 25687
rect 13185 25653 13219 25687
rect 14013 25653 14047 25687
rect 14933 25653 14967 25687
rect 15485 25653 15519 25687
rect 15853 25653 15887 25687
rect 16037 25653 16071 25687
rect 20545 25653 20579 25687
rect 21005 25653 21039 25687
rect 22385 25653 22419 25687
rect 22661 25653 22695 25687
rect 23029 25653 23063 25687
rect 23397 25653 23431 25687
rect 31953 25653 31987 25687
rect 34529 25653 34563 25687
rect 13645 25449 13679 25483
rect 14289 25449 14323 25483
rect 15025 25449 15059 25483
rect 16681 25449 16715 25483
rect 23029 25449 23063 25483
rect 23765 25449 23799 25483
rect 24869 25449 24903 25483
rect 30573 25449 30607 25483
rect 32045 25449 32079 25483
rect 8401 25381 8435 25415
rect 21097 25381 21131 25415
rect 9873 25313 9907 25347
rect 11345 25313 11379 25347
rect 15163 25313 15197 25347
rect 15577 25313 15611 25347
rect 16313 25313 16347 25347
rect 21833 25313 21867 25347
rect 22569 25313 22603 25347
rect 24961 25313 24995 25347
rect 27537 25313 27571 25347
rect 31953 25313 31987 25347
rect 32137 25313 32171 25347
rect 34069 25313 34103 25347
rect 9321 25245 9355 25279
rect 9505 25245 9539 25279
rect 10057 25245 10091 25279
rect 10241 25245 10275 25279
rect 10888 25223 10922 25257
rect 10977 25245 11011 25279
rect 11161 25245 11195 25279
rect 11253 25245 11287 25279
rect 11621 25245 11655 25279
rect 11713 25245 11747 25279
rect 11805 25245 11839 25279
rect 11989 25245 12023 25279
rect 12265 25245 12299 25279
rect 12357 25245 12391 25279
rect 12541 25245 12575 25279
rect 12633 25245 12667 25279
rect 13093 25245 13127 25279
rect 13185 25245 13219 25279
rect 13369 25245 13403 25279
rect 13461 25245 13495 25279
rect 13553 25245 13587 25279
rect 13737 25245 13771 25279
rect 15301 25245 15335 25279
rect 16129 25245 16163 25279
rect 16589 25245 16623 25279
rect 16773 25245 16807 25279
rect 21373 25245 21407 25279
rect 21649 25245 21683 25279
rect 21925 25245 21959 25279
rect 23213 25245 23247 25279
rect 23397 25245 23431 25279
rect 23673 25245 23707 25279
rect 23949 25245 23983 25279
rect 24041 25245 24075 25279
rect 24409 25245 24443 25279
rect 24685 25245 24719 25279
rect 25973 25245 26007 25279
rect 27629 25245 27663 25279
rect 27721 25245 27755 25279
rect 30481 25245 30515 25279
rect 31861 25245 31895 25279
rect 34529 25245 34563 25279
rect 9597 25177 9631 25211
rect 10425 25177 10459 25211
rect 15669 25177 15703 25211
rect 23305 25177 23339 25211
rect 23535 25177 23569 25211
rect 8769 25109 8803 25143
rect 10149 25109 10183 25143
rect 10701 25109 10735 25143
rect 12081 25109 12115 25143
rect 12909 25109 12943 25143
rect 15761 25109 15795 25143
rect 16221 25109 16255 25143
rect 20085 25109 20119 25143
rect 20453 25109 20487 25143
rect 20821 25109 20855 25143
rect 21281 25109 21315 25143
rect 21465 25109 21499 25143
rect 22293 25109 22327 25143
rect 24501 25109 24535 25143
rect 27353 25109 27387 25143
rect 30389 25109 30423 25143
rect 11345 24905 11379 24939
rect 15945 24905 15979 24939
rect 21373 24905 21407 24939
rect 21649 24905 21683 24939
rect 22845 24905 22879 24939
rect 23305 24905 23339 24939
rect 24869 24905 24903 24939
rect 29653 24905 29687 24939
rect 34897 24905 34931 24939
rect 20729 24837 20763 24871
rect 21281 24837 21315 24871
rect 22661 24837 22695 24871
rect 22937 24837 22971 24871
rect 24685 24837 24719 24871
rect 8033 24769 8067 24803
rect 8217 24769 8251 24803
rect 8677 24769 8711 24803
rect 9045 24769 9079 24803
rect 9413 24769 9447 24803
rect 11161 24769 11195 24803
rect 12081 24769 12115 24803
rect 15669 24769 15703 24803
rect 15761 24769 15795 24803
rect 16037 24769 16071 24803
rect 19165 24769 19199 24803
rect 19993 24769 20027 24803
rect 21465 24769 21499 24803
rect 23029 24769 23063 24803
rect 23489 24769 23523 24803
rect 23765 24769 23799 24803
rect 23949 24769 23983 24803
rect 24041 24769 24075 24803
rect 24225 24769 24259 24803
rect 24317 24769 24351 24803
rect 25145 24769 25179 24803
rect 25329 24769 25363 24803
rect 25697 24769 25731 24803
rect 25881 24769 25915 24803
rect 26249 24769 26283 24803
rect 26433 24769 26467 24803
rect 32321 24769 32355 24803
rect 32781 24769 32815 24803
rect 32973 24769 33007 24803
rect 10977 24701 11011 24735
rect 13461 24701 13495 24735
rect 15853 24701 15887 24735
rect 19073 24701 19107 24735
rect 19533 24701 19567 24735
rect 19809 24701 19843 24735
rect 23213 24701 23247 24735
rect 25513 24701 25547 24735
rect 32413 24701 32447 24735
rect 32873 24701 32907 24735
rect 33149 24701 33183 24735
rect 33425 24701 33459 24735
rect 8769 24633 8803 24667
rect 21097 24633 21131 24667
rect 22109 24633 22143 24667
rect 25145 24633 25179 24667
rect 32689 24633 32723 24667
rect 10701 24565 10735 24599
rect 11805 24565 11839 24599
rect 13829 24565 13863 24599
rect 22477 24565 22511 24599
rect 24225 24565 24259 24599
rect 24685 24565 24719 24599
rect 26617 24565 26651 24599
rect 10517 24361 10551 24395
rect 11437 24361 11471 24395
rect 14105 24361 14139 24395
rect 15301 24361 15335 24395
rect 16589 24361 16623 24395
rect 17049 24361 17083 24395
rect 17233 24361 17267 24395
rect 22569 24361 22603 24395
rect 28181 24361 28215 24395
rect 31585 24361 31619 24395
rect 34253 24361 34287 24395
rect 12173 24293 12207 24327
rect 12909 24293 12943 24327
rect 14565 24293 14599 24327
rect 20637 24293 20671 24327
rect 21005 24293 21039 24327
rect 27077 24293 27111 24327
rect 27997 24293 28031 24327
rect 9229 24225 9263 24259
rect 10425 24225 10459 24259
rect 11529 24225 11563 24259
rect 15669 24225 15703 24259
rect 16405 24225 16439 24259
rect 18245 24225 18279 24259
rect 27169 24225 27203 24259
rect 28549 24225 28583 24259
rect 29101 24225 29135 24259
rect 29837 24225 29871 24259
rect 1409 24157 1443 24191
rect 3065 24157 3099 24191
rect 3985 24157 4019 24191
rect 10609 24157 10643 24191
rect 10885 24157 10919 24191
rect 10977 24157 11011 24191
rect 11161 24157 11195 24191
rect 11253 24157 11287 24191
rect 11805 24157 11839 24191
rect 11897 24157 11931 24191
rect 12265 24157 12299 24191
rect 12633 24157 12667 24191
rect 12909 24157 12943 24191
rect 13001 24157 13035 24191
rect 13486 24157 13520 24191
rect 14381 24157 14415 24191
rect 14473 24157 14507 24191
rect 14657 24157 14691 24191
rect 15485 24157 15519 24191
rect 15761 24157 15795 24191
rect 16497 24157 16531 24191
rect 17141 24157 17175 24191
rect 17325 24157 17359 24191
rect 25605 24157 25639 24191
rect 25789 24157 25823 24191
rect 26065 24157 26099 24191
rect 26249 24157 26283 24191
rect 26341 24157 26375 24191
rect 26709 24157 26743 24191
rect 26985 24157 27019 24191
rect 27445 24157 27479 24191
rect 27721 24157 27755 24191
rect 27905 24157 27939 24191
rect 28089 24157 28123 24191
rect 28365 24157 28399 24191
rect 28457 24157 28491 24191
rect 28641 24157 28675 24191
rect 29009 24157 29043 24191
rect 34161 24157 34195 24191
rect 10057 24089 10091 24123
rect 10333 24089 10367 24123
rect 10793 24089 10827 24123
rect 13277 24089 13311 24123
rect 14105 24089 14139 24123
rect 17417 24089 17451 24123
rect 21373 24089 21407 24123
rect 27261 24089 27295 24123
rect 30113 24089 30147 24123
rect 1593 24021 1627 24055
rect 2973 24021 3007 24055
rect 3433 24021 3467 24055
rect 8309 24021 8343 24055
rect 8585 24021 8619 24055
rect 11989 24021 12023 24055
rect 12725 24021 12759 24055
rect 13369 24021 13403 24055
rect 13645 24021 13679 24055
rect 14289 24021 14323 24055
rect 20177 24021 20211 24055
rect 21741 24021 21775 24055
rect 22201 24021 22235 24055
rect 23029 24021 23063 24055
rect 23397 24021 23431 24055
rect 27629 24021 27663 24055
rect 29377 24021 29411 24055
rect 32965 24021 32999 24055
rect 34069 24021 34103 24055
rect 11713 23817 11747 23851
rect 15301 23817 15335 23851
rect 17877 23817 17911 23851
rect 21557 23817 21591 23851
rect 22201 23817 22235 23851
rect 22569 23817 22603 23851
rect 24777 23817 24811 23851
rect 26985 23817 27019 23851
rect 27153 23817 27187 23851
rect 29009 23817 29043 23851
rect 29377 23817 29411 23851
rect 30849 23817 30883 23851
rect 1869 23749 1903 23783
rect 3709 23749 3743 23783
rect 9413 23749 9447 23783
rect 12633 23749 12667 23783
rect 17509 23749 17543 23783
rect 20361 23749 20395 23783
rect 20729 23749 20763 23783
rect 20821 23749 20855 23783
rect 24961 23749 24995 23783
rect 25145 23749 25179 23783
rect 27353 23749 27387 23783
rect 27537 23749 27571 23783
rect 28365 23749 28399 23783
rect 3433 23681 3467 23715
rect 5457 23681 5491 23715
rect 6193 23681 6227 23715
rect 6469 23681 6503 23715
rect 8585 23681 8619 23715
rect 9781 23681 9815 23715
rect 9965 23681 9999 23715
rect 11529 23681 11563 23715
rect 11713 23681 11747 23715
rect 12817 23681 12851 23715
rect 12909 23681 12943 23715
rect 13737 23681 13771 23715
rect 13829 23681 13863 23715
rect 15485 23681 15519 23715
rect 15577 23681 15611 23715
rect 15761 23681 15795 23715
rect 15853 23681 15887 23715
rect 16865 23681 16899 23715
rect 17693 23681 17727 23715
rect 17877 23681 17911 23715
rect 20269 23681 20303 23715
rect 20453 23681 20487 23715
rect 20545 23681 20579 23715
rect 20913 23681 20947 23715
rect 22201 23681 22235 23715
rect 22477 23681 22511 23715
rect 22661 23681 22695 23715
rect 22753 23681 22787 23715
rect 22937 23681 22971 23715
rect 23213 23681 23247 23715
rect 24593 23681 24627 23715
rect 24869 23681 24903 23715
rect 27629 23681 27663 23715
rect 28549 23681 28583 23715
rect 28825 23681 28859 23715
rect 29009 23681 29043 23715
rect 29101 23681 29135 23715
rect 29285 23681 29319 23715
rect 29377 23681 29411 23715
rect 29561 23681 29595 23715
rect 30757 23681 30791 23715
rect 1593 23613 1627 23647
rect 5365 23613 5399 23647
rect 6745 23613 6779 23647
rect 8217 23613 8251 23647
rect 14013 23613 14047 23647
rect 16773 23613 16807 23647
rect 18153 23613 18187 23647
rect 21833 23613 21867 23647
rect 22385 23613 22419 23647
rect 28733 23613 28767 23647
rect 5825 23545 5859 23579
rect 12909 23545 12943 23579
rect 21097 23545 21131 23579
rect 29101 23545 29135 23579
rect 3341 23477 3375 23511
rect 5181 23477 5215 23511
rect 9781 23477 9815 23511
rect 10425 23477 10459 23511
rect 10793 23477 10827 23511
rect 11161 23477 11195 23511
rect 12081 23477 12115 23511
rect 13921 23477 13955 23511
rect 17141 23477 17175 23511
rect 19901 23477 19935 23511
rect 22845 23477 22879 23511
rect 23581 23477 23615 23511
rect 24409 23477 24443 23511
rect 25329 23477 25363 23511
rect 27169 23477 27203 23511
rect 30665 23477 30699 23511
rect 3433 23273 3467 23307
rect 4537 23273 4571 23307
rect 8309 23273 8343 23307
rect 13829 23273 13863 23307
rect 15117 23273 15151 23307
rect 16221 23273 16255 23307
rect 19717 23273 19751 23307
rect 20177 23273 20211 23307
rect 22017 23273 22051 23307
rect 22201 23273 22235 23307
rect 22293 23273 22327 23307
rect 22569 23273 22603 23307
rect 23397 23273 23431 23307
rect 24501 23273 24535 23307
rect 24593 23273 24627 23307
rect 4261 23205 4295 23239
rect 15669 23205 15703 23239
rect 17601 23205 17635 23239
rect 21097 23205 21131 23239
rect 1685 23137 1719 23171
rect 5273 23137 5307 23171
rect 6377 23137 6411 23171
rect 8125 23137 8159 23171
rect 9137 23137 9171 23171
rect 15025 23137 15059 23171
rect 15853 23137 15887 23171
rect 17141 23137 17175 23171
rect 18245 23137 18279 23171
rect 20821 23137 20855 23171
rect 21465 23137 21499 23171
rect 22109 23107 22143 23141
rect 23029 23137 23063 23171
rect 23765 23137 23799 23171
rect 24409 23137 24443 23171
rect 25789 23137 25823 23171
rect 34069 23137 34103 23171
rect 1409 23069 1443 23103
rect 4445 23069 4479 23103
rect 5181 23069 5215 23103
rect 8401 23069 8435 23103
rect 8677 23069 8711 23103
rect 8953 23069 8987 23103
rect 10057 23069 10091 23103
rect 10241 23069 10275 23103
rect 15544 23069 15578 23103
rect 15945 23069 15979 23103
rect 17233 23069 17267 23103
rect 18429 23069 18463 23103
rect 18613 23069 18647 23103
rect 19533 23069 19567 23103
rect 20729 23069 20763 23103
rect 20913 23069 20947 23103
rect 21005 23069 21039 23103
rect 21189 23069 21223 23103
rect 21649 23069 21683 23103
rect 22385 23069 22419 23103
rect 22753 23069 22787 23103
rect 22845 23069 22879 23103
rect 23121 23069 23155 23103
rect 23949 23069 23983 23103
rect 24225 23069 24259 23103
rect 24685 23069 24719 23103
rect 24869 23069 24903 23103
rect 25053 23069 25087 23103
rect 34529 23069 34563 23103
rect 6653 23001 6687 23035
rect 18705 23001 18739 23035
rect 18889 23001 18923 23035
rect 19073 23001 19107 23035
rect 19257 23001 19291 23035
rect 23213 23001 23247 23035
rect 24133 23001 24167 23035
rect 3157 22933 3191 22967
rect 5549 22933 5583 22967
rect 13093 22933 13127 22967
rect 14381 22933 14415 22967
rect 15485 22933 15519 22967
rect 19349 22933 19383 22967
rect 20637 22933 20671 22967
rect 21557 22933 21591 22967
rect 23413 22933 23447 22967
rect 23581 22933 23615 22967
rect 2237 22729 2271 22763
rect 7573 22729 7607 22763
rect 8125 22729 8159 22763
rect 10977 22729 11011 22763
rect 12449 22729 12483 22763
rect 15117 22729 15151 22763
rect 15393 22729 15427 22763
rect 15853 22729 15887 22763
rect 21005 22729 21039 22763
rect 21833 22729 21867 22763
rect 22661 22729 22695 22763
rect 23505 22729 23539 22763
rect 24961 22729 24995 22763
rect 29929 22729 29963 22763
rect 32689 22729 32723 22763
rect 34897 22729 34931 22763
rect 2881 22661 2915 22695
rect 13553 22661 13587 22695
rect 13645 22661 13679 22695
rect 22477 22661 22511 22695
rect 23305 22661 23339 22695
rect 23949 22661 23983 22695
rect 33425 22661 33459 22695
rect 2145 22593 2179 22627
rect 7389 22593 7423 22627
rect 7665 22593 7699 22627
rect 9045 22593 9079 22627
rect 9873 22593 9907 22627
rect 10149 22593 10183 22627
rect 12725 22593 12759 22627
rect 12817 22593 12851 22627
rect 13461 22593 13495 22627
rect 13829 22593 13863 22627
rect 13921 22593 13955 22627
rect 14105 22593 14139 22627
rect 15301 22593 15335 22627
rect 15485 22593 15519 22627
rect 18613 22593 18647 22627
rect 20729 22593 20763 22627
rect 22109 22593 22143 22627
rect 22569 22593 22603 22627
rect 22753 22593 22787 22627
rect 24593 22593 24627 22627
rect 27721 22593 27755 22627
rect 30113 22593 30147 22627
rect 32321 22593 32355 22627
rect 32781 22593 32815 22627
rect 32965 22593 32999 22627
rect 2605 22525 2639 22559
rect 4353 22525 4387 22559
rect 18521 22525 18555 22559
rect 22017 22525 22051 22559
rect 22385 22525 22419 22559
rect 24501 22525 24535 22559
rect 27997 22525 28031 22559
rect 30389 22525 30423 22559
rect 31861 22525 31895 22559
rect 32413 22525 32447 22559
rect 32873 22525 32907 22559
rect 33149 22525 33183 22559
rect 9965 22457 9999 22491
rect 11989 22457 12023 22491
rect 12541 22457 12575 22491
rect 14565 22457 14599 22491
rect 18981 22457 19015 22491
rect 21557 22457 21591 22491
rect 23673 22457 23707 22491
rect 2053 22389 2087 22423
rect 4721 22389 4755 22423
rect 8677 22389 8711 22423
rect 9413 22389 9447 22423
rect 9781 22389 9815 22423
rect 10609 22389 10643 22423
rect 13277 22389 13311 22423
rect 14289 22389 14323 22423
rect 23121 22389 23155 22423
rect 23489 22389 23523 22423
rect 27537 22389 27571 22423
rect 27905 22389 27939 22423
rect 3893 22185 3927 22219
rect 4813 22185 4847 22219
rect 5181 22185 5215 22219
rect 5825 22185 5859 22219
rect 10425 22185 10459 22219
rect 15117 22185 15151 22219
rect 23029 22185 23063 22219
rect 30389 22185 30423 22219
rect 30941 22185 30975 22219
rect 34253 22185 34287 22219
rect 5089 22117 5123 22151
rect 8769 22117 8803 22151
rect 10793 22117 10827 22151
rect 13093 22117 13127 22151
rect 18061 22117 18095 22151
rect 26249 22117 26283 22151
rect 26341 22117 26375 22151
rect 5273 22049 5307 22083
rect 10149 22049 10183 22083
rect 10701 22049 10735 22083
rect 17601 22049 17635 22083
rect 20545 22049 20579 22083
rect 21741 22049 21775 22083
rect 22477 22049 22511 22083
rect 25973 22049 26007 22083
rect 27537 22049 27571 22083
rect 28365 22049 28399 22083
rect 28825 22049 28859 22083
rect 31861 22049 31895 22083
rect 1409 21981 1443 22015
rect 3985 21981 4019 22015
rect 4261 21981 4295 22015
rect 4997 21981 5031 22015
rect 5365 21981 5399 22015
rect 5549 21981 5583 22015
rect 5641 21981 5675 22015
rect 5825 21981 5859 22015
rect 5917 21981 5951 22015
rect 7757 21981 7791 22015
rect 8033 21981 8067 22015
rect 9137 21981 9171 22015
rect 9413 21981 9447 22015
rect 9689 21981 9723 22015
rect 9873 21981 9907 22015
rect 10241 21981 10275 22015
rect 10885 21981 10919 22015
rect 11161 21981 11195 22015
rect 11529 21981 11563 22015
rect 11897 21981 11931 22015
rect 11989 21981 12023 22015
rect 12449 21981 12483 22015
rect 12817 21981 12851 22015
rect 14105 21981 14139 22015
rect 14197 21981 14231 22015
rect 14565 21981 14599 22015
rect 15117 21981 15151 22015
rect 15393 21981 15427 22015
rect 17693 21981 17727 22015
rect 19533 21981 19567 22015
rect 19901 21981 19935 22015
rect 21189 21981 21223 22015
rect 21281 21981 21315 22015
rect 26433 21981 26467 22015
rect 26709 21981 26743 22015
rect 26893 21981 26927 22015
rect 27353 21981 27387 22015
rect 27813 21981 27847 22015
rect 27905 21981 27939 22015
rect 28089 21981 28123 22015
rect 28181 21981 28215 22015
rect 28457 21981 28491 22015
rect 30113 21981 30147 22015
rect 30205 21981 30239 22015
rect 30849 21981 30883 22015
rect 32045 21981 32079 22015
rect 34161 21981 34195 22015
rect 13461 21913 13495 21947
rect 13921 21913 13955 21947
rect 14381 21913 14415 21947
rect 14473 21913 14507 21947
rect 21373 21913 21407 21947
rect 27031 21913 27065 21947
rect 27169 21913 27203 21947
rect 27261 21913 27295 21947
rect 27629 21913 27663 21947
rect 29745 21913 29779 21947
rect 29929 21913 29963 21947
rect 32229 21913 32263 21947
rect 1593 21845 1627 21879
rect 6193 21845 6227 21879
rect 7665 21845 7699 21879
rect 7849 21845 7883 21879
rect 8125 21845 8159 21879
rect 9229 21845 9263 21879
rect 9597 21845 9631 21879
rect 11069 21845 11103 21879
rect 14749 21845 14783 21879
rect 15301 21845 15335 21879
rect 26617 21845 26651 21879
rect 30665 21845 30699 21879
rect 32965 21845 32999 21879
rect 34069 21845 34103 21879
rect 4629 21641 4663 21675
rect 10977 21641 11011 21675
rect 12173 21641 12207 21675
rect 13553 21641 13587 21675
rect 14657 21641 14691 21675
rect 23121 21641 23155 21675
rect 26801 21641 26835 21675
rect 27169 21641 27203 21675
rect 27813 21641 27847 21675
rect 27997 21641 28031 21675
rect 29101 21641 29135 21675
rect 29370 21641 29404 21675
rect 3157 21573 3191 21607
rect 4813 21573 4847 21607
rect 4997 21573 5031 21607
rect 13185 21573 13219 21607
rect 14565 21573 14599 21607
rect 23397 21573 23431 21607
rect 28365 21573 28399 21607
rect 28733 21573 28767 21607
rect 28949 21573 28983 21607
rect 29469 21573 29503 21607
rect 2145 21505 2179 21539
rect 4905 21505 4939 21539
rect 5181 21505 5215 21539
rect 5273 21505 5307 21539
rect 5549 21505 5583 21539
rect 6009 21505 6043 21539
rect 6193 21505 6227 21539
rect 6377 21505 6411 21539
rect 6561 21505 6595 21539
rect 8861 21505 8895 21539
rect 9965 21505 9999 21539
rect 10793 21505 10827 21539
rect 10977 21505 11011 21539
rect 11529 21505 11563 21539
rect 11713 21505 11747 21539
rect 11897 21505 11931 21539
rect 11989 21505 12023 21539
rect 14841 21505 14875 21539
rect 15209 21505 15243 21539
rect 15393 21505 15427 21539
rect 15669 21505 15703 21539
rect 16865 21505 16899 21539
rect 19349 21505 19383 21539
rect 22937 21505 22971 21539
rect 23121 21505 23155 21539
rect 26525 21505 26559 21539
rect 27905 21505 27939 21539
rect 28181 21505 28215 21539
rect 29193 21505 29227 21539
rect 29285 21505 29319 21539
rect 2881 21437 2915 21471
rect 4997 21437 5031 21471
rect 5457 21437 5491 21471
rect 6101 21437 6135 21471
rect 7021 21437 7055 21471
rect 7297 21437 7331 21471
rect 8769 21437 8803 21471
rect 9505 21437 9539 21471
rect 10149 21437 10183 21471
rect 11805 21437 11839 21471
rect 15577 21437 15611 21471
rect 16957 21437 16991 21471
rect 17233 21437 17267 21471
rect 19441 21437 19475 21471
rect 22661 21437 22695 21471
rect 26341 21437 26375 21471
rect 26433 21437 26467 21471
rect 26617 21437 26651 21471
rect 19717 21369 19751 21403
rect 2237 21301 2271 21335
rect 2697 21301 2731 21335
rect 5825 21301 5859 21335
rect 6745 21301 6779 21335
rect 12633 21301 12667 21335
rect 15025 21301 15059 21335
rect 27445 21301 27479 21335
rect 27537 21301 27571 21335
rect 27629 21301 27663 21335
rect 28917 21301 28951 21335
rect 3433 21097 3467 21131
rect 4997 21097 5031 21131
rect 6653 21097 6687 21131
rect 8493 21097 8527 21131
rect 10241 21097 10275 21131
rect 10517 21097 10551 21131
rect 10793 21097 10827 21131
rect 11989 21097 12023 21131
rect 13093 21097 13127 21131
rect 13829 21097 13863 21131
rect 14289 21097 14323 21131
rect 20637 21097 20671 21131
rect 21833 21097 21867 21131
rect 22385 21097 22419 21131
rect 23581 21097 23615 21131
rect 24225 21097 24259 21131
rect 24869 21097 24903 21131
rect 26249 21097 26283 21131
rect 26709 21097 26743 21131
rect 11713 21029 11747 21063
rect 20085 21029 20119 21063
rect 22937 21029 22971 21063
rect 1685 20961 1719 20995
rect 10793 20961 10827 20995
rect 12909 20961 12943 20995
rect 13645 20961 13679 20995
rect 17785 20961 17819 20995
rect 18429 20961 18463 20995
rect 22109 20961 22143 20995
rect 22661 20961 22695 20995
rect 23397 20961 23431 20995
rect 23765 20961 23799 20995
rect 24501 20961 24535 20995
rect 26065 20961 26099 20995
rect 34069 20961 34103 20995
rect 1409 20893 1443 20927
rect 6469 20893 6503 20927
rect 6745 20893 6779 20927
rect 10885 20893 10919 20927
rect 11161 20893 11195 20927
rect 11253 20893 11287 20927
rect 11437 20893 11471 20927
rect 11805 20893 11839 20927
rect 11897 20893 11931 20927
rect 13277 20893 13311 20927
rect 13461 20893 13495 20927
rect 13553 20893 13587 20927
rect 13921 20893 13955 20927
rect 16681 20893 16715 20927
rect 16865 20893 16899 20927
rect 17141 20893 17175 20927
rect 17325 20893 17359 20927
rect 17417 20893 17451 20927
rect 17509 20893 17543 20927
rect 17877 20893 17911 20927
rect 18061 20893 18095 20927
rect 19809 20893 19843 20927
rect 20177 20893 20211 20927
rect 20545 20893 20579 20927
rect 20637 20893 20671 20927
rect 20729 20893 20763 20927
rect 22187 20893 22221 20927
rect 22577 20895 22611 20929
rect 22753 20893 22787 20927
rect 22845 20893 22879 20927
rect 23029 20893 23063 20927
rect 23673 20893 23707 20927
rect 23857 20893 23891 20927
rect 23981 20893 24015 20927
rect 24593 20893 24627 20927
rect 25789 20893 25823 20927
rect 25881 20893 25915 20927
rect 25973 20893 26007 20927
rect 26341 20893 26375 20927
rect 26525 20893 26559 20927
rect 34529 20893 34563 20927
rect 7021 20825 7055 20859
rect 13645 20825 13679 20859
rect 14257 20825 14291 20859
rect 14473 20825 14507 20859
rect 17049 20825 17083 20859
rect 23397 20825 23431 20859
rect 3157 20757 3191 20791
rect 9137 20757 9171 20791
rect 11069 20757 11103 20791
rect 12541 20757 12575 20791
rect 14105 20757 14139 20791
rect 18337 20757 18371 20791
rect 21005 20757 21039 20791
rect 25513 20757 25547 20791
rect 11345 20553 11379 20587
rect 13921 20553 13955 20587
rect 14013 20553 14047 20587
rect 17601 20553 17635 20587
rect 22477 20553 22511 20587
rect 23121 20553 23155 20587
rect 23581 20553 23615 20587
rect 24501 20553 24535 20587
rect 25329 20553 25363 20587
rect 28917 20553 28951 20587
rect 10977 20485 11011 20519
rect 11805 20485 11839 20519
rect 13461 20485 13495 20519
rect 14381 20485 14415 20519
rect 16497 20485 16531 20519
rect 16681 20485 16715 20519
rect 16865 20485 16899 20519
rect 24041 20485 24075 20519
rect 2237 20417 2271 20451
rect 3065 20417 3099 20451
rect 12081 20417 12115 20451
rect 12265 20417 12299 20451
rect 12541 20417 12575 20451
rect 13185 20417 13219 20451
rect 14289 20417 14323 20451
rect 14473 20417 14507 20451
rect 15301 20417 15335 20451
rect 17233 20417 17267 20451
rect 17417 20417 17451 20451
rect 20177 20417 20211 20451
rect 23581 20417 23615 20451
rect 25697 20417 25731 20451
rect 25973 20417 26007 20451
rect 27905 20417 27939 20451
rect 28457 20417 28491 20451
rect 11529 20349 11563 20383
rect 14749 20349 14783 20383
rect 15393 20349 15427 20383
rect 15669 20349 15703 20383
rect 20453 20349 20487 20383
rect 23857 20349 23891 20383
rect 27997 20349 28031 20383
rect 3341 20281 3375 20315
rect 13461 20281 13495 20315
rect 17049 20281 17083 20315
rect 20361 20281 20395 20315
rect 23673 20281 23707 20315
rect 24317 20281 24351 20315
rect 26249 20281 26283 20315
rect 2329 20213 2363 20247
rect 2789 20213 2823 20247
rect 2973 20213 3007 20247
rect 8677 20213 8711 20247
rect 9781 20213 9815 20247
rect 10241 20213 10275 20247
rect 10609 20213 10643 20247
rect 12725 20213 12759 20247
rect 13093 20213 13127 20247
rect 14197 20213 14231 20247
rect 16865 20213 16899 20247
rect 20269 20213 20303 20247
rect 22845 20213 22879 20247
rect 25881 20213 25915 20247
rect 28181 20213 28215 20247
rect 28549 20213 28583 20247
rect 10701 20009 10735 20043
rect 11069 20009 11103 20043
rect 11529 20009 11563 20043
rect 13185 20009 13219 20043
rect 13369 20009 13403 20043
rect 15301 20009 15335 20043
rect 15577 20009 15611 20043
rect 16681 20009 16715 20043
rect 17141 20009 17175 20043
rect 17601 20009 17635 20043
rect 17877 20009 17911 20043
rect 22661 20009 22695 20043
rect 23857 20009 23891 20043
rect 25789 20009 25823 20043
rect 34529 20009 34563 20043
rect 12633 19941 12667 19975
rect 14749 19941 14783 19975
rect 18613 19941 18647 19975
rect 20453 19941 20487 19975
rect 24041 19941 24075 19975
rect 27905 19941 27939 19975
rect 32597 19941 32631 19975
rect 2053 19873 2087 19907
rect 4261 19873 4295 19907
rect 4997 19873 5031 19907
rect 8493 19873 8527 19907
rect 11345 19873 11379 19907
rect 11713 19873 11747 19907
rect 12173 19873 12207 19907
rect 15117 19873 15151 19907
rect 17233 19873 17267 19907
rect 20269 19873 20303 19907
rect 20361 19873 20395 19907
rect 23121 19873 23155 19907
rect 23581 19873 23615 19907
rect 27077 19873 27111 19907
rect 28733 19873 28767 19907
rect 29745 19873 29779 19907
rect 31493 19873 31527 19907
rect 31861 19873 31895 19907
rect 32781 19873 32815 19907
rect 1409 19805 1443 19839
rect 1777 19805 1811 19839
rect 4169 19805 4203 19839
rect 5181 19805 5215 19839
rect 5273 19805 5307 19839
rect 7573 19805 7607 19839
rect 8585 19805 8619 19839
rect 10241 19805 10275 19839
rect 11253 19805 11287 19839
rect 11437 19805 11471 19839
rect 11805 19805 11839 19839
rect 12357 19805 12391 19839
rect 12449 19805 12483 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 13829 19805 13863 19839
rect 13921 19805 13955 19839
rect 15209 19805 15243 19839
rect 15393 19805 15427 19839
rect 15485 19805 15519 19839
rect 15669 19805 15703 19839
rect 16221 19805 16255 19839
rect 16497 19805 16531 19839
rect 16773 19805 16807 19839
rect 16957 19805 16991 19839
rect 17693 19805 17727 19839
rect 17785 19805 17819 19839
rect 19533 19805 19567 19839
rect 19809 19805 19843 19839
rect 20085 19805 20119 19839
rect 20637 19805 20671 19839
rect 20729 19805 20763 19839
rect 23029 19805 23063 19839
rect 23213 19805 23247 19839
rect 23489 19805 23523 19839
rect 23949 19805 23983 19839
rect 24133 19805 24167 19839
rect 25145 19805 25179 19839
rect 25421 19805 25455 19839
rect 25605 19805 25639 19839
rect 25697 19805 25731 19839
rect 25881 19805 25915 19839
rect 26065 19805 26099 19839
rect 26249 19805 26283 19839
rect 27632 19783 27666 19817
rect 28825 19805 28859 19839
rect 31953 19805 31987 19839
rect 34713 19805 34747 19839
rect 9045 19737 9079 19771
rect 9873 19737 9907 19771
rect 12633 19737 12667 19771
rect 17969 19737 18003 19771
rect 20453 19737 20487 19771
rect 24593 19737 24627 19771
rect 25513 19737 25547 19771
rect 27905 19737 27939 19771
rect 30021 19737 30055 19771
rect 33057 19737 33091 19771
rect 34805 19737 34839 19771
rect 1593 19669 1627 19703
rect 3525 19669 3559 19703
rect 4537 19669 4571 19703
rect 4997 19669 5031 19703
rect 7665 19669 7699 19703
rect 8033 19669 8067 19703
rect 8769 19669 8803 19703
rect 10149 19669 10183 19703
rect 14289 19669 14323 19703
rect 16129 19669 16163 19703
rect 16313 19669 16347 19703
rect 27721 19669 27755 19703
rect 29193 19669 29227 19703
rect 32321 19669 32355 19703
rect 4261 19465 4295 19499
rect 4721 19465 4755 19499
rect 5273 19465 5307 19499
rect 11805 19465 11839 19499
rect 12817 19465 12851 19499
rect 13277 19465 13311 19499
rect 16129 19465 16163 19499
rect 18245 19465 18279 19499
rect 18613 19465 18647 19499
rect 20177 19465 20211 19499
rect 20913 19465 20947 19499
rect 21649 19465 21683 19499
rect 22033 19465 22067 19499
rect 22845 19465 22879 19499
rect 23581 19465 23615 19499
rect 26157 19465 26191 19499
rect 29653 19465 29687 19499
rect 30757 19465 30791 19499
rect 31953 19465 31987 19499
rect 32505 19465 32539 19499
rect 8493 19397 8527 19431
rect 9137 19397 9171 19431
rect 11253 19397 11287 19431
rect 12449 19397 12483 19431
rect 16405 19397 16439 19431
rect 21281 19397 21315 19431
rect 21833 19397 21867 19431
rect 22385 19397 22419 19431
rect 25605 19397 25639 19431
rect 1409 19329 1443 19363
rect 3985 19329 4019 19363
rect 4353 19329 4387 19363
rect 5089 19329 5123 19363
rect 5549 19329 5583 19363
rect 6561 19329 6595 19363
rect 8585 19329 8619 19363
rect 10885 19329 10919 19363
rect 17417 19329 17451 19363
rect 18797 19329 18831 19363
rect 18889 19329 18923 19363
rect 18981 19329 19015 19363
rect 19165 19329 19199 19363
rect 19533 19329 19567 19363
rect 19717 19329 19751 19363
rect 19809 19329 19843 19363
rect 19901 19329 19935 19363
rect 20821 19329 20855 19363
rect 21097 19329 21131 19363
rect 21373 19329 21407 19363
rect 21557 19329 21591 19363
rect 21649 19329 21683 19363
rect 22293 19329 22327 19363
rect 22569 19329 22603 19363
rect 25237 19329 25271 19363
rect 25881 19329 25915 19363
rect 30665 19329 30699 19363
rect 31677 19329 31711 19363
rect 32137 19329 32171 19363
rect 1685 19261 1719 19295
rect 4261 19261 4295 19295
rect 4445 19261 4479 19295
rect 4905 19261 4939 19295
rect 5641 19261 5675 19295
rect 6837 19261 6871 19295
rect 8861 19261 8895 19295
rect 15117 19261 15151 19295
rect 17049 19261 17083 19295
rect 18429 19261 18463 19295
rect 18521 19261 18555 19295
rect 25605 19261 25639 19295
rect 26525 19261 26559 19295
rect 31953 19261 31987 19295
rect 32229 19261 32263 19295
rect 3617 19193 3651 19227
rect 4077 19193 4111 19227
rect 5917 19193 5951 19227
rect 17693 19193 17727 19227
rect 19073 19193 19107 19227
rect 24777 19193 24811 19227
rect 31769 19193 31803 19227
rect 3157 19125 3191 19159
rect 4445 19125 4479 19159
rect 8309 19125 8343 19159
rect 18153 19125 18187 19159
rect 22017 19125 22051 19159
rect 22201 19125 22235 19159
rect 22569 19125 22603 19159
rect 24317 19125 24351 19159
rect 25789 19125 25823 19159
rect 30481 19125 30515 19159
rect 32137 19125 32171 19159
rect 34253 19125 34287 19159
rect 34529 19125 34563 19159
rect 5549 18921 5583 18955
rect 8309 18921 8343 18955
rect 10977 18921 11011 18955
rect 17601 18921 17635 18955
rect 22477 18921 22511 18955
rect 23397 18921 23431 18955
rect 24869 18921 24903 18955
rect 26709 18921 26743 18955
rect 12817 18853 12851 18887
rect 18889 18853 18923 18887
rect 21925 18853 21959 18887
rect 22937 18853 22971 18887
rect 23765 18853 23799 18887
rect 28457 18853 28491 18887
rect 6837 18785 6871 18819
rect 17141 18785 17175 18819
rect 18337 18785 18371 18819
rect 22385 18785 22419 18819
rect 23489 18785 23523 18819
rect 25814 18785 25848 18819
rect 26985 18785 27019 18819
rect 27997 18785 28031 18819
rect 28365 18785 28399 18819
rect 28825 18785 28859 18819
rect 31309 18785 31343 18819
rect 32045 18785 32079 18819
rect 32505 18785 32539 18819
rect 32781 18785 32815 18819
rect 3341 18717 3375 18751
rect 3433 18717 3467 18751
rect 4261 18717 4295 18751
rect 5273 18717 5307 18751
rect 5365 18717 5399 18751
rect 6561 18717 6595 18751
rect 9321 18717 9355 18751
rect 10609 18717 10643 18751
rect 11437 18717 11471 18751
rect 11621 18717 11655 18751
rect 12081 18717 12115 18751
rect 13277 18717 13311 18751
rect 13553 18717 13587 18751
rect 13645 18717 13679 18751
rect 17233 18717 17267 18751
rect 17325 18717 17359 18751
rect 17417 18717 17451 18751
rect 17693 18717 17727 18751
rect 17877 18717 17911 18751
rect 18153 18717 18187 18751
rect 18521 18717 18555 18751
rect 20637 18717 20671 18751
rect 20913 18717 20947 18751
rect 21281 18717 21315 18751
rect 21649 18717 21683 18751
rect 22017 18717 22051 18751
rect 22661 18717 22695 18751
rect 22753 18717 22787 18751
rect 23268 18717 23302 18751
rect 24409 18717 24443 18751
rect 24501 18717 24535 18751
rect 24685 18717 24719 18751
rect 25329 18717 25363 18751
rect 26065 18717 26099 18751
rect 26249 18717 26283 18751
rect 26525 18717 26559 18751
rect 27905 18717 27939 18751
rect 29377 18717 29411 18751
rect 29561 18717 29595 18751
rect 31953 18717 31987 18751
rect 32413 18717 32447 18751
rect 32597 18717 32631 18751
rect 34713 18717 34747 18751
rect 3617 18649 3651 18683
rect 4077 18649 4111 18683
rect 9873 18649 9907 18683
rect 11713 18649 11747 18683
rect 13369 18649 13403 18683
rect 23121 18649 23155 18683
rect 29837 18649 29871 18683
rect 33057 18649 33091 18683
rect 34805 18649 34839 18683
rect 3065 18581 3099 18615
rect 8677 18581 8711 18615
rect 10241 18581 10275 18615
rect 12449 18581 12483 18615
rect 24133 18581 24167 18615
rect 25237 18581 25271 18615
rect 25605 18581 25639 18615
rect 25697 18581 25731 18615
rect 25973 18581 26007 18615
rect 28273 18581 28307 18615
rect 32321 18581 32355 18615
rect 34529 18581 34563 18615
rect 14105 18377 14139 18411
rect 17877 18377 17911 18411
rect 21649 18377 21683 18411
rect 23397 18377 23431 18411
rect 24225 18377 24259 18411
rect 24869 18377 24903 18411
rect 25697 18377 25731 18411
rect 30297 18377 30331 18411
rect 13185 18309 13219 18343
rect 13645 18309 13679 18343
rect 13737 18309 13771 18343
rect 14013 18309 14047 18343
rect 15669 18309 15703 18343
rect 17693 18309 17727 18343
rect 18245 18309 18279 18343
rect 23857 18309 23891 18343
rect 24073 18309 24107 18343
rect 25789 18309 25823 18343
rect 4813 18241 4847 18275
rect 5273 18241 5307 18275
rect 5457 18241 5491 18275
rect 10517 18241 10551 18275
rect 10977 18241 11011 18275
rect 11253 18241 11287 18275
rect 11345 18241 11379 18275
rect 12817 18241 12851 18275
rect 13001 18241 13035 18275
rect 13093 18241 13127 18275
rect 13277 18241 13311 18275
rect 13507 18241 13541 18275
rect 13829 18241 13863 18275
rect 14289 18241 14323 18275
rect 14565 18241 14599 18275
rect 14657 18241 14691 18275
rect 14841 18241 14875 18275
rect 15209 18241 15243 18275
rect 15301 18241 15335 18275
rect 15485 18241 15519 18275
rect 15761 18241 15795 18275
rect 15853 18241 15887 18275
rect 16037 18241 16071 18275
rect 16221 18241 16255 18275
rect 17049 18241 17083 18275
rect 17233 18241 17267 18275
rect 17509 18241 17543 18275
rect 17601 18241 17635 18275
rect 17969 18241 18003 18275
rect 19717 18241 19751 18275
rect 20361 18241 20395 18275
rect 21373 18241 21407 18275
rect 21465 18241 21499 18275
rect 24317 18241 24351 18275
rect 24501 18241 24535 18275
rect 25881 18241 25915 18275
rect 30205 18241 30239 18275
rect 34713 18241 34747 18275
rect 4905 18173 4939 18207
rect 5365 18173 5399 18207
rect 11805 18173 11839 18207
rect 12633 18173 12667 18207
rect 13369 18173 13403 18207
rect 14381 18173 14415 18207
rect 15025 18173 15059 18207
rect 17141 18173 17175 18207
rect 18061 18173 18095 18207
rect 18245 18173 18279 18207
rect 25421 18173 25455 18207
rect 34437 18173 34471 18207
rect 5181 18105 5215 18139
rect 8401 18105 8435 18139
rect 10885 18105 10919 18139
rect 12909 18105 12943 18139
rect 17325 18105 17359 18139
rect 20729 18105 20763 18139
rect 23765 18105 23799 18139
rect 8769 18037 8803 18071
rect 9137 18037 9171 18071
rect 14289 18037 14323 18071
rect 24041 18037 24075 18071
rect 24409 18037 24443 18071
rect 25237 18037 25271 18071
rect 26157 18037 26191 18071
rect 30021 18037 30055 18071
rect 32689 18037 32723 18071
rect 5181 17833 5215 17867
rect 13645 17833 13679 17867
rect 14197 17833 14231 17867
rect 14657 17833 14691 17867
rect 15209 17833 15243 17867
rect 15393 17833 15427 17867
rect 16497 17833 16531 17867
rect 16773 17833 16807 17867
rect 17141 17833 17175 17867
rect 20637 17833 20671 17867
rect 23213 17833 23247 17867
rect 23765 17833 23799 17867
rect 24225 17833 24259 17867
rect 25145 17833 25179 17867
rect 25881 17833 25915 17867
rect 26617 17833 26651 17867
rect 1685 17697 1719 17731
rect 6469 17697 6503 17731
rect 9229 17697 9263 17731
rect 11437 17697 11471 17731
rect 13553 17697 13587 17731
rect 18153 17697 18187 17731
rect 19073 17697 19107 17731
rect 20361 17697 20395 17731
rect 1409 17629 1443 17663
rect 8493 17629 8527 17663
rect 8953 17629 8987 17663
rect 11713 17629 11747 17663
rect 13737 17629 13771 17663
rect 13829 17629 13863 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 14933 17629 14967 17663
rect 15301 17629 15335 17663
rect 15577 17629 15611 17663
rect 15669 17629 15703 17663
rect 15853 17629 15887 17663
rect 15945 17629 15979 17663
rect 16037 17629 16071 17663
rect 16313 17629 16347 17663
rect 16773 17629 16807 17663
rect 16957 17629 16991 17663
rect 18337 17629 18371 17663
rect 19349 17629 19383 17663
rect 19533 17629 19567 17663
rect 20545 17629 20579 17663
rect 20729 17629 20763 17663
rect 4997 17561 5031 17595
rect 6745 17561 6779 17595
rect 8401 17561 8435 17595
rect 10977 17561 11011 17595
rect 16129 17561 16163 17595
rect 3157 17493 3191 17527
rect 3433 17493 3467 17527
rect 5197 17493 5231 17527
rect 5365 17493 5399 17527
rect 8217 17493 8251 17527
rect 10701 17493 10735 17527
rect 12357 17493 12391 17527
rect 12725 17493 12759 17527
rect 13461 17493 13495 17527
rect 15025 17493 15059 17527
rect 15117 17493 15151 17527
rect 22937 17493 22971 17527
rect 25513 17493 25547 17527
rect 26249 17493 26283 17527
rect 2329 17289 2363 17323
rect 4353 17289 4387 17323
rect 9965 17289 9999 17323
rect 15945 17289 15979 17323
rect 17601 17289 17635 17323
rect 21833 17289 21867 17323
rect 8769 17221 8803 17255
rect 11345 17221 11379 17255
rect 17417 17221 17451 17255
rect 22385 17221 22419 17255
rect 23305 17221 23339 17255
rect 25237 17221 25271 17255
rect 26249 17221 26283 17255
rect 26709 17221 26743 17255
rect 1409 17153 1443 17187
rect 2237 17153 2271 17187
rect 3433 17153 3467 17187
rect 3893 17153 3927 17187
rect 4169 17153 4203 17187
rect 5273 17153 5307 17187
rect 6377 17153 6411 17187
rect 8217 17153 8251 17187
rect 8493 17153 8527 17187
rect 9873 17153 9907 17187
rect 10333 17153 10367 17187
rect 10793 17153 10827 17187
rect 11069 17153 11103 17187
rect 11161 17153 11195 17187
rect 11621 17153 11655 17187
rect 13645 17153 13679 17187
rect 14013 17153 14047 17187
rect 14289 17153 14323 17187
rect 14657 17153 14691 17187
rect 14933 17153 14967 17187
rect 15209 17153 15243 17187
rect 15577 17153 15611 17187
rect 16037 17153 16071 17187
rect 16221 17153 16255 17187
rect 16773 17153 16807 17187
rect 16957 17153 16991 17187
rect 17233 17153 17267 17187
rect 17785 17153 17819 17187
rect 18153 17153 18187 17187
rect 20821 17153 20855 17187
rect 22109 17153 22143 17187
rect 22569 17153 22603 17187
rect 22753 17153 22787 17187
rect 22937 17153 22971 17187
rect 23213 17153 23247 17187
rect 23397 17153 23431 17187
rect 23673 17153 23707 17187
rect 23765 17153 23799 17187
rect 23857 17153 23891 17187
rect 23995 17153 24029 17187
rect 24593 17153 24627 17187
rect 25973 17153 26007 17187
rect 26157 17153 26191 17187
rect 26341 17153 26375 17187
rect 26525 17153 26559 17187
rect 26801 17153 26835 17187
rect 26985 17153 27019 17187
rect 27077 17153 27111 17187
rect 27261 17153 27295 17187
rect 3525 17085 3559 17119
rect 4077 17085 4111 17119
rect 5365 17085 5399 17119
rect 5641 17085 5675 17119
rect 6653 17085 6687 17119
rect 8125 17085 8159 17119
rect 9505 17085 9539 17119
rect 12173 17085 12207 17119
rect 15485 17085 15519 17119
rect 15669 17085 15703 17119
rect 15761 17085 15795 17119
rect 16405 17085 16439 17119
rect 17509 17085 17543 17119
rect 18245 17085 18279 17119
rect 20729 17085 20763 17119
rect 21649 17085 21683 17119
rect 22017 17085 22051 17119
rect 22477 17085 22511 17119
rect 23489 17085 23523 17119
rect 24133 17085 24167 17119
rect 24501 17085 24535 17119
rect 3801 17017 3835 17051
rect 1593 16949 1627 16983
rect 2789 16949 2823 16983
rect 4169 16949 4203 16983
rect 13277 16949 13311 16983
rect 17785 16949 17819 16983
rect 24225 16949 24259 16983
rect 26801 16949 26835 16983
rect 27445 16949 27479 16983
rect 3801 16745 3835 16779
rect 7481 16745 7515 16779
rect 11529 16745 11563 16779
rect 11989 16745 12023 16779
rect 14749 16745 14783 16779
rect 16957 16745 16991 16779
rect 18061 16745 18095 16779
rect 19441 16745 19475 16779
rect 23765 16745 23799 16779
rect 24869 16745 24903 16779
rect 26065 16745 26099 16779
rect 27813 16745 27847 16779
rect 4169 16677 4203 16711
rect 10701 16677 10735 16711
rect 11161 16677 11195 16711
rect 17049 16677 17083 16711
rect 24685 16677 24719 16711
rect 26709 16677 26743 16711
rect 27445 16677 27479 16711
rect 13921 16609 13955 16643
rect 16589 16609 16623 16643
rect 22109 16609 22143 16643
rect 23397 16609 23431 16643
rect 27077 16609 27111 16643
rect 30021 16609 30055 16643
rect 3985 16541 4019 16575
rect 4077 16541 4111 16575
rect 4261 16541 4295 16575
rect 7389 16541 7423 16575
rect 14105 16541 14139 16575
rect 14197 16541 14231 16575
rect 14381 16541 14415 16575
rect 14565 16541 14599 16575
rect 16773 16541 16807 16575
rect 17233 16541 17267 16575
rect 17509 16541 17543 16575
rect 17693 16541 17727 16575
rect 19257 16541 19291 16575
rect 22385 16541 22419 16575
rect 23949 16541 23983 16575
rect 24133 16541 24167 16575
rect 25053 16541 25087 16575
rect 25237 16541 25271 16575
rect 25329 16541 25363 16575
rect 25421 16541 25455 16575
rect 25605 16541 25639 16575
rect 25881 16541 25915 16575
rect 25973 16541 26007 16575
rect 26157 16541 26191 16575
rect 26249 16541 26283 16575
rect 26433 16541 26467 16575
rect 29745 16541 29779 16575
rect 34529 16541 34563 16575
rect 11069 16473 11103 16507
rect 11529 16473 11563 16507
rect 14473 16473 14507 16507
rect 33609 16473 33643 16507
rect 7941 16405 7975 16439
rect 8309 16405 8343 16439
rect 9873 16405 9907 16439
rect 10333 16405 10367 16439
rect 11713 16405 11747 16439
rect 12449 16405 12483 16439
rect 13369 16405 13403 16439
rect 23029 16405 23063 16439
rect 25789 16405 25823 16439
rect 26249 16405 26283 16439
rect 29653 16405 29687 16439
rect 10609 16201 10643 16235
rect 11345 16201 11379 16235
rect 13737 16201 13771 16235
rect 15301 16201 15335 16235
rect 17325 16201 17359 16235
rect 18521 16201 18555 16235
rect 19165 16201 19199 16235
rect 19901 16201 19935 16235
rect 32505 16201 32539 16235
rect 33057 16201 33091 16235
rect 34897 16201 34931 16235
rect 8493 16133 8527 16167
rect 10149 16133 10183 16167
rect 12541 16133 12575 16167
rect 13553 16133 13587 16167
rect 19533 16133 19567 16167
rect 19625 16133 19659 16167
rect 20085 16133 20119 16167
rect 21005 16133 21039 16167
rect 28641 16133 28675 16167
rect 4445 16065 4479 16099
rect 5089 16065 5123 16099
rect 5365 16065 5399 16099
rect 10241 16065 10275 16099
rect 11713 16065 11747 16099
rect 11897 16065 11931 16099
rect 12265 16065 12299 16099
rect 12817 16065 12851 16099
rect 13921 16065 13955 16099
rect 14105 16065 14139 16099
rect 15209 16065 15243 16099
rect 15393 16065 15427 16099
rect 17785 16065 17819 16099
rect 17969 16065 18003 16099
rect 18061 16065 18095 16099
rect 18153 16065 18187 16099
rect 18337 16065 18371 16099
rect 18429 16065 18463 16099
rect 18705 16065 18739 16099
rect 18797 16065 18831 16099
rect 18889 16065 18923 16099
rect 19257 16065 19291 16099
rect 19405 16065 19439 16099
rect 19763 16065 19797 16099
rect 20269 16065 20303 16099
rect 20545 16065 20579 16099
rect 21189 16065 21223 16099
rect 21373 16065 21407 16099
rect 22017 16065 22051 16099
rect 23305 16065 23339 16099
rect 25421 16065 25455 16099
rect 25605 16065 25639 16099
rect 25973 16065 26007 16099
rect 26249 16065 26283 16099
rect 32137 16065 32171 16099
rect 32321 16065 32355 16099
rect 33149 16065 33183 16099
rect 4537 15997 4571 16031
rect 4905 15997 4939 16031
rect 8217 15997 8251 16031
rect 11989 15997 12023 16031
rect 12081 15997 12115 16031
rect 12725 15997 12759 16031
rect 13185 15997 13219 16031
rect 20453 15997 20487 16031
rect 21925 15997 21959 16031
rect 25513 15997 25547 16031
rect 26801 15997 26835 16031
rect 28273 15997 28307 16031
rect 28365 15997 28399 16031
rect 33425 15997 33459 16031
rect 5273 15929 5307 15963
rect 10977 15929 11011 15963
rect 12449 15929 12483 15963
rect 17693 15929 17727 15963
rect 18705 15929 18739 15963
rect 21373 15929 21407 15963
rect 4813 15861 4847 15895
rect 9965 15861 9999 15895
rect 16865 15861 16899 15895
rect 18981 15861 19015 15895
rect 20637 15861 20671 15895
rect 22385 15861 22419 15895
rect 24961 15861 24995 15895
rect 25237 15861 25271 15895
rect 30113 15861 30147 15895
rect 3341 15657 3375 15691
rect 5273 15657 5307 15691
rect 12265 15657 12299 15691
rect 12633 15657 12667 15691
rect 13185 15657 13219 15691
rect 13553 15657 13587 15691
rect 14749 15657 14783 15691
rect 15209 15657 15243 15691
rect 17509 15657 17543 15691
rect 18613 15657 18647 15691
rect 19441 15657 19475 15691
rect 25513 15657 25547 15691
rect 29285 15657 29319 15691
rect 32229 15657 32263 15691
rect 34161 15657 34195 15691
rect 13093 15589 13127 15623
rect 31309 15589 31343 15623
rect 6285 15521 6319 15555
rect 9597 15521 9631 15555
rect 9873 15521 9907 15555
rect 13277 15521 13311 15555
rect 13829 15521 13863 15555
rect 14381 15521 14415 15555
rect 14473 15521 14507 15555
rect 15209 15521 15243 15555
rect 16497 15521 16531 15555
rect 29561 15521 29595 15555
rect 32045 15521 32079 15555
rect 32505 15521 32539 15555
rect 1593 15453 1627 15487
rect 3617 15453 3651 15487
rect 4629 15453 4663 15487
rect 4813 15453 4847 15487
rect 6009 15453 6043 15487
rect 8033 15453 8067 15487
rect 12081 15453 12115 15487
rect 12909 15453 12943 15487
rect 13001 15453 13035 15487
rect 13369 15453 13403 15487
rect 14105 15453 14139 15487
rect 14289 15453 14323 15487
rect 14565 15453 14599 15487
rect 15025 15453 15059 15487
rect 15669 15453 15703 15487
rect 16129 15453 16163 15487
rect 17693 15453 17727 15487
rect 17877 15453 17911 15487
rect 19349 15453 19383 15487
rect 19533 15453 19567 15487
rect 19625 15453 19659 15487
rect 19809 15453 19843 15487
rect 23305 15453 23339 15487
rect 23581 15453 23615 15487
rect 26899 15453 26933 15487
rect 27077 15453 27111 15487
rect 31401 15453 31435 15487
rect 31953 15453 31987 15487
rect 32413 15453 32447 15487
rect 32597 15453 32631 15487
rect 34069 15453 34103 15487
rect 1869 15385 1903 15419
rect 3525 15385 3559 15419
rect 4997 15385 5031 15419
rect 5181 15385 5215 15419
rect 7941 15385 7975 15419
rect 11805 15385 11839 15419
rect 11897 15385 11931 15419
rect 12817 15385 12851 15419
rect 15301 15385 15335 15419
rect 18337 15385 18371 15419
rect 18981 15385 19015 15419
rect 20085 15385 20119 15419
rect 29837 15385 29871 15419
rect 31493 15385 31527 15419
rect 3985 15317 4019 15351
rect 7757 15317 7791 15351
rect 8401 15317 8435 15351
rect 8769 15317 8803 15351
rect 11345 15317 11379 15351
rect 14841 15317 14875 15351
rect 17049 15317 17083 15351
rect 17877 15317 17911 15351
rect 19717 15317 19751 15351
rect 21005 15317 21039 15351
rect 21373 15317 21407 15351
rect 23397 15317 23431 15351
rect 23765 15317 23799 15351
rect 25053 15317 25087 15351
rect 25973 15317 26007 15351
rect 27077 15317 27111 15351
rect 33885 15317 33919 15351
rect 1593 15113 1627 15147
rect 10701 15113 10735 15147
rect 14105 15113 14139 15147
rect 14289 15113 14323 15147
rect 22135 15113 22169 15147
rect 27629 15113 27663 15147
rect 32229 15113 32263 15147
rect 11253 15045 11287 15079
rect 15301 15045 15335 15079
rect 16497 15045 16531 15079
rect 19165 15045 19199 15079
rect 21465 15045 21499 15079
rect 21925 15045 21959 15079
rect 24409 15045 24443 15079
rect 1409 14977 1443 15011
rect 8125 14977 8159 15011
rect 10609 14977 10643 15011
rect 11621 14977 11655 15011
rect 12265 14977 12299 15011
rect 13737 14977 13771 15011
rect 14381 14977 14415 15011
rect 14933 14977 14967 15011
rect 15117 14977 15151 15011
rect 15485 14977 15519 15011
rect 16681 14977 16715 15011
rect 16773 14977 16807 15011
rect 16957 14977 16991 15011
rect 20729 14977 20763 15011
rect 21097 14977 21131 15011
rect 21281 14977 21315 15011
rect 22385 14977 22419 15011
rect 22477 14977 22511 15011
rect 22661 14977 22695 15011
rect 22753 14977 22787 15011
rect 23489 14977 23523 15011
rect 23857 14977 23891 15011
rect 24317 14977 24351 15011
rect 24593 14977 24627 15011
rect 24777 14977 24811 15011
rect 25145 14977 25179 15011
rect 26525 14977 26559 15011
rect 26709 14977 26743 15011
rect 26801 14977 26835 15011
rect 27169 14977 27203 15011
rect 27261 14977 27295 15011
rect 27721 14977 27755 15011
rect 27905 14977 27939 15011
rect 28181 14977 28215 15011
rect 28365 14977 28399 15011
rect 29837 14977 29871 15011
rect 31217 14977 31251 15011
rect 32413 14977 32447 15011
rect 32689 14977 32723 15011
rect 8953 14909 8987 14943
rect 13645 14909 13679 14943
rect 14841 14909 14875 14943
rect 23765 14909 23799 14943
rect 25053 14909 25087 14943
rect 26341 14909 26375 14943
rect 28089 14909 28123 14943
rect 10517 14841 10551 14875
rect 24225 14841 24259 14875
rect 26985 14841 27019 14875
rect 3525 14773 3559 14807
rect 17509 14773 17543 14807
rect 20453 14773 20487 14807
rect 22109 14773 22143 14807
rect 22293 14773 22327 14807
rect 22937 14773 22971 14807
rect 23029 14773 23063 14807
rect 23213 14773 23247 14807
rect 25513 14773 25547 14807
rect 28273 14773 28307 14807
rect 29653 14773 29687 14807
rect 29929 14773 29963 14807
rect 5089 14569 5123 14603
rect 5273 14569 5307 14603
rect 10701 14569 10735 14603
rect 12633 14569 12667 14603
rect 13921 14569 13955 14603
rect 16589 14569 16623 14603
rect 18889 14569 18923 14603
rect 21373 14569 21407 14603
rect 23949 14569 23983 14603
rect 32137 14569 32171 14603
rect 32965 14569 32999 14603
rect 4353 14501 4387 14535
rect 13001 14501 13035 14535
rect 13369 14501 13403 14535
rect 14565 14501 14599 14535
rect 15761 14501 15795 14535
rect 20913 14501 20947 14535
rect 22569 14501 22603 14535
rect 29285 14501 29319 14535
rect 4997 14433 5031 14467
rect 6561 14433 6595 14467
rect 8309 14433 8343 14467
rect 9229 14433 9263 14467
rect 16681 14433 16715 14467
rect 17877 14433 17911 14467
rect 20821 14433 20855 14467
rect 21741 14433 21775 14467
rect 22661 14433 22695 14467
rect 23029 14433 23063 14467
rect 26985 14433 27019 14467
rect 28089 14433 28123 14467
rect 29561 14433 29595 14467
rect 31677 14433 31711 14467
rect 31861 14433 31895 14467
rect 34069 14433 34103 14467
rect 3985 14365 4019 14399
rect 5089 14365 5123 14399
rect 8585 14365 8619 14399
rect 8953 14365 8987 14399
rect 16865 14365 16899 14399
rect 17233 14365 17267 14399
rect 17417 14365 17451 14399
rect 20177 14365 20211 14399
rect 20729 14365 20763 14399
rect 21005 14365 21039 14399
rect 21373 14365 21407 14399
rect 21557 14365 21591 14399
rect 21833 14365 21867 14399
rect 22293 14365 22327 14399
rect 23121 14365 23155 14399
rect 23397 14365 23431 14399
rect 23489 14365 23523 14399
rect 23673 14365 23707 14399
rect 23765 14365 23799 14399
rect 25513 14365 25547 14399
rect 25789 14365 25823 14399
rect 27169 14365 27203 14399
rect 27997 14365 28031 14399
rect 31585 14365 31619 14399
rect 34529 14365 34563 14399
rect 4813 14297 4847 14331
rect 6837 14297 6871 14331
rect 8493 14297 8527 14331
rect 17601 14297 17635 14331
rect 20269 14297 20303 14331
rect 20453 14297 20487 14331
rect 22569 14297 22603 14331
rect 29837 14297 29871 14331
rect 3893 14229 3927 14263
rect 11161 14229 11195 14263
rect 11529 14229 11563 14263
rect 15393 14229 15427 14263
rect 16129 14229 16163 14263
rect 17049 14229 17083 14263
rect 19441 14229 19475 14263
rect 20085 14229 20119 14263
rect 20354 14229 20388 14263
rect 20545 14229 20579 14263
rect 21189 14229 21223 14263
rect 22109 14229 22143 14263
rect 22385 14229 22419 14263
rect 23305 14229 23339 14263
rect 25697 14229 25731 14263
rect 25973 14229 26007 14263
rect 27353 14229 27387 14263
rect 28365 14229 28399 14263
rect 31309 14229 31343 14263
rect 31861 14229 31895 14263
rect 4353 14025 4387 14059
rect 9045 14025 9079 14059
rect 9781 14025 9815 14059
rect 10241 14025 10275 14059
rect 13645 14025 13679 14059
rect 14749 14025 14783 14059
rect 16129 14025 16163 14059
rect 23121 14025 23155 14059
rect 25145 14025 25179 14059
rect 26525 14025 26559 14059
rect 29285 14025 29319 14059
rect 34805 14025 34839 14059
rect 2881 13957 2915 13991
rect 17049 13957 17083 13991
rect 22017 13957 22051 13991
rect 22753 13957 22787 13991
rect 25237 13957 25271 13991
rect 22983 13923 23017 13957
rect 2605 13889 2639 13923
rect 5089 13889 5123 13923
rect 5365 13889 5399 13923
rect 5733 13889 5767 13923
rect 6561 13889 6595 13923
rect 6745 13889 6779 13923
rect 6837 13889 6871 13923
rect 9873 13889 9907 13923
rect 12449 13889 12483 13923
rect 14657 13889 14691 13923
rect 15945 13889 15979 13923
rect 16681 13889 16715 13923
rect 16865 13889 16899 13923
rect 17417 13889 17451 13923
rect 17601 13889 17635 13923
rect 19257 13889 19291 13923
rect 19441 13889 19475 13923
rect 19809 13889 19843 13923
rect 19993 13889 20027 13923
rect 20361 13889 20395 13923
rect 20453 13889 20487 13923
rect 20729 13889 20763 13923
rect 21005 13889 21039 13923
rect 21557 13889 21591 13923
rect 24961 13889 24995 13923
rect 25421 13889 25455 13923
rect 25513 13889 25547 13923
rect 25697 13889 25731 13923
rect 25789 13889 25823 13923
rect 26065 13889 26099 13923
rect 26249 13889 26283 13923
rect 26341 13889 26375 13923
rect 26709 13889 26743 13923
rect 27169 13889 27203 13923
rect 27445 13889 27479 13923
rect 27629 13889 27663 13923
rect 27721 13889 27755 13923
rect 27905 13889 27939 13923
rect 29469 13889 29503 13923
rect 31493 13889 31527 13923
rect 31585 13889 31619 13923
rect 32321 13889 32355 13923
rect 33057 13889 33091 13923
rect 4629 13821 4663 13855
rect 5825 13821 5859 13855
rect 6377 13821 6411 13855
rect 12817 13821 12851 13855
rect 14105 13821 14139 13855
rect 15761 13821 15795 13855
rect 19533 13821 19567 13855
rect 19625 13821 19659 13855
rect 20177 13821 20211 13855
rect 20637 13821 20671 13855
rect 20821 13821 20855 13855
rect 21281 13821 21315 13855
rect 21465 13821 21499 13855
rect 25881 13821 25915 13855
rect 27813 13821 27847 13855
rect 32229 13821 32263 13855
rect 5181 13753 5215 13787
rect 5273 13753 5307 13787
rect 6101 13753 6135 13787
rect 15209 13753 15243 13787
rect 15577 13753 15611 13787
rect 18429 13753 18463 13787
rect 26157 13753 26191 13787
rect 27261 13753 27295 13787
rect 27353 13753 27387 13787
rect 31861 13753 31895 13787
rect 4905 13685 4939 13719
rect 8769 13685 8803 13719
rect 14565 13685 14599 13719
rect 21189 13685 21223 13719
rect 22937 13685 22971 13719
rect 26985 13685 27019 13719
rect 29726 13685 29760 13719
rect 31217 13685 31251 13719
rect 31493 13685 31527 13719
rect 32597 13685 32631 13719
rect 33314 13685 33348 13719
rect 3157 13481 3191 13515
rect 12173 13481 12207 13515
rect 13553 13481 13587 13515
rect 13829 13481 13863 13515
rect 15761 13481 15795 13515
rect 18705 13481 18739 13515
rect 18981 13481 19015 13515
rect 19625 13481 19659 13515
rect 19717 13481 19751 13515
rect 21833 13481 21867 13515
rect 22661 13481 22695 13515
rect 26341 13481 26375 13515
rect 28273 13481 28307 13515
rect 30389 13481 30423 13515
rect 30573 13481 30607 13515
rect 34161 13481 34195 13515
rect 15117 13413 15151 13447
rect 17601 13413 17635 13447
rect 20821 13413 20855 13447
rect 25697 13413 25731 13447
rect 26249 13413 26283 13447
rect 27537 13413 27571 13447
rect 1409 13345 1443 13379
rect 4813 13345 4847 13379
rect 5089 13345 5123 13379
rect 7297 13345 7331 13379
rect 8769 13345 8803 13379
rect 10149 13345 10183 13379
rect 15393 13345 15427 13379
rect 16221 13345 16255 13379
rect 19533 13345 19567 13379
rect 21373 13345 21407 13379
rect 23305 13345 23339 13379
rect 27261 13345 27295 13379
rect 27905 13345 27939 13379
rect 32137 13345 32171 13379
rect 32597 13345 32631 13379
rect 4721 13277 4755 13311
rect 7021 13277 7055 13311
rect 9137 13277 9171 13311
rect 9321 13277 9355 13311
rect 10425 13277 10459 13311
rect 12449 13277 12483 13311
rect 14197 13277 14231 13311
rect 14381 13277 14415 13311
rect 16313 13277 16347 13311
rect 16681 13277 16715 13311
rect 16957 13277 16991 13311
rect 17233 13277 17267 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 18889 13277 18923 13311
rect 19073 13277 19107 13311
rect 19257 13277 19291 13311
rect 20453 13277 20487 13311
rect 20729 13277 20763 13311
rect 21189 13277 21223 13311
rect 22937 13277 22971 13311
rect 23397 13277 23431 13311
rect 24685 13277 24719 13311
rect 24961 13277 24995 13311
rect 25237 13277 25271 13311
rect 25513 13277 25547 13311
rect 25789 13277 25823 13311
rect 26065 13277 26099 13311
rect 26525 13277 26559 13311
rect 27169 13277 27203 13311
rect 27997 13277 28031 13311
rect 30481 13277 30515 13311
rect 32045 13277 32079 13311
rect 32505 13277 32539 13311
rect 32689 13277 32723 13311
rect 32965 13277 32999 13311
rect 34069 13277 34103 13311
rect 34529 13277 34563 13311
rect 1685 13209 1719 13243
rect 9045 13209 9079 13243
rect 10701 13209 10735 13243
rect 12357 13209 12391 13243
rect 14565 13209 14599 13243
rect 23121 13209 23155 13243
rect 33609 13209 33643 13243
rect 33885 13209 33919 13243
rect 3525 13141 3559 13175
rect 12725 13141 12759 13175
rect 13185 13141 13219 13175
rect 17417 13141 17451 13175
rect 17877 13141 17911 13175
rect 18153 13141 18187 13175
rect 19349 13141 19383 13175
rect 19993 13141 20027 13175
rect 20269 13141 20303 13175
rect 20637 13141 20671 13175
rect 21281 13141 21315 13175
rect 23029 13141 23063 13175
rect 24869 13141 24903 13175
rect 25145 13141 25179 13175
rect 25421 13141 25455 13175
rect 25973 13141 26007 13175
rect 32413 13141 32447 13175
rect 34437 13141 34471 13175
rect 1593 12937 1627 12971
rect 2329 12937 2363 12971
rect 4537 12937 4571 12971
rect 5657 12937 5691 12971
rect 10333 12937 10367 12971
rect 12449 12937 12483 12971
rect 13829 12937 13863 12971
rect 14105 12937 14139 12971
rect 17417 12937 17451 12971
rect 18705 12937 18739 12971
rect 19165 12937 19199 12971
rect 19549 12937 19583 12971
rect 19717 12937 19751 12971
rect 23857 12937 23891 12971
rect 24501 12937 24535 12971
rect 24777 12937 24811 12971
rect 25145 12937 25179 12971
rect 25697 12937 25731 12971
rect 25973 12937 26007 12971
rect 27813 12937 27847 12971
rect 28549 12937 28583 12971
rect 32965 12937 32999 12971
rect 3065 12869 3099 12903
rect 4721 12869 4755 12903
rect 5089 12869 5123 12903
rect 5457 12869 5491 12903
rect 19349 12869 19383 12903
rect 19993 12869 20027 12903
rect 20545 12869 20579 12903
rect 26801 12869 26835 12903
rect 27077 12869 27111 12903
rect 33333 12869 33367 12903
rect 1409 12801 1443 12835
rect 2237 12801 2271 12835
rect 4813 12801 4847 12835
rect 8033 12801 8067 12835
rect 12633 12801 12667 12835
rect 12817 12801 12851 12835
rect 14013 12801 14047 12835
rect 14289 12801 14323 12835
rect 14473 12801 14507 12835
rect 14565 12801 14599 12835
rect 14749 12801 14783 12835
rect 14933 12801 14967 12835
rect 15117 12801 15151 12835
rect 15945 12801 15979 12835
rect 16129 12801 16163 12835
rect 16313 12801 16347 12835
rect 16773 12801 16807 12835
rect 16957 12801 16991 12835
rect 23397 12801 23431 12835
rect 24593 12801 24627 12835
rect 24869 12801 24903 12835
rect 24961 12801 24995 12835
rect 25605 12801 25639 12835
rect 25881 12801 25915 12835
rect 26157 12801 26191 12835
rect 26433 12801 26467 12835
rect 26617 12801 26651 12835
rect 26985 12801 27019 12835
rect 27261 12801 27295 12835
rect 27537 12801 27571 12835
rect 27629 12801 27663 12835
rect 28641 12801 28675 12835
rect 33057 12801 33091 12835
rect 2789 12733 2823 12767
rect 14841 12733 14875 12767
rect 20821 12733 20855 12767
rect 23305 12733 23339 12767
rect 24133 12733 24167 12767
rect 25053 12733 25087 12767
rect 27445 12733 27479 12767
rect 27813 12733 27847 12767
rect 28917 12733 28951 12767
rect 8861 12665 8895 12699
rect 13461 12665 13495 12699
rect 15669 12665 15703 12699
rect 17877 12665 17911 12699
rect 21189 12665 21223 12699
rect 23765 12665 23799 12699
rect 25421 12665 25455 12699
rect 2145 12597 2179 12631
rect 5641 12597 5675 12631
rect 5825 12597 5859 12631
rect 8125 12597 8159 12631
rect 8585 12597 8619 12631
rect 9229 12597 9263 12631
rect 12633 12597 12667 12631
rect 15301 12597 15335 12631
rect 16221 12597 16255 12631
rect 16957 12597 16991 12631
rect 18337 12597 18371 12631
rect 19533 12597 19567 12631
rect 24225 12597 24259 12631
rect 24317 12597 24351 12631
rect 25145 12597 25179 12631
rect 30389 12597 30423 12631
rect 34805 12597 34839 12631
rect 4629 12393 4663 12427
rect 17877 12393 17911 12427
rect 19533 12393 19567 12427
rect 19993 12393 20027 12427
rect 20729 12393 20763 12427
rect 25237 12393 25271 12427
rect 29745 12393 29779 12427
rect 30205 12393 30239 12427
rect 31677 12393 31711 12427
rect 16129 12325 16163 12359
rect 17509 12325 17543 12359
rect 21005 12325 21039 12359
rect 25329 12325 25363 12359
rect 5825 12257 5859 12291
rect 6285 12257 6319 12291
rect 7297 12257 7331 12291
rect 8769 12257 8803 12291
rect 10977 12257 11011 12291
rect 20085 12257 20119 12291
rect 22017 12257 22051 12291
rect 22293 12257 22327 12291
rect 31033 12257 31067 12291
rect 31401 12257 31435 12291
rect 34069 12257 34103 12291
rect 5917 12189 5951 12223
rect 6745 12189 6779 12223
rect 7021 12189 7055 12223
rect 10425 12189 10459 12223
rect 12449 12189 12483 12223
rect 12817 12189 12851 12223
rect 14565 12189 14599 12223
rect 14841 12189 14875 12223
rect 16313 12189 16347 12223
rect 16773 12189 16807 12223
rect 16957 12189 16991 12223
rect 17233 12189 17267 12223
rect 17325 12189 17359 12223
rect 18153 12189 18187 12223
rect 18245 12189 18279 12223
rect 18705 12189 18739 12223
rect 20223 12189 20257 12223
rect 20361 12189 20395 12223
rect 20453 12189 20487 12223
rect 20545 12189 20579 12223
rect 21189 12189 21223 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 21925 12189 21959 12223
rect 24041 12189 24075 12223
rect 24501 12189 24535 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 25513 12189 25547 12223
rect 27813 12189 27847 12223
rect 28365 12189 28399 12223
rect 29653 12189 29687 12223
rect 31125 12189 31159 12223
rect 31217 12189 31251 12223
rect 34437 12189 34471 12223
rect 16497 12121 16531 12155
rect 17141 12121 17175 12155
rect 17509 12121 17543 12155
rect 6929 12053 6963 12087
rect 9137 12053 9171 12087
rect 16405 12053 16439 12087
rect 16681 12053 16715 12087
rect 17969 12053 18003 12087
rect 18429 12053 18463 12087
rect 18521 12053 18555 12087
rect 24225 12053 24259 12087
rect 24685 12053 24719 12087
rect 24961 12053 24995 12087
rect 27905 12053 27939 12087
rect 28641 12053 28675 12087
rect 31401 12053 31435 12087
rect 4629 11849 4663 11883
rect 5181 11849 5215 11883
rect 8401 11849 8435 11883
rect 12541 11849 12575 11883
rect 13553 11849 13587 11883
rect 13921 11849 13955 11883
rect 14289 11849 14323 11883
rect 15209 11849 15243 11883
rect 15577 11849 15611 11883
rect 19441 11849 19475 11883
rect 23673 11849 23707 11883
rect 23857 11849 23891 11883
rect 24501 11849 24535 11883
rect 24593 11849 24627 11883
rect 32413 11849 32447 11883
rect 3157 11781 3191 11815
rect 4813 11781 4847 11815
rect 5549 11781 5583 11815
rect 8769 11781 8803 11815
rect 10425 11781 10459 11815
rect 12725 11781 12759 11815
rect 14841 11781 14875 11815
rect 23489 11781 23523 11815
rect 24685 11781 24719 11815
rect 26341 11781 26375 11815
rect 28733 11781 28767 11815
rect 34437 11781 34471 11815
rect 2145 11713 2179 11747
rect 4905 11713 4939 11747
rect 6009 11713 6043 11747
rect 6377 11713 6411 11747
rect 8217 11713 8251 11747
rect 8493 11713 8527 11747
rect 10517 11713 10551 11747
rect 10701 11713 10735 11747
rect 12817 11713 12851 11747
rect 13001 11713 13035 11747
rect 14473 11713 14507 11747
rect 14657 11713 14691 11747
rect 15761 11713 15795 11747
rect 15853 11713 15887 11747
rect 16037 11713 16071 11747
rect 16129 11713 16163 11747
rect 16865 11713 16899 11747
rect 17049 11713 17083 11747
rect 17141 11713 17175 11747
rect 17325 11713 17359 11747
rect 17417 11713 17451 11747
rect 18337 11713 18371 11747
rect 18705 11713 18739 11747
rect 18889 11713 18923 11747
rect 18981 11713 19015 11747
rect 19073 11713 19107 11747
rect 19257 11713 19291 11747
rect 19717 11713 19751 11747
rect 19809 11713 19843 11747
rect 19947 11713 19981 11747
rect 20085 11713 20119 11747
rect 20177 11713 20211 11747
rect 20361 11713 20395 11747
rect 20637 11713 20671 11747
rect 21005 11713 21039 11747
rect 21189 11713 21223 11747
rect 21465 11713 21499 11747
rect 24041 11713 24075 11747
rect 24133 11713 24167 11747
rect 24317 11713 24351 11747
rect 24593 11713 24627 11747
rect 24869 11713 24903 11747
rect 25329 11713 25363 11747
rect 25513 11713 25547 11747
rect 25789 11713 25823 11747
rect 26249 11713 26283 11747
rect 26433 11713 26467 11747
rect 26709 11713 26743 11747
rect 26985 11713 27019 11747
rect 30849 11713 30883 11747
rect 31493 11713 31527 11747
rect 31585 11713 31619 11747
rect 31769 11713 31803 11747
rect 32505 11713 32539 11747
rect 34529 11713 34563 11747
rect 34897 11713 34931 11747
rect 2881 11645 2915 11679
rect 8125 11645 8159 11679
rect 10241 11645 10275 11679
rect 11253 11645 11287 11679
rect 18153 11645 18187 11679
rect 18245 11645 18279 11679
rect 18429 11645 18463 11679
rect 18613 11645 18647 11679
rect 21281 11645 21315 11679
rect 25421 11645 25455 11679
rect 25697 11645 25731 11679
rect 28825 11645 28859 11679
rect 29101 11645 29135 11679
rect 30573 11645 30607 11679
rect 30941 11645 30975 11679
rect 31309 11645 31343 11679
rect 32781 11645 32815 11679
rect 2697 11577 2731 11611
rect 19533 11577 19567 11611
rect 21189 11577 21223 11611
rect 25145 11577 25179 11611
rect 31677 11577 31711 11611
rect 2237 11509 2271 11543
rect 6193 11509 6227 11543
rect 12173 11509 12207 11543
rect 16313 11509 16347 11543
rect 21649 11509 21683 11543
rect 23673 11509 23707 11543
rect 26157 11509 26191 11543
rect 31217 11509 31251 11543
rect 34253 11509 34287 11543
rect 3157 11305 3191 11339
rect 15393 11305 15427 11339
rect 15761 11305 15795 11339
rect 16129 11305 16163 11339
rect 17141 11305 17175 11339
rect 17785 11305 17819 11339
rect 18153 11305 18187 11339
rect 18613 11305 18647 11339
rect 20913 11305 20947 11339
rect 21281 11305 21315 11339
rect 25237 11305 25271 11339
rect 29837 11305 29871 11339
rect 30113 11305 30147 11339
rect 30757 11305 30791 11339
rect 31217 11305 31251 11339
rect 31861 11305 31895 11339
rect 3525 11237 3559 11271
rect 4537 11237 4571 11271
rect 17555 11237 17589 11271
rect 23857 11237 23891 11271
rect 24225 11237 24259 11271
rect 26065 11237 26099 11271
rect 32597 11237 32631 11271
rect 6837 11169 6871 11203
rect 8309 11169 8343 11203
rect 11069 11169 11103 11203
rect 27077 11169 27111 11203
rect 28549 11169 28583 11203
rect 30849 11169 30883 11203
rect 31493 11169 31527 11203
rect 33057 11169 33091 11203
rect 34529 11169 34563 11203
rect 1409 11101 1443 11135
rect 4169 11101 4203 11135
rect 6561 11101 6595 11135
rect 8585 11101 8619 11135
rect 8953 11101 8987 11135
rect 9781 11101 9815 11135
rect 17417 11101 17451 11135
rect 17693 11101 17727 11135
rect 17969 11101 18003 11135
rect 18061 11101 18095 11135
rect 18429 11101 18463 11135
rect 18889 11101 18923 11135
rect 18981 11101 19015 11135
rect 19257 11101 19291 11135
rect 19809 11101 19843 11135
rect 19993 11101 20027 11135
rect 20361 11101 20395 11135
rect 20821 11101 20855 11135
rect 21097 11101 21131 11135
rect 21649 11101 21683 11135
rect 22753 11101 22787 11135
rect 23213 11101 23247 11135
rect 23673 11101 23707 11135
rect 26617 11101 26651 11135
rect 26801 11101 26835 11135
rect 30205 11101 30239 11135
rect 30757 11101 30791 11135
rect 31033 11101 31067 11135
rect 31585 11101 31619 11135
rect 32781 11101 32815 11135
rect 34713 11101 34747 11135
rect 1685 11033 1719 11067
rect 4077 11033 4111 11067
rect 8493 11033 8527 11067
rect 16957 11033 16991 11067
rect 17157 11033 17191 11067
rect 20637 11033 20671 11067
rect 22293 11033 22327 11067
rect 34805 11033 34839 11067
rect 10701 10965 10735 10999
rect 17325 10965 17359 10999
rect 17969 10965 18003 10999
rect 18705 10965 18739 10999
rect 21741 10965 21775 10999
rect 28825 10965 28859 10999
rect 1593 10761 1627 10795
rect 4629 10761 4663 10795
rect 5733 10761 5767 10795
rect 8309 10761 8343 10795
rect 21097 10761 21131 10795
rect 21931 10761 21965 10795
rect 23489 10761 23523 10795
rect 31769 10761 31803 10795
rect 34529 10761 34563 10795
rect 8677 10693 8711 10727
rect 9137 10693 9171 10727
rect 21005 10693 21039 10727
rect 21281 10693 21315 10727
rect 21833 10693 21867 10727
rect 22937 10693 22971 10727
rect 1409 10625 1443 10659
rect 5549 10625 5583 10659
rect 17785 10625 17819 10659
rect 17969 10625 18003 10659
rect 22017 10625 22051 10659
rect 22109 10625 22143 10659
rect 22293 10625 22327 10659
rect 22569 10625 22603 10659
rect 22661 10625 22695 10659
rect 23489 10625 23523 10659
rect 23949 10625 23983 10659
rect 24225 10625 24259 10659
rect 30849 10625 30883 10659
rect 31309 10625 31343 10659
rect 31493 10625 31527 10659
rect 2881 10557 2915 10591
rect 3157 10557 3191 10591
rect 23213 10557 23247 10591
rect 30941 10557 30975 10591
rect 31401 10557 31435 10591
rect 17969 10489 18003 10523
rect 31217 10489 31251 10523
rect 4905 10421 4939 10455
rect 21557 10421 21591 10455
rect 3157 10217 3191 10251
rect 16037 10217 16071 10251
rect 17233 10217 17267 10251
rect 22293 10217 22327 10251
rect 3525 10149 3559 10183
rect 17049 10149 17083 10183
rect 20729 10149 20763 10183
rect 31493 10149 31527 10183
rect 1409 10081 1443 10115
rect 16129 10081 16163 10115
rect 16313 10081 16347 10115
rect 20453 10081 20487 10115
rect 21649 10081 21683 10115
rect 21833 10081 21867 10115
rect 34069 10081 34103 10115
rect 15669 10013 15703 10047
rect 16221 10013 16255 10047
rect 16589 10013 16623 10047
rect 16681 10013 16715 10047
rect 16773 10013 16807 10047
rect 16957 10013 16991 10047
rect 17601 10013 17635 10047
rect 17785 10013 17819 10047
rect 18153 10013 18187 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 18555 10013 18589 10047
rect 20361 10013 20395 10047
rect 21925 10013 21959 10047
rect 26065 10013 26099 10047
rect 28089 10013 28123 10047
rect 31309 10013 31343 10047
rect 32045 10013 32079 10047
rect 32689 10013 32723 10047
rect 34437 10013 34471 10047
rect 1685 9945 1719 9979
rect 17217 9945 17251 9979
rect 17417 9945 17451 9979
rect 18797 9945 18831 9979
rect 32597 9945 32631 9979
rect 15761 9877 15795 9911
rect 17693 9877 17727 9911
rect 27353 9877 27387 9911
rect 32229 9877 32263 9911
rect 32781 9877 32815 9911
rect 17509 9673 17543 9707
rect 18153 9673 18187 9707
rect 2421 9605 2455 9639
rect 16865 9605 16899 9639
rect 32413 9605 32447 9639
rect 2329 9537 2363 9571
rect 2789 9537 2823 9571
rect 17233 9537 17267 9571
rect 17325 9537 17359 9571
rect 17863 9537 17897 9571
rect 18429 9537 18463 9571
rect 18613 9537 18647 9571
rect 18705 9537 18739 9571
rect 18889 9537 18923 9571
rect 19441 9537 19475 9571
rect 27169 9537 27203 9571
rect 34161 9537 34195 9571
rect 34437 9537 34471 9571
rect 17693 9469 17727 9503
rect 18245 9469 18279 9503
rect 27445 9469 27479 9503
rect 31953 9469 31987 9503
rect 32137 9469 32171 9503
rect 16957 9333 16991 9367
rect 33885 9333 33919 9367
rect 34069 9333 34103 9367
rect 1593 9129 1627 9163
rect 17693 9129 17727 9163
rect 19533 9129 19567 9163
rect 32045 9129 32079 9163
rect 32137 8993 32171 9027
rect 1409 8925 1443 8959
rect 17509 8925 17543 8959
rect 17693 8925 17727 8959
rect 19349 8925 19383 8959
rect 19533 8925 19567 8959
rect 32413 8857 32447 8891
rect 33885 8789 33919 8823
rect 34069 7905 34103 7939
rect 34345 7837 34379 7871
rect 1409 6749 1443 6783
rect 1593 6613 1627 6647
rect 33333 5661 33367 5695
rect 34345 5593 34379 5627
rect 1593 4777 1627 4811
rect 1409 4573 1443 4607
rect 33333 3485 33367 3519
rect 34345 3417 34379 3451
rect 1593 2601 1627 2635
rect 27353 2601 27387 2635
rect 9597 2465 9631 2499
rect 1409 2397 1443 2431
rect 9137 2397 9171 2431
rect 27537 2397 27571 2431
<< metal1 >>
rect 1104 36474 35248 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 35248 36474
rect 1104 36400 35248 36422
rect 934 36116 940 36168
rect 992 36156 998 36168
rect 1397 36159 1455 36165
rect 1397 36156 1409 36159
rect 992 36128 1409 36156
rect 992 36116 998 36128
rect 1397 36125 1409 36128
rect 1443 36125 1455 36159
rect 1397 36119 1455 36125
rect 33321 36159 33379 36165
rect 33321 36125 33333 36159
rect 33367 36156 33379 36159
rect 33870 36156 33876 36168
rect 33367 36128 33876 36156
rect 33367 36125 33379 36128
rect 33321 36119 33379 36125
rect 33870 36116 33876 36128
rect 33928 36116 33934 36168
rect 34330 36048 34336 36100
rect 34388 36048 34394 36100
rect 1578 35980 1584 36032
rect 1636 35980 1642 36032
rect 1104 35930 35236 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 35236 35930
rect 1104 35856 35236 35878
rect 1104 35386 35248 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 35248 35386
rect 1104 35312 35248 35334
rect 934 35028 940 35080
rect 992 35068 998 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 992 35040 1409 35068
rect 992 35028 998 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 2866 34932 2872 34944
rect 1627 34904 2872 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 2866 34892 2872 34904
rect 2924 34892 2930 34944
rect 1104 34842 35236 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 35236 34842
rect 1104 34768 35236 34790
rect 1104 34298 35248 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 35248 34298
rect 1104 34224 35248 34246
rect 34057 34051 34115 34057
rect 34057 34017 34069 34051
rect 34103 34048 34115 34051
rect 34103 34020 34652 34048
rect 34103 34017 34115 34020
rect 34057 34011 34115 34017
rect 34517 33983 34575 33989
rect 34517 33949 34529 33983
rect 34563 33949 34575 33983
rect 34517 33943 34575 33949
rect 34532 33844 34560 33943
rect 34624 33924 34652 34020
rect 34606 33872 34612 33924
rect 34664 33872 34670 33924
rect 34698 33844 34704 33856
rect 34532 33816 34704 33844
rect 34698 33804 34704 33816
rect 34756 33804 34762 33856
rect 1104 33754 35236 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 35236 33754
rect 1104 33680 35236 33702
rect 1104 33210 35248 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 35248 33210
rect 1104 33136 35248 33158
rect 934 32852 940 32904
rect 992 32892 998 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 992 32864 1409 32892
rect 992 32852 998 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1578 32716 1584 32768
rect 1636 32716 1642 32768
rect 1104 32666 35236 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 35236 32666
rect 1104 32592 35236 32614
rect 1104 32122 35248 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 35248 32122
rect 1104 32048 35248 32070
rect 34057 31875 34115 31881
rect 34057 31841 34069 31875
rect 34103 31841 34115 31875
rect 34057 31835 34115 31841
rect 34072 31680 34100 31835
rect 34514 31764 34520 31816
rect 34572 31764 34578 31816
rect 34054 31628 34060 31680
rect 34112 31628 34118 31680
rect 1104 31578 35236 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 35236 31578
rect 1104 31504 35236 31526
rect 1104 31034 35248 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 35248 31034
rect 1104 30960 35248 30982
rect 1394 30676 1400 30728
rect 1452 30676 1458 30728
rect 32861 30719 32919 30725
rect 32861 30685 32873 30719
rect 32907 30716 32919 30719
rect 32907 30688 32941 30716
rect 32907 30685 32919 30688
rect 32861 30679 32919 30685
rect 32769 30651 32827 30657
rect 32769 30617 32781 30651
rect 32815 30648 32827 30651
rect 32876 30648 32904 30679
rect 32815 30620 34468 30648
rect 32815 30617 32827 30620
rect 32769 30611 32827 30617
rect 34440 30592 34468 30620
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 3694 30580 3700 30592
rect 1627 30552 3700 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 3694 30540 3700 30552
rect 3752 30540 3758 30592
rect 32953 30583 33011 30589
rect 32953 30549 32965 30583
rect 32999 30580 33011 30583
rect 33134 30580 33140 30592
rect 32999 30552 33140 30580
rect 32999 30549 33011 30552
rect 32953 30543 33011 30549
rect 33134 30540 33140 30552
rect 33192 30540 33198 30592
rect 34422 30540 34428 30592
rect 34480 30540 34486 30592
rect 1104 30490 35236 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 35236 30490
rect 1104 30416 35236 30438
rect 29270 30268 29276 30320
rect 29328 30268 29334 30320
rect 33134 30268 33140 30320
rect 33192 30268 33198 30320
rect 30929 30243 30987 30249
rect 30929 30240 30941 30243
rect 30300 30212 30941 30240
rect 28537 30175 28595 30181
rect 28537 30141 28549 30175
rect 28583 30141 28595 30175
rect 28537 30135 28595 30141
rect 28445 30039 28503 30045
rect 28445 30005 28457 30039
rect 28491 30036 28503 30039
rect 28552 30036 28580 30135
rect 28810 30132 28816 30184
rect 28868 30132 28874 30184
rect 30300 30181 30328 30212
rect 30929 30209 30941 30212
rect 30975 30209 30987 30243
rect 30929 30203 30987 30209
rect 31846 30200 31852 30252
rect 31904 30240 31910 30252
rect 32125 30243 32183 30249
rect 32125 30240 32137 30243
rect 31904 30212 32137 30240
rect 31904 30200 31910 30212
rect 32125 30209 32137 30212
rect 32171 30209 32183 30243
rect 32125 30203 32183 30209
rect 34333 30243 34391 30249
rect 34333 30209 34345 30243
rect 34379 30240 34391 30243
rect 34379 30212 34468 30240
rect 34379 30209 34391 30212
rect 34333 30203 34391 30209
rect 30285 30175 30343 30181
rect 30285 30141 30297 30175
rect 30331 30141 30343 30175
rect 30285 30135 30343 30141
rect 31018 30132 31024 30184
rect 31076 30132 31082 30184
rect 32401 30175 32459 30181
rect 32401 30172 32413 30175
rect 32232 30144 32413 30172
rect 31297 30107 31355 30113
rect 31297 30073 31309 30107
rect 31343 30104 31355 30107
rect 32232 30104 32260 30144
rect 32401 30141 32413 30144
rect 32447 30141 32459 30175
rect 32401 30135 32459 30141
rect 31343 30076 32260 30104
rect 31343 30073 31355 30076
rect 31297 30067 31355 30073
rect 33870 30064 33876 30116
rect 33928 30064 33934 30116
rect 34440 30048 34468 30212
rect 29822 30036 29828 30048
rect 28491 30008 29828 30036
rect 28491 30005 28503 30008
rect 28445 29999 28503 30005
rect 29822 29996 29828 30008
rect 29880 30036 29886 30048
rect 31846 30036 31852 30048
rect 29880 30008 31852 30036
rect 29880 29996 29886 30008
rect 31846 29996 31852 30008
rect 31904 29996 31910 30048
rect 34238 29996 34244 30048
rect 34296 29996 34302 30048
rect 34422 29996 34428 30048
rect 34480 30036 34486 30048
rect 34609 30039 34667 30045
rect 34609 30036 34621 30039
rect 34480 30008 34621 30036
rect 34480 29996 34486 30008
rect 34609 30005 34621 30008
rect 34655 30005 34667 30039
rect 34609 29999 34667 30005
rect 1104 29946 35248 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 35248 29946
rect 1104 29872 35248 29894
rect 26513 29835 26571 29841
rect 26513 29801 26525 29835
rect 26559 29832 26571 29835
rect 28810 29832 28816 29844
rect 26559 29804 28816 29832
rect 26559 29801 26571 29804
rect 26513 29795 26571 29801
rect 28810 29792 28816 29804
rect 28868 29792 28874 29844
rect 29270 29792 29276 29844
rect 29328 29792 29334 29844
rect 34514 29792 34520 29844
rect 34572 29792 34578 29844
rect 25409 29767 25467 29773
rect 25409 29733 25421 29767
rect 25455 29764 25467 29767
rect 34238 29764 34244 29776
rect 25455 29736 27844 29764
rect 25455 29733 25467 29736
rect 25409 29727 25467 29733
rect 25130 29656 25136 29708
rect 25188 29656 25194 29708
rect 27816 29705 27844 29736
rect 34164 29736 34244 29764
rect 27801 29699 27859 29705
rect 27801 29665 27813 29699
rect 27847 29665 27859 29699
rect 27801 29659 27859 29665
rect 29549 29699 29607 29705
rect 29549 29665 29561 29699
rect 29595 29696 29607 29699
rect 29822 29696 29828 29708
rect 29595 29668 29828 29696
rect 29595 29665 29607 29668
rect 29549 29659 29607 29665
rect 29822 29656 29828 29668
rect 29880 29656 29886 29708
rect 31297 29699 31355 29705
rect 31297 29665 31309 29699
rect 31343 29696 31355 29699
rect 31343 29668 31754 29696
rect 31343 29665 31355 29668
rect 31297 29659 31355 29665
rect 31726 29640 31754 29668
rect 32214 29656 32220 29708
rect 32272 29656 32278 29708
rect 24029 29631 24087 29637
rect 24029 29628 24041 29631
rect 23400 29600 24041 29628
rect 23400 29504 23428 29600
rect 24029 29597 24041 29600
rect 24075 29597 24087 29631
rect 24029 29591 24087 29597
rect 24213 29631 24271 29637
rect 24213 29597 24225 29631
rect 24259 29628 24271 29631
rect 24259 29600 24440 29628
rect 24259 29597 24271 29600
rect 24213 29591 24271 29597
rect 24412 29504 24440 29600
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 25041 29631 25099 29637
rect 25041 29628 25053 29631
rect 24912 29600 25053 29628
rect 24912 29588 24918 29600
rect 25041 29597 25053 29600
rect 25087 29597 25099 29631
rect 25041 29591 25099 29597
rect 26145 29631 26203 29637
rect 26145 29597 26157 29631
rect 26191 29597 26203 29631
rect 26145 29591 26203 29597
rect 26237 29631 26295 29637
rect 26237 29597 26249 29631
rect 26283 29597 26295 29631
rect 26237 29591 26295 29597
rect 26329 29631 26387 29637
rect 26329 29597 26341 29631
rect 26375 29628 26387 29631
rect 26970 29628 26976 29640
rect 26375 29600 26976 29628
rect 26375 29597 26387 29600
rect 26329 29591 26387 29597
rect 24670 29520 24676 29572
rect 24728 29560 24734 29572
rect 26160 29560 26188 29591
rect 24728 29532 26188 29560
rect 26252 29560 26280 29591
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 27893 29631 27951 29637
rect 27893 29597 27905 29631
rect 27939 29628 27951 29631
rect 28350 29628 28356 29640
rect 27939 29600 28356 29628
rect 27939 29597 27951 29600
rect 27893 29591 27951 29597
rect 28350 29588 28356 29600
rect 28408 29588 28414 29640
rect 29178 29588 29184 29640
rect 29236 29588 29242 29640
rect 31662 29588 31668 29640
rect 31720 29628 31754 29640
rect 32125 29631 32183 29637
rect 32125 29628 32137 29631
rect 31720 29600 32137 29628
rect 31720 29588 31726 29600
rect 32125 29597 32137 29600
rect 32171 29597 32183 29631
rect 32582 29628 32588 29640
rect 32125 29591 32183 29597
rect 32416 29600 32588 29628
rect 27062 29560 27068 29572
rect 26252 29532 27068 29560
rect 24728 29520 24734 29532
rect 27062 29520 27068 29532
rect 27120 29520 27126 29572
rect 29825 29563 29883 29569
rect 29825 29560 29837 29563
rect 28276 29532 29837 29560
rect 23382 29452 23388 29504
rect 23440 29452 23446 29504
rect 24213 29495 24271 29501
rect 24213 29461 24225 29495
rect 24259 29492 24271 29495
rect 24302 29492 24308 29504
rect 24259 29464 24308 29492
rect 24259 29461 24271 29464
rect 24213 29455 24271 29461
rect 24302 29452 24308 29464
rect 24360 29452 24366 29504
rect 24394 29452 24400 29504
rect 24452 29452 24458 29504
rect 28276 29501 28304 29532
rect 29825 29529 29837 29532
rect 29871 29529 29883 29563
rect 29825 29523 29883 29529
rect 30374 29520 30380 29572
rect 30432 29520 30438 29572
rect 31846 29520 31852 29572
rect 31904 29560 31910 29572
rect 32416 29560 32444 29600
rect 32582 29588 32588 29600
rect 32640 29628 32646 29640
rect 32769 29631 32827 29637
rect 32769 29628 32781 29631
rect 32640 29600 32781 29628
rect 32640 29588 32646 29600
rect 32769 29597 32781 29600
rect 32815 29597 32827 29631
rect 34164 29614 34192 29736
rect 34238 29724 34244 29736
rect 34296 29724 34302 29776
rect 32769 29591 32827 29597
rect 33045 29563 33103 29569
rect 33045 29560 33057 29563
rect 31904 29532 32444 29560
rect 32508 29532 33057 29560
rect 31904 29520 31910 29532
rect 28261 29495 28319 29501
rect 28261 29461 28273 29495
rect 28307 29461 28319 29495
rect 28261 29455 28319 29461
rect 29089 29495 29147 29501
rect 29089 29461 29101 29495
rect 29135 29492 29147 29495
rect 29178 29492 29184 29504
rect 29135 29464 29184 29492
rect 29135 29461 29147 29464
rect 29089 29455 29147 29461
rect 29178 29452 29184 29464
rect 29236 29492 29242 29504
rect 30190 29492 30196 29504
rect 29236 29464 30196 29492
rect 29236 29452 29242 29464
rect 30190 29452 30196 29464
rect 30248 29452 30254 29504
rect 32508 29501 32536 29532
rect 33045 29529 33057 29532
rect 33091 29529 33103 29563
rect 33045 29523 33103 29529
rect 32493 29495 32551 29501
rect 32493 29461 32505 29495
rect 32539 29461 32551 29495
rect 32493 29455 32551 29461
rect 1104 29402 35236 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 35236 29402
rect 1104 29328 35236 29350
rect 23293 29291 23351 29297
rect 23293 29257 23305 29291
rect 23339 29288 23351 29291
rect 23658 29288 23664 29300
rect 23339 29260 23664 29288
rect 23339 29257 23351 29260
rect 23293 29251 23351 29257
rect 23658 29248 23664 29260
rect 23716 29248 23722 29300
rect 24854 29288 24860 29300
rect 24136 29260 24860 29288
rect 23934 29220 23940 29232
rect 23216 29192 23940 29220
rect 23216 29161 23244 29192
rect 23934 29180 23940 29192
rect 23992 29180 23998 29232
rect 23201 29155 23259 29161
rect 23201 29121 23213 29155
rect 23247 29121 23259 29155
rect 23201 29115 23259 29121
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23492 29016 23520 29115
rect 23566 29112 23572 29164
rect 23624 29112 23630 29164
rect 23753 29155 23811 29161
rect 23753 29121 23765 29155
rect 23799 29152 23811 29155
rect 24136 29152 24164 29260
rect 24854 29248 24860 29260
rect 24912 29248 24918 29300
rect 25130 29248 25136 29300
rect 25188 29248 25194 29300
rect 29457 29291 29515 29297
rect 29457 29257 29469 29291
rect 29503 29288 29515 29291
rect 29822 29288 29828 29300
rect 29503 29260 29828 29288
rect 29503 29257 29515 29260
rect 29457 29251 29515 29257
rect 29822 29248 29828 29260
rect 29880 29248 29886 29300
rect 30374 29248 30380 29300
rect 30432 29248 30438 29300
rect 32582 29248 32588 29300
rect 32640 29288 32646 29300
rect 32953 29291 33011 29297
rect 32953 29288 32965 29291
rect 32640 29260 32965 29288
rect 32640 29248 32646 29260
rect 32953 29257 32965 29260
rect 32999 29257 33011 29291
rect 32953 29251 33011 29257
rect 24302 29180 24308 29232
rect 24360 29220 24366 29232
rect 24360 29192 24992 29220
rect 24360 29180 24366 29192
rect 23799 29124 24164 29152
rect 24213 29155 24271 29161
rect 23799 29121 23811 29124
rect 23753 29115 23811 29121
rect 24213 29121 24225 29155
rect 24259 29121 24271 29155
rect 24213 29115 24271 29121
rect 23584 29084 23612 29112
rect 24228 29084 24256 29115
rect 24394 29112 24400 29164
rect 24452 29112 24458 29164
rect 24673 29155 24731 29161
rect 24673 29152 24685 29155
rect 24504 29124 24685 29152
rect 24504 29084 24532 29124
rect 24673 29121 24685 29124
rect 24719 29121 24731 29155
rect 24673 29115 24731 29121
rect 24854 29112 24860 29164
rect 24912 29112 24918 29164
rect 24964 29161 24992 29192
rect 25056 29192 25728 29220
rect 25056 29164 25084 29192
rect 24949 29155 25007 29161
rect 24949 29121 24961 29155
rect 24995 29121 25007 29155
rect 24949 29115 25007 29121
rect 25038 29112 25044 29164
rect 25096 29112 25102 29164
rect 25130 29112 25136 29164
rect 25188 29152 25194 29164
rect 25700 29161 25728 29192
rect 25501 29155 25559 29161
rect 25188 29124 25268 29152
rect 25188 29112 25194 29124
rect 23584 29056 24532 29084
rect 24581 29087 24639 29093
rect 24581 29053 24593 29087
rect 24627 29084 24639 29087
rect 25240 29084 25268 29124
rect 25501 29121 25513 29155
rect 25547 29121 25559 29155
rect 25501 29115 25559 29121
rect 25685 29155 25743 29161
rect 25685 29121 25697 29155
rect 25731 29121 25743 29155
rect 30285 29155 30343 29161
rect 30285 29152 30297 29155
rect 25685 29115 25743 29121
rect 30208 29124 30297 29152
rect 24627 29056 25268 29084
rect 24627 29053 24639 29056
rect 24581 29047 24639 29053
rect 24857 29019 24915 29025
rect 24857 29016 24869 29019
rect 23492 28988 24869 29016
rect 24857 28985 24869 28988
rect 24903 29016 24915 29019
rect 25516 29016 25544 29115
rect 24903 28988 25544 29016
rect 25593 29019 25651 29025
rect 24903 28985 24915 28988
rect 24857 28979 24915 28985
rect 25593 28985 25605 29019
rect 25639 29016 25651 29019
rect 26970 29016 26976 29028
rect 25639 28988 26976 29016
rect 25639 28985 25651 28988
rect 25593 28979 25651 28985
rect 26970 28976 26976 28988
rect 27028 28976 27034 29028
rect 30208 28960 30236 29124
rect 30285 29121 30297 29124
rect 30331 29121 30343 29155
rect 32968 29152 32996 29251
rect 34698 29248 34704 29300
rect 34756 29288 34762 29300
rect 34885 29291 34943 29297
rect 34885 29288 34897 29291
rect 34756 29260 34897 29288
rect 34756 29248 34762 29260
rect 34885 29257 34897 29260
rect 34931 29257 34943 29291
rect 34885 29251 34943 29257
rect 34790 29220 34796 29232
rect 34638 29192 34796 29220
rect 34790 29180 34796 29192
rect 34848 29180 34854 29232
rect 33137 29155 33195 29161
rect 33137 29152 33149 29155
rect 32968 29124 33149 29152
rect 30285 29115 30343 29121
rect 33137 29121 33149 29124
rect 33183 29121 33195 29155
rect 33137 29115 33195 29121
rect 23474 28908 23480 28960
rect 23532 28908 23538 28960
rect 26234 28908 26240 28960
rect 26292 28948 26298 28960
rect 27982 28948 27988 28960
rect 26292 28920 27988 28948
rect 26292 28908 26298 28920
rect 27982 28908 27988 28920
rect 28040 28948 28046 28960
rect 28534 28948 28540 28960
rect 28040 28920 28540 28948
rect 28040 28908 28046 28920
rect 28534 28908 28540 28920
rect 28592 28908 28598 28960
rect 30190 28908 30196 28960
rect 30248 28908 30254 28960
rect 33042 28908 33048 28960
rect 33100 28948 33106 28960
rect 33394 28951 33452 28957
rect 33394 28948 33406 28951
rect 33100 28920 33406 28948
rect 33100 28908 33106 28920
rect 33394 28917 33406 28920
rect 33440 28917 33452 28951
rect 33394 28911 33452 28917
rect 1104 28858 35248 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 35248 28858
rect 1104 28784 35248 28806
rect 23934 28704 23940 28756
rect 23992 28744 23998 28756
rect 24029 28747 24087 28753
rect 24029 28744 24041 28747
rect 23992 28716 24041 28744
rect 23992 28704 23998 28716
rect 24029 28713 24041 28716
rect 24075 28713 24087 28747
rect 28350 28744 28356 28756
rect 24029 28707 24087 28713
rect 26896 28716 28356 28744
rect 24762 28636 24768 28688
rect 24820 28636 24826 28688
rect 25915 28679 25973 28685
rect 25915 28645 25927 28679
rect 25961 28676 25973 28679
rect 26510 28676 26516 28688
rect 25961 28648 26516 28676
rect 25961 28645 25973 28648
rect 25915 28639 25973 28645
rect 26510 28636 26516 28648
rect 26568 28636 26574 28688
rect 24486 28608 24492 28620
rect 23860 28580 24492 28608
rect 934 28500 940 28552
rect 992 28540 998 28552
rect 1397 28543 1455 28549
rect 1397 28540 1409 28543
rect 992 28512 1409 28540
rect 992 28500 998 28512
rect 1397 28509 1409 28512
rect 1443 28509 1455 28543
rect 1397 28503 1455 28509
rect 23474 28500 23480 28552
rect 23532 28540 23538 28552
rect 23860 28549 23888 28580
rect 24486 28568 24492 28580
rect 24544 28568 24550 28620
rect 25130 28568 25136 28620
rect 25188 28608 25194 28620
rect 26896 28617 26924 28716
rect 28350 28704 28356 28716
rect 28408 28704 28414 28756
rect 31018 28704 31024 28756
rect 31076 28744 31082 28756
rect 31389 28747 31447 28753
rect 31389 28744 31401 28747
rect 31076 28716 31401 28744
rect 31076 28704 31082 28716
rect 31389 28713 31401 28716
rect 31435 28713 31447 28747
rect 31389 28707 31447 28713
rect 32493 28747 32551 28753
rect 32493 28713 32505 28747
rect 32539 28744 32551 28747
rect 33042 28744 33048 28756
rect 32539 28716 33048 28744
rect 32539 28713 32551 28716
rect 32493 28707 32551 28713
rect 33042 28704 33048 28716
rect 33100 28704 33106 28756
rect 34790 28704 34796 28756
rect 34848 28704 34854 28756
rect 28258 28636 28264 28688
rect 28316 28676 28322 28688
rect 28316 28648 28994 28676
rect 28316 28636 28322 28648
rect 25317 28611 25375 28617
rect 25317 28608 25329 28611
rect 25188 28580 25329 28608
rect 25188 28568 25194 28580
rect 25317 28577 25329 28580
rect 25363 28577 25375 28611
rect 25317 28571 25375 28577
rect 25777 28611 25835 28617
rect 25777 28577 25789 28611
rect 25823 28608 25835 28611
rect 26881 28611 26939 28617
rect 25823 28580 26372 28608
rect 25823 28577 25835 28580
rect 25777 28571 25835 28577
rect 23753 28543 23811 28549
rect 23753 28540 23765 28543
rect 23532 28512 23765 28540
rect 23532 28500 23538 28512
rect 23753 28509 23765 28512
rect 23799 28509 23811 28543
rect 23753 28503 23811 28509
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28509 23903 28543
rect 23845 28503 23903 28509
rect 24121 28543 24179 28549
rect 24121 28509 24133 28543
rect 24167 28509 24179 28543
rect 24121 28503 24179 28509
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28540 24455 28543
rect 24504 28540 24532 28568
rect 26344 28552 26372 28580
rect 26881 28577 26893 28611
rect 26927 28577 26939 28611
rect 26881 28571 26939 28577
rect 26970 28568 26976 28620
rect 27028 28568 27034 28620
rect 27617 28611 27675 28617
rect 27617 28577 27629 28611
rect 27663 28608 27675 28611
rect 28074 28608 28080 28620
rect 27663 28580 28080 28608
rect 27663 28577 27675 28580
rect 27617 28571 27675 28577
rect 28074 28568 28080 28580
rect 28132 28568 28138 28620
rect 24443 28512 24532 28540
rect 24581 28543 24639 28549
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 24581 28509 24593 28543
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 25501 28543 25559 28549
rect 25501 28509 25513 28543
rect 25547 28540 25559 28543
rect 25593 28543 25651 28549
rect 25593 28540 25605 28543
rect 25547 28512 25605 28540
rect 25547 28509 25559 28512
rect 25501 28503 25559 28509
rect 25593 28509 25605 28512
rect 25639 28509 25651 28543
rect 25593 28503 25651 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28540 26111 28543
rect 26234 28540 26240 28552
rect 26099 28512 26240 28540
rect 26099 28509 26111 28512
rect 26053 28503 26111 28509
rect 23658 28432 23664 28484
rect 23716 28432 23722 28484
rect 24136 28472 24164 28503
rect 24489 28475 24547 28481
rect 24489 28472 24501 28475
rect 24136 28444 24501 28472
rect 24489 28441 24501 28444
rect 24535 28441 24547 28475
rect 24489 28435 24547 28441
rect 24596 28472 24624 28503
rect 26234 28500 26240 28512
rect 26292 28500 26298 28552
rect 26326 28500 26332 28552
rect 26384 28500 26390 28552
rect 27062 28500 27068 28552
rect 27120 28540 27126 28552
rect 27341 28543 27399 28549
rect 27341 28540 27353 28543
rect 27120 28512 27353 28540
rect 27120 28500 27126 28512
rect 27341 28509 27353 28512
rect 27387 28540 27399 28543
rect 27709 28543 27767 28549
rect 27709 28540 27721 28543
rect 27387 28512 27721 28540
rect 27387 28509 27399 28512
rect 27341 28503 27399 28509
rect 27709 28509 27721 28512
rect 27755 28509 27767 28543
rect 27893 28543 27951 28549
rect 27893 28540 27905 28543
rect 27709 28503 27767 28509
rect 27816 28512 27905 28540
rect 24765 28475 24823 28481
rect 24765 28472 24777 28475
rect 24596 28444 24777 28472
rect 1578 28364 1584 28416
rect 1636 28364 1642 28416
rect 23566 28364 23572 28416
rect 23624 28364 23630 28416
rect 23676 28404 23704 28432
rect 24596 28404 24624 28444
rect 24765 28441 24777 28444
rect 24811 28472 24823 28475
rect 25038 28472 25044 28484
rect 24811 28444 25044 28472
rect 24811 28441 24823 28444
rect 24765 28435 24823 28441
rect 25038 28432 25044 28444
rect 25096 28472 25102 28484
rect 25406 28472 25412 28484
rect 25096 28444 25412 28472
rect 25096 28432 25102 28444
rect 25406 28432 25412 28444
rect 25464 28432 25470 28484
rect 25685 28475 25743 28481
rect 25685 28441 25697 28475
rect 25731 28472 25743 28475
rect 27249 28475 27307 28481
rect 27249 28472 27261 28475
rect 25731 28444 27261 28472
rect 25731 28441 25743 28444
rect 25685 28435 25743 28441
rect 27249 28441 27261 28444
rect 27295 28441 27307 28475
rect 27816 28472 27844 28512
rect 27893 28509 27905 28512
rect 27939 28509 27951 28543
rect 27893 28503 27951 28509
rect 27982 28500 27988 28552
rect 28040 28500 28046 28552
rect 28166 28500 28172 28552
rect 28224 28500 28230 28552
rect 28261 28543 28319 28549
rect 28261 28509 28273 28543
rect 28307 28509 28319 28543
rect 28629 28543 28687 28549
rect 28629 28540 28641 28543
rect 28261 28503 28319 28509
rect 28460 28512 28641 28540
rect 27249 28435 27307 28441
rect 27724 28444 27844 28472
rect 27724 28416 27752 28444
rect 28074 28432 28080 28484
rect 28132 28472 28138 28484
rect 28276 28472 28304 28503
rect 28353 28475 28411 28481
rect 28353 28472 28365 28475
rect 28132 28444 28365 28472
rect 28132 28432 28138 28444
rect 28353 28441 28365 28444
rect 28399 28441 28411 28475
rect 28353 28435 28411 28441
rect 23676 28376 24624 28404
rect 24854 28364 24860 28416
rect 24912 28404 24918 28416
rect 25225 28407 25283 28413
rect 25225 28404 25237 28407
rect 24912 28376 25237 28404
rect 24912 28364 24918 28376
rect 25225 28373 25237 28376
rect 25271 28373 25283 28407
rect 25225 28367 25283 28373
rect 26234 28364 26240 28416
rect 26292 28404 26298 28416
rect 27157 28407 27215 28413
rect 27157 28404 27169 28407
rect 26292 28376 27169 28404
rect 26292 28364 26298 28376
rect 27157 28373 27169 28376
rect 27203 28373 27215 28407
rect 27157 28367 27215 28373
rect 27706 28364 27712 28416
rect 27764 28404 27770 28416
rect 28460 28404 28488 28512
rect 28629 28509 28641 28512
rect 28675 28509 28687 28543
rect 28629 28503 28687 28509
rect 28534 28432 28540 28484
rect 28592 28432 28598 28484
rect 28966 28472 28994 28648
rect 31662 28636 31668 28688
rect 31720 28636 31726 28688
rect 32214 28636 32220 28688
rect 32272 28676 32278 28688
rect 32769 28679 32827 28685
rect 32769 28676 32781 28679
rect 32272 28648 32781 28676
rect 32272 28636 32278 28648
rect 32769 28645 32781 28648
rect 32815 28645 32827 28679
rect 32769 28639 32827 28645
rect 29365 28611 29423 28617
rect 29365 28577 29377 28611
rect 29411 28608 29423 28611
rect 29549 28611 29607 28617
rect 29549 28608 29561 28611
rect 29411 28580 29561 28608
rect 29411 28577 29423 28580
rect 29365 28571 29423 28577
rect 29549 28577 29561 28580
rect 29595 28608 29607 28611
rect 29822 28608 29828 28620
rect 29595 28580 29828 28608
rect 29595 28577 29607 28580
rect 29549 28571 29607 28577
rect 29822 28568 29828 28580
rect 29880 28568 29886 28620
rect 31297 28611 31355 28617
rect 31297 28577 31309 28611
rect 31343 28577 31355 28611
rect 31297 28571 31355 28577
rect 31312 28540 31340 28571
rect 32306 28568 32312 28620
rect 32364 28568 32370 28620
rect 34054 28568 34060 28620
rect 34112 28568 34118 28620
rect 31573 28543 31631 28549
rect 31573 28540 31585 28543
rect 31312 28512 31585 28540
rect 31573 28509 31585 28512
rect 31619 28509 31631 28543
rect 31573 28503 31631 28509
rect 29825 28475 29883 28481
rect 29825 28472 29837 28475
rect 28966 28444 29837 28472
rect 29825 28441 29837 28444
rect 29871 28441 29883 28475
rect 29825 28435 29883 28441
rect 30282 28432 30288 28484
rect 30340 28432 30346 28484
rect 31588 28472 31616 28503
rect 31754 28500 31760 28552
rect 31812 28500 31818 28552
rect 31849 28543 31907 28549
rect 31849 28509 31861 28543
rect 31895 28540 31907 28543
rect 32030 28540 32036 28552
rect 31895 28512 32036 28540
rect 31895 28509 31907 28512
rect 31849 28503 31907 28509
rect 32030 28500 32036 28512
rect 32088 28500 32094 28552
rect 32217 28543 32275 28549
rect 32217 28509 32229 28543
rect 32263 28509 32275 28543
rect 32217 28503 32275 28509
rect 32677 28543 32735 28549
rect 32677 28509 32689 28543
rect 32723 28509 32735 28543
rect 32861 28543 32919 28549
rect 32861 28540 32873 28543
rect 32677 28503 32735 28509
rect 32784 28512 32873 28540
rect 32232 28472 32260 28503
rect 31588 28444 32260 28472
rect 27764 28376 28488 28404
rect 27764 28364 27770 28376
rect 31754 28364 31760 28416
rect 31812 28404 31818 28416
rect 32692 28404 32720 28503
rect 32784 28416 32812 28512
rect 32861 28509 32873 28512
rect 32907 28509 32919 28543
rect 32861 28503 32919 28509
rect 34514 28500 34520 28552
rect 34572 28500 34578 28552
rect 34701 28543 34759 28549
rect 34701 28509 34713 28543
rect 34747 28509 34759 28543
rect 34701 28503 34759 28509
rect 34716 28472 34744 28503
rect 34440 28444 34744 28472
rect 34440 28416 34468 28444
rect 31812 28376 32720 28404
rect 31812 28364 31818 28376
rect 32766 28364 32772 28416
rect 32824 28364 32830 28416
rect 34422 28364 34428 28416
rect 34480 28364 34486 28416
rect 1104 28314 35236 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 35236 28314
rect 1104 28240 35236 28262
rect 27706 28160 27712 28212
rect 27764 28160 27770 28212
rect 27893 28203 27951 28209
rect 27893 28169 27905 28203
rect 27939 28200 27951 28203
rect 28074 28200 28080 28212
rect 27939 28172 28080 28200
rect 27939 28169 27951 28172
rect 27893 28163 27951 28169
rect 28074 28160 28080 28172
rect 28132 28160 28138 28212
rect 30282 28160 30288 28212
rect 30340 28160 30346 28212
rect 32306 28160 32312 28212
rect 32364 28200 32370 28212
rect 32401 28203 32459 28209
rect 32401 28200 32413 28203
rect 32364 28172 32413 28200
rect 32364 28160 32370 28172
rect 32401 28169 32413 28172
rect 32447 28169 32459 28203
rect 32401 28163 32459 28169
rect 27540 28104 28028 28132
rect 27540 28076 27568 28104
rect 27522 28024 27528 28076
rect 27580 28024 27586 28076
rect 27706 28024 27712 28076
rect 27764 28064 27770 28076
rect 28000 28073 28028 28104
rect 27801 28067 27859 28073
rect 27801 28064 27813 28067
rect 27764 28036 27813 28064
rect 27764 28024 27770 28036
rect 27801 28033 27813 28036
rect 27847 28033 27859 28067
rect 27801 28027 27859 28033
rect 27985 28067 28043 28073
rect 27985 28033 27997 28067
rect 28031 28033 28043 28067
rect 27985 28027 28043 28033
rect 30190 28024 30196 28076
rect 30248 28024 30254 28076
rect 31662 28024 31668 28076
rect 31720 28064 31726 28076
rect 32125 28067 32183 28073
rect 32125 28064 32137 28067
rect 31720 28036 32137 28064
rect 31720 28024 31726 28036
rect 32125 28033 32137 28036
rect 32171 28033 32183 28067
rect 32125 28027 32183 28033
rect 23566 27956 23572 28008
rect 23624 27996 23630 28008
rect 28166 27996 28172 28008
rect 23624 27968 28172 27996
rect 23624 27956 23630 27968
rect 28166 27956 28172 27968
rect 28224 27956 28230 28008
rect 30101 27863 30159 27869
rect 30101 27829 30113 27863
rect 30147 27860 30159 27863
rect 30208 27860 30236 28024
rect 32030 27956 32036 28008
rect 32088 27996 32094 28008
rect 32401 27999 32459 28005
rect 32401 27996 32413 27999
rect 32088 27968 32413 27996
rect 32088 27956 32094 27968
rect 32324 27872 32352 27968
rect 32401 27965 32413 27968
rect 32447 27996 32459 27999
rect 32766 27996 32772 28008
rect 32447 27968 32772 27996
rect 32447 27965 32459 27968
rect 32401 27959 32459 27965
rect 32766 27956 32772 27968
rect 32824 27956 32830 28008
rect 31294 27860 31300 27872
rect 30147 27832 31300 27860
rect 30147 27829 30159 27832
rect 30101 27823 30159 27829
rect 31294 27820 31300 27832
rect 31352 27820 31358 27872
rect 31754 27820 31760 27872
rect 31812 27860 31818 27872
rect 32217 27863 32275 27869
rect 32217 27860 32229 27863
rect 31812 27832 32229 27860
rect 31812 27820 31818 27832
rect 32217 27829 32229 27832
rect 32263 27829 32275 27863
rect 32217 27823 32275 27829
rect 32306 27820 32312 27872
rect 32364 27820 32370 27872
rect 34241 27863 34299 27869
rect 34241 27829 34253 27863
rect 34287 27860 34299 27863
rect 34422 27860 34428 27872
rect 34287 27832 34428 27860
rect 34287 27829 34299 27832
rect 34241 27823 34299 27829
rect 34422 27820 34428 27832
rect 34480 27860 34486 27872
rect 34517 27863 34575 27869
rect 34517 27860 34529 27863
rect 34480 27832 34529 27860
rect 34480 27820 34486 27832
rect 34517 27829 34529 27832
rect 34563 27829 34575 27863
rect 34517 27823 34575 27829
rect 1104 27770 35248 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 35248 27770
rect 1104 27696 35248 27718
rect 19797 27659 19855 27665
rect 19797 27625 19809 27659
rect 19843 27656 19855 27659
rect 21358 27656 21364 27668
rect 19843 27628 21364 27656
rect 19843 27625 19855 27628
rect 19797 27619 19855 27625
rect 21358 27616 21364 27628
rect 21416 27616 21422 27668
rect 24394 27616 24400 27668
rect 24452 27656 24458 27668
rect 24581 27659 24639 27665
rect 24581 27656 24593 27659
rect 24452 27628 24593 27656
rect 24452 27616 24458 27628
rect 24581 27625 24593 27628
rect 24627 27625 24639 27659
rect 24581 27619 24639 27625
rect 24762 27616 24768 27668
rect 24820 27616 24826 27668
rect 26234 27616 26240 27668
rect 26292 27616 26298 27668
rect 26326 27616 26332 27668
rect 26384 27616 26390 27668
rect 31754 27616 31760 27668
rect 31812 27616 31818 27668
rect 34514 27616 34520 27668
rect 34572 27616 34578 27668
rect 22649 27591 22707 27597
rect 22649 27557 22661 27591
rect 22695 27588 22707 27591
rect 23382 27588 23388 27600
rect 22695 27560 23388 27588
rect 22695 27557 22707 27560
rect 22649 27551 22707 27557
rect 23382 27548 23388 27560
rect 23440 27548 23446 27600
rect 20257 27523 20315 27529
rect 20257 27520 20269 27523
rect 19352 27492 20269 27520
rect 19352 27464 19380 27492
rect 20257 27489 20269 27492
rect 20303 27489 20315 27523
rect 20257 27483 20315 27489
rect 22373 27523 22431 27529
rect 22373 27489 22385 27523
rect 22419 27520 22431 27523
rect 22462 27520 22468 27532
rect 22419 27492 22468 27520
rect 22419 27489 22431 27492
rect 22373 27483 22431 27489
rect 22462 27480 22468 27492
rect 22520 27480 22526 27532
rect 25225 27523 25283 27529
rect 24320 27492 25176 27520
rect 19242 27412 19248 27464
rect 19300 27412 19306 27464
rect 19334 27412 19340 27464
rect 19392 27412 19398 27464
rect 19426 27412 19432 27464
rect 19484 27452 19490 27464
rect 19521 27455 19579 27461
rect 19521 27452 19533 27455
rect 19484 27424 19533 27452
rect 19484 27412 19490 27424
rect 19521 27421 19533 27424
rect 19567 27421 19579 27455
rect 19521 27415 19579 27421
rect 19613 27455 19671 27461
rect 19613 27421 19625 27455
rect 19659 27421 19671 27455
rect 19613 27415 19671 27421
rect 18966 27384 18972 27396
rect 17604 27356 18972 27384
rect 17604 27328 17632 27356
rect 18966 27344 18972 27356
rect 19024 27384 19030 27396
rect 19628 27384 19656 27415
rect 19978 27412 19984 27464
rect 20036 27412 20042 27464
rect 20070 27412 20076 27464
rect 20128 27412 20134 27464
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27452 20223 27455
rect 22281 27455 22339 27461
rect 22281 27452 22293 27455
rect 20211 27424 20300 27452
rect 20211 27421 20223 27424
rect 20165 27415 20223 27421
rect 19024 27356 19656 27384
rect 19024 27344 19030 27356
rect 20272 27328 20300 27424
rect 22204 27424 22293 27452
rect 22204 27328 22232 27424
rect 22281 27421 22293 27424
rect 22327 27421 22339 27455
rect 22281 27415 22339 27421
rect 17586 27276 17592 27328
rect 17644 27276 17650 27328
rect 20254 27276 20260 27328
rect 20312 27276 20318 27328
rect 20438 27276 20444 27328
rect 20496 27276 20502 27328
rect 22186 27276 22192 27328
rect 22244 27276 22250 27328
rect 23198 27276 23204 27328
rect 23256 27316 23262 27328
rect 24320 27316 24348 27492
rect 24486 27412 24492 27464
rect 24544 27452 24550 27464
rect 24857 27455 24915 27461
rect 24857 27452 24869 27455
rect 24544 27424 24869 27452
rect 24544 27412 24550 27424
rect 24857 27421 24869 27424
rect 24903 27421 24915 27455
rect 24857 27415 24915 27421
rect 25041 27455 25099 27461
rect 25041 27421 25053 27455
rect 25087 27421 25099 27455
rect 25041 27415 25099 27421
rect 24397 27387 24455 27393
rect 24397 27353 24409 27387
rect 24443 27384 24455 27387
rect 25056 27384 25084 27415
rect 24443 27356 25084 27384
rect 25148 27384 25176 27492
rect 25225 27489 25237 27523
rect 25271 27520 25283 27523
rect 27706 27520 27712 27532
rect 25271 27492 27712 27520
rect 25271 27489 25283 27492
rect 25225 27483 25283 27489
rect 27706 27480 27712 27492
rect 27764 27520 27770 27532
rect 28077 27523 28135 27529
rect 27764 27492 28028 27520
rect 27764 27480 27770 27492
rect 25406 27412 25412 27464
rect 25464 27452 25470 27464
rect 25685 27455 25743 27461
rect 25685 27452 25697 27455
rect 25464 27424 25697 27452
rect 25464 27412 25470 27424
rect 25685 27421 25697 27424
rect 25731 27421 25743 27455
rect 25685 27415 25743 27421
rect 25777 27455 25835 27461
rect 25777 27421 25789 27455
rect 25823 27421 25835 27455
rect 25777 27415 25835 27421
rect 25792 27384 25820 27415
rect 25958 27412 25964 27464
rect 26016 27412 26022 27464
rect 26053 27455 26111 27461
rect 26053 27421 26065 27455
rect 26099 27452 26111 27455
rect 26142 27452 26148 27464
rect 26099 27424 26148 27452
rect 26099 27421 26111 27424
rect 26053 27415 26111 27421
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 28000 27461 28028 27492
rect 28077 27489 28089 27523
rect 28123 27489 28135 27523
rect 28077 27483 28135 27489
rect 28353 27523 28411 27529
rect 28353 27489 28365 27523
rect 28399 27520 28411 27523
rect 28629 27523 28687 27529
rect 28629 27520 28641 27523
rect 28399 27492 28641 27520
rect 28399 27489 28411 27492
rect 28353 27483 28411 27489
rect 28629 27489 28641 27492
rect 28675 27489 28687 27523
rect 31662 27520 31668 27532
rect 28629 27483 28687 27489
rect 31404 27492 31668 27520
rect 26605 27455 26663 27461
rect 26605 27421 26617 27455
rect 26651 27421 26663 27455
rect 26605 27415 26663 27421
rect 27985 27455 28043 27461
rect 27985 27421 27997 27455
rect 28031 27421 28043 27455
rect 27985 27415 28043 27421
rect 26326 27384 26332 27396
rect 25148 27356 26332 27384
rect 24443 27353 24455 27356
rect 24397 27347 24455 27353
rect 25056 27328 25084 27356
rect 26326 27344 26332 27356
rect 26384 27344 26390 27396
rect 26418 27344 26424 27396
rect 26476 27384 26482 27396
rect 26620 27384 26648 27415
rect 27522 27384 27528 27396
rect 26476 27356 27528 27384
rect 26476 27344 26482 27356
rect 27522 27344 27528 27356
rect 27580 27384 27586 27396
rect 28092 27384 28120 27483
rect 28534 27412 28540 27464
rect 28592 27452 28598 27464
rect 31404 27461 31432 27492
rect 31662 27480 31668 27492
rect 31720 27480 31726 27532
rect 32122 27480 32128 27532
rect 32180 27480 32186 27532
rect 32582 27480 32588 27532
rect 32640 27520 32646 27532
rect 32769 27523 32827 27529
rect 32769 27520 32781 27523
rect 32640 27492 32781 27520
rect 32640 27480 32646 27492
rect 32769 27489 32781 27492
rect 32815 27489 32827 27523
rect 32769 27483 32827 27489
rect 28721 27455 28779 27461
rect 28721 27452 28733 27455
rect 28592 27424 28733 27452
rect 28592 27412 28598 27424
rect 28721 27421 28733 27424
rect 28767 27421 28779 27455
rect 28721 27415 28779 27421
rect 31389 27455 31447 27461
rect 31389 27421 31401 27455
rect 31435 27421 31447 27455
rect 32033 27455 32091 27461
rect 32033 27452 32045 27455
rect 31389 27415 31447 27421
rect 31726 27424 32045 27452
rect 27580 27356 28120 27384
rect 31573 27387 31631 27393
rect 27580 27344 27586 27356
rect 31573 27353 31585 27387
rect 31619 27384 31631 27387
rect 31726 27384 31754 27424
rect 32033 27421 32045 27424
rect 32079 27421 32091 27455
rect 32033 27415 32091 27421
rect 34514 27412 34520 27464
rect 34572 27452 34578 27464
rect 34701 27455 34759 27461
rect 34701 27452 34713 27455
rect 34572 27424 34713 27452
rect 34572 27412 34578 27424
rect 34701 27421 34713 27424
rect 34747 27421 34759 27455
rect 34701 27415 34759 27421
rect 33045 27387 33103 27393
rect 33045 27384 33057 27387
rect 31619 27356 31754 27384
rect 32416 27356 33057 27384
rect 31619 27353 31631 27356
rect 31573 27347 31631 27353
rect 24597 27319 24655 27325
rect 24597 27316 24609 27319
rect 23256 27288 24609 27316
rect 23256 27276 23262 27288
rect 24597 27285 24609 27288
rect 24643 27285 24655 27319
rect 24597 27279 24655 27285
rect 25038 27276 25044 27328
rect 25096 27276 25102 27328
rect 25866 27276 25872 27328
rect 25924 27316 25930 27328
rect 26513 27319 26571 27325
rect 26513 27316 26525 27319
rect 25924 27288 26525 27316
rect 25924 27276 25930 27288
rect 26513 27285 26525 27288
rect 26559 27285 26571 27319
rect 26513 27279 26571 27285
rect 29086 27276 29092 27328
rect 29144 27276 29150 27328
rect 31478 27276 31484 27328
rect 31536 27316 31542 27328
rect 31588 27316 31616 27347
rect 32416 27325 32444 27356
rect 33045 27353 33057 27356
rect 33091 27353 33103 27387
rect 34793 27387 34851 27393
rect 34793 27384 34805 27387
rect 34270 27356 34805 27384
rect 33045 27347 33103 27353
rect 34793 27353 34805 27356
rect 34839 27353 34851 27387
rect 34793 27347 34851 27353
rect 31536 27288 31616 27316
rect 32401 27319 32459 27325
rect 31536 27276 31542 27288
rect 32401 27285 32413 27319
rect 32447 27285 32459 27319
rect 32401 27279 32459 27285
rect 1104 27226 35236 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 35236 27226
rect 1104 27152 35236 27174
rect 17586 27072 17592 27124
rect 17644 27072 17650 27124
rect 18966 27072 18972 27124
rect 19024 27072 19030 27124
rect 19242 27072 19248 27124
rect 19300 27112 19306 27124
rect 19429 27115 19487 27121
rect 19429 27112 19441 27115
rect 19300 27084 19441 27112
rect 19300 27072 19306 27084
rect 19429 27081 19441 27084
rect 19475 27081 19487 27115
rect 19429 27075 19487 27081
rect 19978 27072 19984 27124
rect 20036 27112 20042 27124
rect 20165 27115 20223 27121
rect 20165 27112 20177 27115
rect 20036 27084 20177 27112
rect 20036 27072 20042 27084
rect 20165 27081 20177 27084
rect 20211 27081 20223 27115
rect 20165 27075 20223 27081
rect 20438 27072 20444 27124
rect 20496 27072 20502 27124
rect 20625 27115 20683 27121
rect 20625 27081 20637 27115
rect 20671 27112 20683 27115
rect 24394 27112 24400 27124
rect 20671 27084 24400 27112
rect 20671 27081 20683 27084
rect 20625 27075 20683 27081
rect 24394 27072 24400 27084
rect 24452 27072 24458 27124
rect 24486 27072 24492 27124
rect 24544 27072 24550 27124
rect 25130 27112 25136 27124
rect 24688 27084 25136 27112
rect 18984 27044 19012 27072
rect 20254 27044 20260 27056
rect 18892 27016 19012 27044
rect 19076 27016 20260 27044
rect 13354 26936 13360 26988
rect 13412 26936 13418 26988
rect 17405 26979 17463 26985
rect 17405 26976 17417 26979
rect 17236 26948 17417 26976
rect 13170 26868 13176 26920
rect 13228 26868 13234 26920
rect 17236 26908 17264 26948
rect 17405 26945 17417 26948
rect 17451 26945 17463 26979
rect 17405 26939 17463 26945
rect 17494 26936 17500 26988
rect 17552 26976 17558 26988
rect 17589 26979 17647 26985
rect 17589 26976 17601 26979
rect 17552 26948 17601 26976
rect 17552 26936 17558 26948
rect 17589 26945 17601 26948
rect 17635 26976 17647 26979
rect 17681 26979 17739 26985
rect 17681 26976 17693 26979
rect 17635 26948 17693 26976
rect 17635 26945 17647 26948
rect 17589 26939 17647 26945
rect 17681 26945 17693 26948
rect 17727 26945 17739 26979
rect 17681 26939 17739 26945
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26945 17923 26979
rect 17865 26939 17923 26945
rect 17880 26908 17908 26939
rect 18782 26936 18788 26988
rect 18840 26936 18846 26988
rect 18892 26976 18920 27016
rect 19076 26988 19104 27016
rect 18964 26979 19022 26985
rect 18964 26976 18976 26979
rect 18892 26948 18976 26976
rect 18964 26945 18976 26948
rect 19010 26945 19022 26979
rect 18964 26939 19022 26945
rect 19058 26936 19064 26988
rect 19116 26936 19122 26988
rect 19812 26985 19840 27016
rect 20254 27004 20260 27016
rect 20312 27004 20318 27056
rect 19153 26979 19211 26985
rect 19153 26945 19165 26979
rect 19199 26976 19211 26979
rect 19521 26979 19579 26985
rect 19521 26976 19533 26979
rect 19199 26948 19533 26976
rect 19199 26945 19211 26948
rect 19153 26939 19211 26945
rect 19521 26945 19533 26948
rect 19567 26945 19579 26979
rect 19521 26939 19579 26945
rect 19705 26979 19763 26985
rect 19705 26945 19717 26979
rect 19751 26945 19763 26979
rect 19705 26939 19763 26945
rect 19797 26979 19855 26985
rect 19797 26945 19809 26979
rect 19843 26945 19855 26979
rect 19797 26939 19855 26945
rect 19889 26979 19947 26985
rect 19889 26945 19901 26979
rect 19935 26976 19947 26979
rect 20070 26976 20076 26988
rect 19935 26948 20076 26976
rect 19935 26945 19947 26948
rect 19889 26939 19947 26945
rect 17236 26880 17908 26908
rect 17236 26784 17264 26880
rect 18874 26868 18880 26920
rect 18932 26908 18938 26920
rect 19168 26908 19196 26939
rect 18932 26880 19196 26908
rect 18932 26868 18938 26880
rect 17865 26843 17923 26849
rect 17865 26809 17877 26843
rect 17911 26840 17923 26843
rect 19334 26840 19340 26852
rect 17911 26812 19340 26840
rect 17911 26809 17923 26812
rect 17865 26803 17923 26809
rect 19334 26800 19340 26812
rect 19392 26840 19398 26852
rect 19720 26840 19748 26939
rect 19392 26812 19748 26840
rect 19392 26800 19398 26812
rect 13538 26732 13544 26784
rect 13596 26732 13602 26784
rect 15381 26775 15439 26781
rect 15381 26741 15393 26775
rect 15427 26772 15439 26775
rect 15930 26772 15936 26784
rect 15427 26744 15936 26772
rect 15427 26741 15439 26744
rect 15381 26735 15439 26741
rect 15930 26732 15936 26744
rect 15988 26732 15994 26784
rect 16025 26775 16083 26781
rect 16025 26741 16037 26775
rect 16071 26772 16083 26775
rect 16114 26772 16120 26784
rect 16071 26744 16120 26772
rect 16071 26741 16083 26744
rect 16025 26735 16083 26741
rect 16114 26732 16120 26744
rect 16172 26732 16178 26784
rect 17218 26732 17224 26784
rect 17276 26732 17282 26784
rect 18506 26732 18512 26784
rect 18564 26772 18570 26784
rect 18782 26772 18788 26784
rect 18564 26744 18788 26772
rect 18564 26732 18570 26744
rect 18782 26732 18788 26744
rect 18840 26772 18846 26784
rect 19242 26772 19248 26784
rect 18840 26744 19248 26772
rect 18840 26732 18846 26744
rect 19242 26732 19248 26744
rect 19300 26772 19306 26784
rect 19904 26772 19932 26939
rect 20070 26936 20076 26948
rect 20128 26936 20134 26988
rect 20456 26976 20484 27072
rect 20990 27004 20996 27056
rect 21048 27044 21054 27056
rect 22094 27044 22100 27056
rect 21048 27016 22100 27044
rect 21048 27004 21054 27016
rect 22094 27004 22100 27016
rect 22152 27004 22158 27056
rect 24412 27044 24440 27072
rect 24688 27044 24716 27084
rect 25130 27072 25136 27084
rect 25188 27072 25194 27124
rect 25777 27115 25835 27121
rect 25777 27081 25789 27115
rect 25823 27112 25835 27115
rect 26142 27112 26148 27124
rect 25823 27084 26148 27112
rect 25823 27081 25835 27084
rect 25777 27075 25835 27081
rect 26142 27072 26148 27084
rect 26200 27072 26206 27124
rect 26234 27072 26240 27124
rect 26292 27072 26298 27124
rect 26326 27072 26332 27124
rect 26384 27112 26390 27124
rect 26697 27115 26755 27121
rect 26697 27112 26709 27115
rect 26384 27084 26709 27112
rect 26384 27072 26390 27084
rect 26697 27081 26709 27084
rect 26743 27081 26755 27115
rect 26697 27075 26755 27081
rect 27065 27115 27123 27121
rect 27065 27081 27077 27115
rect 27111 27112 27123 27115
rect 28534 27112 28540 27124
rect 27111 27084 28540 27112
rect 27111 27081 27123 27084
rect 27065 27075 27123 27081
rect 28534 27072 28540 27084
rect 28592 27072 28598 27124
rect 29086 27072 29092 27124
rect 29144 27072 29150 27124
rect 29549 27115 29607 27121
rect 29549 27081 29561 27115
rect 29595 27112 29607 27115
rect 29638 27112 29644 27124
rect 29595 27084 29644 27112
rect 29595 27081 29607 27084
rect 29549 27075 29607 27081
rect 29638 27072 29644 27084
rect 29696 27112 29702 27124
rect 29822 27112 29828 27124
rect 29696 27084 29828 27112
rect 29696 27072 29702 27084
rect 29822 27072 29828 27084
rect 29880 27072 29886 27124
rect 31389 27115 31447 27121
rect 31389 27081 31401 27115
rect 31435 27112 31447 27115
rect 31478 27112 31484 27124
rect 31435 27084 31484 27112
rect 31435 27081 31447 27084
rect 31389 27075 31447 27081
rect 31478 27072 31484 27084
rect 31536 27072 31542 27124
rect 32122 27072 32128 27124
rect 32180 27112 32186 27124
rect 32217 27115 32275 27121
rect 32217 27112 32229 27115
rect 32180 27084 32229 27112
rect 32180 27072 32186 27084
rect 32217 27081 32229 27084
rect 32263 27081 32275 27115
rect 32217 27075 32275 27081
rect 32582 27072 32588 27124
rect 32640 27072 32646 27124
rect 25222 27044 25228 27056
rect 24412 27016 24716 27044
rect 24780 27016 25228 27044
rect 24780 26988 24808 27016
rect 25222 27004 25228 27016
rect 25280 27004 25286 27056
rect 25406 27004 25412 27056
rect 25464 27044 25470 27056
rect 25501 27047 25559 27053
rect 25501 27044 25513 27047
rect 25464 27016 25513 27044
rect 25464 27004 25470 27016
rect 25501 27013 25513 27016
rect 25547 27044 25559 27047
rect 25866 27044 25872 27056
rect 25547 27016 25872 27044
rect 25547 27013 25559 27016
rect 25501 27007 25559 27013
rect 25866 27004 25872 27016
rect 25924 27044 25930 27056
rect 25924 27016 26004 27044
rect 25924 27004 25930 27016
rect 20533 26979 20591 26985
rect 20533 26976 20545 26979
rect 20456 26948 20545 26976
rect 20533 26945 20545 26948
rect 20579 26945 20591 26979
rect 20533 26939 20591 26945
rect 21266 26936 21272 26988
rect 21324 26936 21330 26988
rect 21358 26936 21364 26988
rect 21416 26936 21422 26988
rect 22462 26936 22468 26988
rect 22520 26936 22526 26988
rect 23198 26936 23204 26988
rect 23256 26936 23262 26988
rect 24302 26936 24308 26988
rect 24360 26976 24366 26988
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24360 26948 24409 26976
rect 24360 26936 24366 26948
rect 24397 26945 24409 26948
rect 24443 26945 24455 26979
rect 24397 26939 24455 26945
rect 24581 26979 24639 26985
rect 24581 26945 24593 26979
rect 24627 26976 24639 26979
rect 24673 26979 24731 26985
rect 24673 26976 24685 26979
rect 24627 26948 24685 26976
rect 24627 26945 24639 26948
rect 24581 26939 24639 26945
rect 24673 26945 24685 26948
rect 24719 26976 24731 26979
rect 24762 26976 24768 26988
rect 24719 26948 24768 26976
rect 24719 26945 24731 26948
rect 24673 26939 24731 26945
rect 22373 26911 22431 26917
rect 22373 26877 22385 26911
rect 22419 26877 22431 26911
rect 24412 26908 24440 26939
rect 24762 26936 24768 26948
rect 24820 26936 24826 26988
rect 24857 26979 24915 26985
rect 24857 26945 24869 26979
rect 24903 26945 24915 26979
rect 24857 26939 24915 26945
rect 24872 26908 24900 26939
rect 25130 26936 25136 26988
rect 25188 26976 25194 26988
rect 25976 26985 26004 27016
rect 25317 26979 25375 26985
rect 25317 26976 25329 26979
rect 25188 26948 25329 26976
rect 25188 26936 25194 26948
rect 25317 26945 25329 26948
rect 25363 26945 25375 26979
rect 25317 26939 25375 26945
rect 25961 26979 26019 26985
rect 25961 26945 25973 26979
rect 26007 26945 26019 26979
rect 25961 26939 26019 26945
rect 26050 26936 26056 26988
rect 26108 26936 26114 26988
rect 26145 26982 26203 26985
rect 26252 26982 26280 27072
rect 29104 27044 29132 27072
rect 29917 27047 29975 27053
rect 29917 27044 29929 27047
rect 29104 27016 29929 27044
rect 29917 27013 29929 27016
rect 29963 27013 29975 27047
rect 31573 27047 31631 27053
rect 31573 27044 31585 27047
rect 31142 27016 31585 27044
rect 29917 27007 29975 27013
rect 31573 27013 31585 27016
rect 31619 27013 31631 27047
rect 31573 27007 31631 27013
rect 26145 26979 26280 26982
rect 26145 26945 26157 26979
rect 26191 26954 26280 26979
rect 26191 26945 26203 26954
rect 26145 26939 26203 26945
rect 26326 26936 26332 26988
rect 26384 26936 26390 26988
rect 26421 26979 26479 26985
rect 26421 26945 26433 26979
rect 26467 26976 26479 26979
rect 26513 26979 26571 26985
rect 26513 26976 26525 26979
rect 26467 26948 26525 26976
rect 26467 26945 26479 26948
rect 26421 26939 26479 26945
rect 26513 26945 26525 26948
rect 26559 26945 26571 26979
rect 26513 26939 26571 26945
rect 24412 26880 24900 26908
rect 22373 26871 22431 26877
rect 22186 26800 22192 26852
rect 22244 26840 22250 26852
rect 22388 26840 22416 26871
rect 22244 26812 22416 26840
rect 24872 26840 24900 26880
rect 25682 26868 25688 26920
rect 25740 26868 25746 26920
rect 26436 26840 26464 26939
rect 26786 26936 26792 26988
rect 26844 26936 26850 26988
rect 26973 26979 27031 26985
rect 26973 26945 26985 26979
rect 27019 26976 27031 26979
rect 27062 26976 27068 26988
rect 27019 26948 27068 26976
rect 27019 26945 27031 26948
rect 26973 26939 27031 26945
rect 27062 26936 27068 26948
rect 27120 26936 27126 26988
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26976 27215 26979
rect 27246 26976 27252 26988
rect 27203 26948 27252 26976
rect 27203 26945 27215 26948
rect 27157 26939 27215 26945
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 31294 26936 31300 26988
rect 31352 26976 31358 26988
rect 31481 26979 31539 26985
rect 31481 26976 31493 26979
rect 31352 26948 31493 26976
rect 31352 26936 31358 26948
rect 31481 26945 31493 26948
rect 31527 26945 31539 26979
rect 31481 26939 31539 26945
rect 31662 26936 31668 26988
rect 31720 26976 31726 26988
rect 32125 26979 32183 26985
rect 32125 26976 32137 26979
rect 31720 26948 32137 26976
rect 31720 26936 31726 26948
rect 32125 26945 32137 26948
rect 32171 26945 32183 26979
rect 32125 26939 32183 26945
rect 32306 26936 32312 26988
rect 32364 26936 32370 26988
rect 34698 26936 34704 26988
rect 34756 26936 34762 26988
rect 34790 26936 34796 26988
rect 34848 26936 34854 26988
rect 29638 26868 29644 26920
rect 29696 26868 29702 26920
rect 34425 26911 34483 26917
rect 34425 26877 34437 26911
rect 34471 26908 34483 26911
rect 34808 26908 34836 26936
rect 34471 26880 34836 26908
rect 34471 26877 34483 26880
rect 34425 26871 34483 26877
rect 24872 26812 26004 26840
rect 22244 26800 22250 26812
rect 19300 26744 19932 26772
rect 19300 26732 19306 26744
rect 22922 26732 22928 26784
rect 22980 26772 22986 26784
rect 23477 26775 23535 26781
rect 23477 26772 23489 26775
rect 22980 26744 23489 26772
rect 22980 26732 22986 26744
rect 23477 26741 23489 26744
rect 23523 26741 23535 26775
rect 23477 26735 23535 26741
rect 23566 26732 23572 26784
rect 23624 26772 23630 26784
rect 23845 26775 23903 26781
rect 23845 26772 23857 26775
rect 23624 26744 23857 26772
rect 23624 26732 23630 26744
rect 23845 26741 23857 26744
rect 23891 26741 23903 26775
rect 23845 26735 23903 26741
rect 25038 26732 25044 26784
rect 25096 26772 25102 26784
rect 25866 26772 25872 26784
rect 25096 26744 25872 26772
rect 25096 26732 25102 26744
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 25976 26772 26004 26812
rect 26160 26812 26464 26840
rect 26160 26772 26188 26812
rect 26510 26800 26516 26852
rect 26568 26800 26574 26852
rect 25976 26744 26188 26772
rect 1104 26682 35248 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 35248 26682
rect 1104 26608 35248 26630
rect 13081 26571 13139 26577
rect 13081 26537 13093 26571
rect 13127 26537 13139 26571
rect 13081 26531 13139 26537
rect 13096 26500 13124 26531
rect 13170 26528 13176 26580
rect 13228 26568 13234 26580
rect 13357 26571 13415 26577
rect 13357 26568 13369 26571
rect 13228 26540 13369 26568
rect 13228 26528 13234 26540
rect 13357 26537 13369 26540
rect 13403 26537 13415 26571
rect 13357 26531 13415 26537
rect 13538 26528 13544 26580
rect 13596 26528 13602 26580
rect 15381 26571 15439 26577
rect 15381 26537 15393 26571
rect 15427 26568 15439 26571
rect 16390 26568 16396 26580
rect 15427 26540 16396 26568
rect 15427 26537 15439 26540
rect 15381 26531 15439 26537
rect 16390 26528 16396 26540
rect 16448 26528 16454 26580
rect 19981 26571 20039 26577
rect 19981 26537 19993 26571
rect 20027 26568 20039 26571
rect 20990 26568 20996 26580
rect 20027 26540 20996 26568
rect 20027 26537 20039 26540
rect 19981 26531 20039 26537
rect 20990 26528 20996 26540
rect 21048 26528 21054 26580
rect 22186 26528 22192 26580
rect 22244 26528 22250 26580
rect 22462 26528 22468 26580
rect 22520 26528 22526 26580
rect 23845 26571 23903 26577
rect 23845 26537 23857 26571
rect 23891 26568 23903 26571
rect 24670 26568 24676 26580
rect 23891 26540 24676 26568
rect 23891 26537 23903 26540
rect 23845 26531 23903 26537
rect 24670 26528 24676 26540
rect 24728 26528 24734 26580
rect 25958 26528 25964 26580
rect 26016 26568 26022 26580
rect 26237 26571 26295 26577
rect 26237 26568 26249 26571
rect 26016 26540 26249 26568
rect 26016 26528 26022 26540
rect 26237 26537 26249 26540
rect 26283 26537 26295 26571
rect 26237 26531 26295 26537
rect 32582 26528 32588 26580
rect 32640 26528 32646 26580
rect 34517 26571 34575 26577
rect 34517 26537 34529 26571
rect 34563 26568 34575 26571
rect 34698 26568 34704 26580
rect 34563 26540 34704 26568
rect 34563 26537 34575 26540
rect 34517 26531 34575 26537
rect 34698 26528 34704 26540
rect 34756 26528 34762 26580
rect 13262 26500 13268 26512
rect 13096 26472 13268 26500
rect 13262 26460 13268 26472
rect 13320 26460 13326 26512
rect 13556 26500 13584 26528
rect 15565 26503 15623 26509
rect 13556 26472 14596 26500
rect 11992 26404 13676 26432
rect 11992 26376 12020 26404
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 11974 26324 11980 26376
rect 12032 26324 12038 26376
rect 12986 26324 12992 26376
rect 13044 26324 13050 26376
rect 13078 26324 13084 26376
rect 13136 26364 13142 26376
rect 13648 26373 13676 26404
rect 14568 26373 14596 26472
rect 15565 26469 15577 26503
rect 15611 26500 15623 26503
rect 17034 26500 17040 26512
rect 15611 26472 17040 26500
rect 15611 26469 15623 26472
rect 15565 26463 15623 26469
rect 17034 26460 17040 26472
rect 17092 26460 17098 26512
rect 19061 26503 19119 26509
rect 19061 26469 19073 26503
rect 19107 26500 19119 26503
rect 19613 26503 19671 26509
rect 19613 26500 19625 26503
rect 19107 26472 19625 26500
rect 19107 26469 19119 26472
rect 19061 26463 19119 26469
rect 19613 26469 19625 26472
rect 19659 26469 19671 26503
rect 23201 26503 23259 26509
rect 19613 26463 19671 26469
rect 20732 26472 22416 26500
rect 15933 26435 15991 26441
rect 15933 26401 15945 26435
rect 15979 26432 15991 26435
rect 15979 26404 16252 26432
rect 15979 26401 15991 26404
rect 15933 26395 15991 26401
rect 16224 26373 16252 26404
rect 18138 26392 18144 26444
rect 18196 26432 18202 26444
rect 18233 26435 18291 26441
rect 18233 26432 18245 26435
rect 18196 26404 18245 26432
rect 18196 26392 18202 26404
rect 18233 26401 18245 26404
rect 18279 26432 18291 26435
rect 18279 26404 19196 26432
rect 18279 26401 18291 26404
rect 18233 26395 18291 26401
rect 13265 26367 13323 26373
rect 13265 26364 13277 26367
rect 13136 26336 13277 26364
rect 13136 26324 13142 26336
rect 13265 26333 13277 26336
rect 13311 26333 13323 26367
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 13265 26327 13323 26333
rect 13372 26336 13553 26364
rect 11054 26256 11060 26308
rect 11112 26296 11118 26308
rect 12526 26296 12532 26308
rect 11112 26268 12532 26296
rect 11112 26256 11118 26268
rect 12526 26256 12532 26268
rect 12584 26296 12590 26308
rect 13372 26296 13400 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13633 26367 13691 26373
rect 13633 26333 13645 26367
rect 13679 26333 13691 26367
rect 13633 26327 13691 26333
rect 13817 26367 13875 26373
rect 13817 26333 13829 26367
rect 13863 26333 13875 26367
rect 13817 26327 13875 26333
rect 13909 26367 13967 26373
rect 13909 26333 13921 26367
rect 13955 26333 13967 26367
rect 13909 26327 13967 26333
rect 14553 26367 14611 26373
rect 14553 26333 14565 26367
rect 14599 26333 14611 26367
rect 14553 26327 14611 26333
rect 14737 26367 14795 26373
rect 14737 26333 14749 26367
rect 14783 26364 14795 26367
rect 15473 26367 15531 26373
rect 15473 26364 15485 26367
rect 14783 26336 15485 26364
rect 14783 26333 14795 26336
rect 14737 26327 14795 26333
rect 15473 26333 15485 26336
rect 15519 26333 15531 26367
rect 15473 26327 15531 26333
rect 15749 26367 15807 26373
rect 15749 26333 15761 26367
rect 15795 26364 15807 26367
rect 16025 26367 16083 26373
rect 15795 26336 15976 26364
rect 15795 26333 15807 26336
rect 15749 26327 15807 26333
rect 13832 26296 13860 26327
rect 12584 26268 13400 26296
rect 13648 26268 13860 26296
rect 12584 26256 12590 26268
rect 13648 26240 13676 26268
rect 13924 26240 13952 26327
rect 1581 26231 1639 26237
rect 1581 26197 1593 26231
rect 1627 26228 1639 26231
rect 1854 26228 1860 26240
rect 1627 26200 1860 26228
rect 1627 26197 1639 26200
rect 1581 26191 1639 26197
rect 1854 26188 1860 26200
rect 1912 26188 1918 26240
rect 9490 26188 9496 26240
rect 9548 26188 9554 26240
rect 12710 26188 12716 26240
rect 12768 26188 12774 26240
rect 13630 26188 13636 26240
rect 13688 26188 13694 26240
rect 13906 26188 13912 26240
rect 13964 26188 13970 26240
rect 15488 26228 15516 26327
rect 15948 26308 15976 26336
rect 16025 26333 16037 26367
rect 16071 26333 16083 26367
rect 16025 26327 16083 26333
rect 16209 26367 16267 26373
rect 16209 26333 16221 26367
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 15930 26256 15936 26308
rect 15988 26256 15994 26308
rect 16040 26296 16068 26327
rect 16482 26324 16488 26376
rect 16540 26324 16546 26376
rect 16669 26367 16727 26373
rect 16669 26333 16681 26367
rect 16715 26364 16727 26367
rect 17218 26364 17224 26376
rect 16715 26336 17224 26364
rect 16715 26333 16727 26336
rect 16669 26327 16727 26333
rect 17218 26324 17224 26336
rect 17276 26324 17282 26376
rect 17402 26324 17408 26376
rect 17460 26324 17466 26376
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 18506 26364 18512 26376
rect 18463 26336 18512 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 18506 26324 18512 26336
rect 18564 26324 18570 26376
rect 18616 26373 18644 26404
rect 19168 26376 19196 26404
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 19521 26435 19579 26441
rect 19521 26432 19533 26435
rect 19392 26404 19533 26432
rect 19392 26392 19398 26404
rect 19521 26401 19533 26404
rect 19567 26401 19579 26435
rect 19521 26395 19579 26401
rect 18601 26367 18659 26373
rect 18601 26333 18613 26367
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26333 18751 26367
rect 18693 26327 18751 26333
rect 16574 26296 16580 26308
rect 16040 26268 16580 26296
rect 16574 26256 16580 26268
rect 16632 26256 16638 26308
rect 18708 26296 18736 26327
rect 18782 26324 18788 26376
rect 18840 26324 18846 26376
rect 19058 26324 19064 26376
rect 19116 26324 19122 26376
rect 19150 26324 19156 26376
rect 19208 26364 19214 26376
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 19208 26336 19257 26364
rect 19208 26324 19214 26336
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 19426 26324 19432 26376
rect 19484 26324 19490 26376
rect 19705 26367 19763 26373
rect 19705 26333 19717 26367
rect 19751 26333 19763 26367
rect 19705 26327 19763 26333
rect 19076 26296 19104 26324
rect 18708 26268 19104 26296
rect 16298 26228 16304 26240
rect 15488 26200 16304 26228
rect 16298 26188 16304 26200
rect 16356 26188 16362 26240
rect 17037 26231 17095 26237
rect 17037 26197 17049 26231
rect 17083 26228 17095 26231
rect 17126 26228 17132 26240
rect 17083 26200 17132 26228
rect 17083 26197 17095 26200
rect 17037 26191 17095 26197
rect 17126 26188 17132 26200
rect 17184 26188 17190 26240
rect 18230 26188 18236 26240
rect 18288 26228 18294 26240
rect 19720 26228 19748 26327
rect 20732 26240 20760 26472
rect 21082 26392 21088 26444
rect 21140 26392 21146 26444
rect 21468 26404 22324 26432
rect 21468 26308 21496 26404
rect 22296 26373 22324 26404
rect 22388 26373 22416 26472
rect 23201 26469 23213 26503
rect 23247 26500 23259 26503
rect 24302 26500 24308 26512
rect 23247 26472 24308 26500
rect 23247 26469 23259 26472
rect 23201 26463 23259 26469
rect 22833 26435 22891 26441
rect 22833 26432 22845 26435
rect 22572 26404 22845 26432
rect 22572 26373 22600 26404
rect 22833 26401 22845 26404
rect 22879 26432 22891 26435
rect 22922 26432 22928 26444
rect 22879 26404 22928 26432
rect 22879 26401 22891 26404
rect 22833 26395 22891 26401
rect 22922 26392 22928 26404
rect 22980 26392 22986 26444
rect 23385 26435 23443 26441
rect 23385 26401 23397 26435
rect 23431 26432 23443 26435
rect 23750 26432 23756 26444
rect 23431 26404 23756 26432
rect 23431 26401 23443 26404
rect 23385 26395 23443 26401
rect 23750 26392 23756 26404
rect 23808 26392 23814 26444
rect 22097 26367 22155 26373
rect 22097 26364 22109 26367
rect 22020 26336 22109 26364
rect 21450 26256 21456 26308
rect 21508 26256 21514 26308
rect 22020 26296 22048 26336
rect 22097 26333 22109 26336
rect 22143 26333 22155 26367
rect 22097 26327 22155 26333
rect 22281 26367 22339 26373
rect 22281 26333 22293 26367
rect 22327 26333 22339 26367
rect 22281 26327 22339 26333
rect 22373 26367 22431 26373
rect 22373 26333 22385 26367
rect 22419 26333 22431 26367
rect 22373 26327 22431 26333
rect 22557 26367 22615 26373
rect 22557 26333 22569 26367
rect 22603 26333 22615 26367
rect 22557 26327 22615 26333
rect 23017 26367 23075 26373
rect 23017 26333 23029 26367
rect 23063 26333 23075 26367
rect 23017 26327 23075 26333
rect 23032 26296 23060 26327
rect 23290 26324 23296 26376
rect 23348 26364 23354 26376
rect 23477 26367 23535 26373
rect 23477 26364 23489 26367
rect 23348 26336 23489 26364
rect 23348 26324 23354 26336
rect 23477 26333 23489 26336
rect 23523 26333 23535 26367
rect 23477 26327 23535 26333
rect 23566 26324 23572 26376
rect 23624 26324 23630 26376
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26364 23719 26367
rect 23860 26364 23888 26472
rect 24302 26460 24308 26472
rect 24360 26460 24366 26512
rect 32600 26432 32628 26528
rect 32769 26435 32827 26441
rect 32769 26432 32781 26435
rect 32600 26404 32781 26432
rect 32769 26401 32781 26404
rect 32815 26401 32827 26435
rect 32769 26395 32827 26401
rect 23707 26336 23888 26364
rect 23707 26333 23719 26336
rect 23661 26327 23719 26333
rect 25682 26324 25688 26376
rect 25740 26373 25746 26376
rect 25740 26367 25763 26373
rect 25751 26333 25763 26367
rect 25740 26327 25763 26333
rect 25740 26324 25746 26327
rect 25866 26324 25872 26376
rect 25924 26324 25930 26376
rect 26050 26324 26056 26376
rect 26108 26364 26114 26376
rect 27246 26364 27252 26376
rect 26108 26336 27252 26364
rect 26108 26324 26114 26336
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 34514 26324 34520 26376
rect 34572 26364 34578 26376
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 34572 26336 34713 26364
rect 34572 26324 34578 26336
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 24121 26299 24179 26305
rect 24121 26296 24133 26299
rect 22020 26268 24133 26296
rect 18288 26200 19748 26228
rect 18288 26188 18294 26200
rect 20714 26188 20720 26240
rect 20772 26188 20778 26240
rect 21358 26188 21364 26240
rect 21416 26228 21422 26240
rect 21729 26231 21787 26237
rect 21729 26228 21741 26231
rect 21416 26200 21741 26228
rect 21416 26188 21422 26200
rect 21729 26197 21741 26200
rect 21775 26228 21787 26231
rect 22066 26228 22094 26268
rect 24121 26265 24133 26268
rect 24167 26265 24179 26299
rect 25961 26299 26019 26305
rect 24121 26259 24179 26265
rect 24228 26268 25912 26296
rect 21775 26200 22094 26228
rect 21775 26197 21787 26200
rect 21729 26191 21787 26197
rect 22186 26188 22192 26240
rect 22244 26228 22250 26240
rect 24228 26228 24256 26268
rect 22244 26200 24256 26228
rect 25884 26228 25912 26268
rect 25961 26265 25973 26299
rect 26007 26296 26019 26299
rect 26234 26296 26240 26308
rect 26007 26268 26240 26296
rect 26007 26265 26019 26268
rect 25961 26259 26019 26265
rect 26234 26256 26240 26268
rect 26292 26296 26298 26308
rect 27062 26296 27068 26308
rect 26292 26268 27068 26296
rect 26292 26256 26298 26268
rect 27062 26256 27068 26268
rect 27120 26256 27126 26308
rect 33042 26256 33048 26308
rect 33100 26256 33106 26308
rect 34793 26299 34851 26305
rect 34793 26296 34805 26299
rect 34270 26268 34805 26296
rect 34793 26265 34805 26268
rect 34839 26265 34851 26299
rect 34793 26259 34851 26265
rect 26326 26228 26332 26240
rect 25884 26200 26332 26228
rect 22244 26188 22250 26200
rect 26326 26188 26332 26200
rect 26384 26188 26390 26240
rect 30650 26188 30656 26240
rect 30708 26228 30714 26240
rect 31294 26228 31300 26240
rect 30708 26200 31300 26228
rect 30708 26188 30714 26200
rect 31294 26188 31300 26200
rect 31352 26188 31358 26240
rect 1104 26138 35236 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 35236 26138
rect 1104 26064 35236 26086
rect 12713 26027 12771 26033
rect 12713 25993 12725 26027
rect 12759 26024 12771 26027
rect 13354 26024 13360 26036
rect 12759 25996 13360 26024
rect 12759 25993 12771 25996
rect 12713 25987 12771 25993
rect 13354 25984 13360 25996
rect 13412 25984 13418 26036
rect 13722 26024 13728 26036
rect 13556 25996 13728 26024
rect 11241 25959 11299 25965
rect 11241 25925 11253 25959
rect 11287 25956 11299 25959
rect 11287 25928 11652 25956
rect 11287 25925 11299 25928
rect 11241 25919 11299 25925
rect 8665 25891 8723 25897
rect 8665 25857 8677 25891
rect 8711 25888 8723 25891
rect 9398 25888 9404 25900
rect 8711 25860 9404 25888
rect 8711 25857 8723 25860
rect 8665 25851 8723 25857
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 10413 25891 10471 25897
rect 10413 25888 10425 25891
rect 10284 25860 10425 25888
rect 10284 25848 10290 25860
rect 10413 25857 10425 25860
rect 10459 25888 10471 25891
rect 11057 25891 11115 25897
rect 11057 25888 11069 25891
rect 10459 25860 11069 25888
rect 10459 25857 10471 25860
rect 10413 25851 10471 25857
rect 11057 25857 11069 25860
rect 11103 25888 11115 25891
rect 11330 25888 11336 25900
rect 11103 25860 11336 25888
rect 11103 25857 11115 25860
rect 11057 25851 11115 25857
rect 11330 25848 11336 25860
rect 11388 25848 11394 25900
rect 11624 25897 11652 25928
rect 11974 25916 11980 25968
rect 12032 25956 12038 25968
rect 12345 25959 12403 25965
rect 12345 25956 12357 25959
rect 12032 25928 12357 25956
rect 12032 25916 12038 25928
rect 12345 25925 12357 25928
rect 12391 25925 12403 25959
rect 12345 25919 12403 25925
rect 12437 25959 12495 25965
rect 12437 25925 12449 25959
rect 12483 25956 12495 25959
rect 12897 25959 12955 25965
rect 12897 25956 12909 25959
rect 12483 25928 12909 25956
rect 12483 25925 12495 25928
rect 12437 25919 12495 25925
rect 12897 25925 12909 25928
rect 12943 25925 12955 25959
rect 12897 25919 12955 25925
rect 13556 25903 13584 25996
rect 13722 25984 13728 25996
rect 13780 25984 13786 26036
rect 16209 26027 16267 26033
rect 16209 26024 16221 26027
rect 15672 25996 16221 26024
rect 15672 25965 15700 25996
rect 16209 25993 16221 25996
rect 16255 26024 16267 26027
rect 16482 26024 16488 26036
rect 16255 25996 16488 26024
rect 16255 25993 16267 25996
rect 16209 25987 16267 25993
rect 16482 25984 16488 25996
rect 16540 25984 16546 26036
rect 16574 25984 16580 26036
rect 16632 26024 16638 26036
rect 16669 26027 16727 26033
rect 16669 26024 16681 26027
rect 16632 25996 16681 26024
rect 16632 25984 16638 25996
rect 16669 25993 16681 25996
rect 16715 25993 16727 26027
rect 16669 25987 16727 25993
rect 18049 26027 18107 26033
rect 18049 25993 18061 26027
rect 18095 26024 18107 26027
rect 18230 26024 18236 26036
rect 18095 25996 18236 26024
rect 18095 25993 18107 25996
rect 18049 25987 18107 25993
rect 18230 25984 18236 25996
rect 18288 25984 18294 26036
rect 19426 25984 19432 26036
rect 19484 25984 19490 26036
rect 21177 26027 21235 26033
rect 21177 25993 21189 26027
rect 21223 26024 21235 26027
rect 21266 26024 21272 26036
rect 21223 25996 21272 26024
rect 21223 25993 21235 25996
rect 21177 25987 21235 25993
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 27246 25984 27252 26036
rect 27304 25984 27310 26036
rect 29089 26027 29147 26033
rect 29089 25993 29101 26027
rect 29135 26024 29147 26027
rect 31573 26027 31631 26033
rect 29135 25996 29868 26024
rect 29135 25993 29147 25996
rect 29089 25987 29147 25993
rect 15657 25959 15715 25965
rect 13740 25928 14872 25956
rect 11517 25891 11575 25897
rect 11517 25857 11529 25891
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11609 25891 11667 25897
rect 11609 25857 11621 25891
rect 11655 25888 11667 25891
rect 11793 25891 11851 25897
rect 11655 25860 11744 25888
rect 11655 25857 11667 25860
rect 11609 25851 11667 25857
rect 10873 25823 10931 25829
rect 10873 25789 10885 25823
rect 10919 25789 10931 25823
rect 10873 25783 10931 25789
rect 9401 25755 9459 25761
rect 9401 25721 9413 25755
rect 9447 25752 9459 25755
rect 9447 25724 9904 25752
rect 9447 25721 9459 25724
rect 9401 25715 9459 25721
rect 9876 25696 9904 25724
rect 8846 25644 8852 25696
rect 8904 25684 8910 25696
rect 8941 25687 8999 25693
rect 8941 25684 8953 25687
rect 8904 25656 8953 25684
rect 8904 25644 8910 25656
rect 8941 25653 8953 25656
rect 8987 25653 8999 25687
rect 8941 25647 8999 25653
rect 9490 25644 9496 25696
rect 9548 25684 9554 25696
rect 9677 25687 9735 25693
rect 9677 25684 9689 25687
rect 9548 25656 9689 25684
rect 9548 25644 9554 25656
rect 9677 25653 9689 25656
rect 9723 25653 9735 25687
rect 9677 25647 9735 25653
rect 9858 25644 9864 25696
rect 9916 25684 9922 25696
rect 10781 25687 10839 25693
rect 10781 25684 10793 25687
rect 9916 25656 10793 25684
rect 9916 25644 9922 25656
rect 10781 25653 10793 25656
rect 10827 25684 10839 25687
rect 10888 25684 10916 25783
rect 11532 25752 11560 25851
rect 11716 25832 11744 25860
rect 11793 25857 11805 25891
rect 11839 25888 11851 25891
rect 12227 25891 12285 25897
rect 11839 25860 11928 25888
rect 11839 25857 11851 25860
rect 11793 25851 11851 25857
rect 11900 25832 11928 25860
rect 12227 25857 12239 25891
rect 12273 25857 12285 25891
rect 12227 25851 12285 25857
rect 11698 25780 11704 25832
rect 11756 25780 11762 25832
rect 11882 25780 11888 25832
rect 11940 25780 11946 25832
rect 11977 25823 12035 25829
rect 11977 25789 11989 25823
rect 12023 25820 12035 25823
rect 12069 25823 12127 25829
rect 12069 25820 12081 25823
rect 12023 25792 12081 25820
rect 12023 25789 12035 25792
rect 11977 25783 12035 25789
rect 12069 25789 12081 25792
rect 12115 25789 12127 25823
rect 12242 25820 12270 25851
rect 12526 25848 12532 25900
rect 12584 25848 12590 25900
rect 12802 25848 12808 25900
rect 12860 25848 12866 25900
rect 12986 25848 12992 25900
rect 13044 25848 13050 25900
rect 13446 25848 13452 25900
rect 13504 25848 13510 25900
rect 13538 25897 13596 25903
rect 13538 25863 13550 25897
rect 13584 25863 13596 25897
rect 13538 25857 13596 25863
rect 13630 25848 13636 25900
rect 13688 25848 13694 25900
rect 12710 25820 12716 25832
rect 12242 25792 12716 25820
rect 12069 25783 12127 25789
rect 12710 25780 12716 25792
rect 12768 25820 12774 25832
rect 13740 25820 13768 25928
rect 13814 25848 13820 25900
rect 13872 25848 13878 25900
rect 13909 25891 13967 25897
rect 13909 25857 13921 25891
rect 13955 25857 13967 25891
rect 13909 25851 13967 25857
rect 12768 25792 13768 25820
rect 13924 25820 13952 25851
rect 14090 25848 14096 25900
rect 14148 25848 14154 25900
rect 14844 25897 14872 25928
rect 15657 25925 15669 25959
rect 15703 25925 15715 25959
rect 15857 25959 15915 25965
rect 15857 25956 15869 25959
rect 15657 25919 15715 25925
rect 15764 25928 15869 25956
rect 14829 25891 14887 25897
rect 14829 25857 14841 25891
rect 14875 25857 14887 25891
rect 14829 25851 14887 25857
rect 15013 25891 15071 25897
rect 15013 25857 15025 25891
rect 15059 25888 15071 25891
rect 15059 25860 15148 25888
rect 15059 25857 15071 25860
rect 15013 25851 15071 25857
rect 15120 25829 15148 25860
rect 15562 25848 15568 25900
rect 15620 25848 15626 25900
rect 15105 25823 15163 25829
rect 13924 25792 14504 25820
rect 12768 25780 12774 25792
rect 12894 25752 12900 25764
rect 11532 25724 12900 25752
rect 12894 25712 12900 25724
rect 12952 25712 12958 25764
rect 13924 25752 13952 25792
rect 14476 25764 14504 25792
rect 15105 25789 15117 25823
rect 15151 25789 15163 25823
rect 15105 25783 15163 25789
rect 13004 25724 13952 25752
rect 13004 25684 13032 25724
rect 14458 25712 14464 25764
rect 14516 25712 14522 25764
rect 15672 25696 15700 25919
rect 15764 25900 15792 25928
rect 15857 25925 15869 25928
rect 15903 25925 15915 25959
rect 15857 25919 15915 25925
rect 16022 25916 16028 25968
rect 16080 25956 16086 25968
rect 17497 25959 17555 25965
rect 17497 25956 17509 25959
rect 16080 25928 17509 25956
rect 16080 25916 16086 25928
rect 15746 25848 15752 25900
rect 15804 25848 15810 25900
rect 16114 25848 16120 25900
rect 16172 25848 16178 25900
rect 16301 25891 16359 25897
rect 16301 25857 16313 25891
rect 16347 25888 16359 25891
rect 16390 25888 16396 25900
rect 16347 25860 16396 25888
rect 16347 25857 16359 25860
rect 16301 25851 16359 25857
rect 16390 25848 16396 25860
rect 16448 25848 16454 25900
rect 16868 25897 16896 25928
rect 17497 25925 17509 25928
rect 17543 25956 17555 25959
rect 17586 25956 17592 25968
rect 17543 25928 17592 25956
rect 17543 25925 17555 25928
rect 17497 25919 17555 25925
rect 17586 25916 17592 25928
rect 17644 25916 17650 25968
rect 18138 25956 18144 25968
rect 18064 25928 18144 25956
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25857 16911 25891
rect 16853 25851 16911 25857
rect 17034 25848 17040 25900
rect 17092 25848 17098 25900
rect 17126 25848 17132 25900
rect 17184 25848 17190 25900
rect 18064 25897 18092 25928
rect 18138 25916 18144 25928
rect 18196 25916 18202 25968
rect 19058 25956 19064 25968
rect 18892 25928 19064 25956
rect 18892 25897 18920 25928
rect 19058 25916 19064 25928
rect 19116 25956 19122 25968
rect 19116 25928 19288 25956
rect 19116 25916 19122 25928
rect 18049 25891 18107 25897
rect 18049 25857 18061 25891
rect 18095 25857 18107 25891
rect 18877 25891 18935 25897
rect 18877 25888 18889 25891
rect 18049 25851 18107 25857
rect 18156 25860 18889 25888
rect 16132 25752 16160 25848
rect 16206 25780 16212 25832
rect 16264 25820 16270 25832
rect 18156 25829 18184 25860
rect 18877 25857 18889 25860
rect 18923 25857 18935 25891
rect 18877 25851 18935 25857
rect 18969 25891 19027 25897
rect 18969 25857 18981 25891
rect 19015 25857 19027 25891
rect 18969 25851 19027 25857
rect 18141 25823 18199 25829
rect 18141 25820 18153 25823
rect 16264 25792 18153 25820
rect 16264 25780 16270 25792
rect 18141 25789 18153 25792
rect 18187 25789 18199 25823
rect 18141 25783 18199 25789
rect 18322 25780 18328 25832
rect 18380 25820 18386 25832
rect 18782 25820 18788 25832
rect 18380 25792 18788 25820
rect 18380 25780 18386 25792
rect 18782 25780 18788 25792
rect 18840 25820 18846 25832
rect 18984 25820 19012 25851
rect 19150 25848 19156 25900
rect 19208 25848 19214 25900
rect 19260 25888 19288 25928
rect 19334 25916 19340 25968
rect 19392 25916 19398 25968
rect 26326 25916 26332 25968
rect 26384 25916 26390 25968
rect 29457 25959 29515 25965
rect 29457 25925 29469 25959
rect 29503 25956 29515 25959
rect 29546 25956 29552 25968
rect 29503 25928 29552 25956
rect 29503 25925 29515 25928
rect 29457 25919 29515 25925
rect 29546 25916 29552 25928
rect 29604 25916 29610 25968
rect 29840 25965 29868 25996
rect 31573 25993 31585 26027
rect 31619 26024 31631 26027
rect 31662 26024 31668 26036
rect 31619 25996 31668 26024
rect 31619 25993 31631 25996
rect 31573 25987 31631 25993
rect 31662 25984 31668 25996
rect 31720 25984 31726 26036
rect 32677 26027 32735 26033
rect 32677 25993 32689 26027
rect 32723 26024 32735 26027
rect 33042 26024 33048 26036
rect 32723 25996 33048 26024
rect 32723 25993 32735 25996
rect 32677 25987 32735 25993
rect 33042 25984 33048 25996
rect 33100 25984 33106 26036
rect 29825 25959 29883 25965
rect 29825 25925 29837 25959
rect 29871 25925 29883 25959
rect 29825 25919 29883 25925
rect 30558 25916 30564 25968
rect 30616 25916 30622 25968
rect 19613 25891 19671 25897
rect 19613 25888 19625 25891
rect 19260 25860 19625 25888
rect 19613 25857 19625 25860
rect 19659 25857 19671 25891
rect 19613 25851 19671 25857
rect 20990 25848 20996 25900
rect 21048 25888 21054 25900
rect 21391 25891 21449 25897
rect 21391 25888 21403 25891
rect 21048 25860 21403 25888
rect 21048 25848 21054 25860
rect 21391 25857 21403 25860
rect 21437 25857 21449 25891
rect 21391 25851 21449 25857
rect 21545 25891 21603 25897
rect 21545 25857 21557 25891
rect 21591 25888 21603 25891
rect 26142 25888 26148 25900
rect 21591 25860 26148 25888
rect 21591 25857 21603 25860
rect 21545 25851 21603 25857
rect 26142 25848 26148 25860
rect 26200 25848 26206 25900
rect 18840 25792 19012 25820
rect 18840 25780 18846 25792
rect 16132 25724 16528 25752
rect 16500 25696 16528 25724
rect 16666 25712 16672 25764
rect 16724 25752 16730 25764
rect 16945 25755 17003 25761
rect 16945 25752 16957 25755
rect 16724 25724 16957 25752
rect 16724 25712 16730 25724
rect 16945 25721 16957 25724
rect 16991 25721 17003 25755
rect 18984 25752 19012 25792
rect 19242 25780 19248 25832
rect 19300 25780 19306 25832
rect 19797 25823 19855 25829
rect 19797 25789 19809 25823
rect 19843 25789 19855 25823
rect 26344 25820 26372 25916
rect 27154 25848 27160 25900
rect 27212 25888 27218 25900
rect 27525 25891 27583 25897
rect 27525 25888 27537 25891
rect 27212 25860 27537 25888
rect 27212 25848 27218 25860
rect 27525 25857 27537 25860
rect 27571 25888 27583 25891
rect 27801 25891 27859 25897
rect 27801 25888 27813 25891
rect 27571 25860 27813 25888
rect 27571 25857 27583 25860
rect 27525 25851 27583 25857
rect 27801 25857 27813 25860
rect 27847 25857 27859 25891
rect 27801 25851 27859 25857
rect 28721 25891 28779 25897
rect 28721 25857 28733 25891
rect 28767 25857 28779 25891
rect 28721 25851 28779 25857
rect 27249 25823 27307 25829
rect 27249 25820 27261 25823
rect 26344 25792 27261 25820
rect 19797 25783 19855 25789
rect 27249 25789 27261 25792
rect 27295 25820 27307 25823
rect 27338 25820 27344 25832
rect 27295 25792 27344 25820
rect 27295 25789 27307 25792
rect 27249 25783 27307 25789
rect 19812 25752 19840 25783
rect 27338 25780 27344 25792
rect 27396 25820 27402 25832
rect 27709 25823 27767 25829
rect 27709 25820 27721 25823
rect 27396 25792 27721 25820
rect 27396 25780 27402 25792
rect 27709 25789 27721 25792
rect 27755 25789 27767 25823
rect 27709 25783 27767 25789
rect 28169 25823 28227 25829
rect 28169 25789 28181 25823
rect 28215 25820 28227 25823
rect 28629 25823 28687 25829
rect 28629 25820 28641 25823
rect 28215 25792 28641 25820
rect 28215 25789 28227 25792
rect 28169 25783 28227 25789
rect 28629 25789 28641 25792
rect 28675 25789 28687 25823
rect 28629 25783 28687 25789
rect 23290 25752 23296 25764
rect 16945 25715 17003 25721
rect 17512 25724 18184 25752
rect 18984 25724 19840 25752
rect 23032 25724 23296 25752
rect 10827 25656 13032 25684
rect 10827 25653 10839 25656
rect 10781 25647 10839 25653
rect 13170 25644 13176 25696
rect 13228 25644 13234 25696
rect 13262 25644 13268 25696
rect 13320 25684 13326 25696
rect 13814 25684 13820 25696
rect 13320 25656 13820 25684
rect 13320 25644 13326 25656
rect 13814 25644 13820 25656
rect 13872 25684 13878 25696
rect 14001 25687 14059 25693
rect 14001 25684 14013 25687
rect 13872 25656 14013 25684
rect 13872 25644 13878 25656
rect 14001 25653 14013 25656
rect 14047 25653 14059 25687
rect 14001 25647 14059 25653
rect 14918 25644 14924 25696
rect 14976 25644 14982 25696
rect 15473 25687 15531 25693
rect 15473 25653 15485 25687
rect 15519 25684 15531 25687
rect 15654 25684 15660 25696
rect 15519 25656 15660 25684
rect 15519 25653 15531 25656
rect 15473 25647 15531 25653
rect 15654 25644 15660 25656
rect 15712 25644 15718 25696
rect 15841 25687 15899 25693
rect 15841 25653 15853 25687
rect 15887 25684 15899 25687
rect 15930 25684 15936 25696
rect 15887 25656 15936 25684
rect 15887 25653 15899 25656
rect 15841 25647 15899 25653
rect 15930 25644 15936 25656
rect 15988 25644 15994 25696
rect 16022 25644 16028 25696
rect 16080 25644 16086 25696
rect 16482 25644 16488 25696
rect 16540 25644 16546 25696
rect 16574 25644 16580 25696
rect 16632 25684 16638 25696
rect 17512 25684 17540 25724
rect 16632 25656 17540 25684
rect 18156 25684 18184 25724
rect 20533 25687 20591 25693
rect 20533 25684 20545 25687
rect 18156 25656 20545 25684
rect 16632 25644 16638 25656
rect 20533 25653 20545 25656
rect 20579 25684 20591 25687
rect 20898 25684 20904 25696
rect 20579 25656 20904 25684
rect 20579 25653 20591 25656
rect 20533 25647 20591 25653
rect 20898 25644 20904 25656
rect 20956 25644 20962 25696
rect 20993 25687 21051 25693
rect 20993 25653 21005 25687
rect 21039 25684 21051 25687
rect 21266 25684 21272 25696
rect 21039 25656 21272 25684
rect 21039 25653 21051 25656
rect 20993 25647 21051 25653
rect 21266 25644 21272 25656
rect 21324 25644 21330 25696
rect 22370 25644 22376 25696
rect 22428 25644 22434 25696
rect 22646 25644 22652 25696
rect 22704 25644 22710 25696
rect 22922 25644 22928 25696
rect 22980 25684 22986 25696
rect 23032 25693 23060 25724
rect 23290 25712 23296 25724
rect 23348 25752 23354 25764
rect 23753 25755 23811 25761
rect 23753 25752 23765 25755
rect 23348 25724 23765 25752
rect 23348 25712 23354 25724
rect 23753 25721 23765 25724
rect 23799 25721 23811 25755
rect 23753 25715 23811 25721
rect 27433 25755 27491 25761
rect 27433 25721 27445 25755
rect 27479 25752 27491 25755
rect 28074 25752 28080 25764
rect 27479 25724 28080 25752
rect 27479 25721 27491 25724
rect 27433 25715 27491 25721
rect 28074 25712 28080 25724
rect 28132 25752 28138 25764
rect 28736 25752 28764 25851
rect 29564 25829 29592 25916
rect 31941 25891 31999 25897
rect 31941 25888 31953 25891
rect 31772 25860 31953 25888
rect 29549 25823 29607 25829
rect 29549 25789 29561 25823
rect 29595 25789 29607 25823
rect 29549 25783 29607 25789
rect 31297 25823 31355 25829
rect 31297 25789 31309 25823
rect 31343 25820 31355 25823
rect 31343 25792 31708 25820
rect 31343 25789 31355 25792
rect 31297 25783 31355 25789
rect 28132 25724 28764 25752
rect 28132 25712 28138 25724
rect 23017 25687 23075 25693
rect 23017 25684 23029 25687
rect 22980 25656 23029 25684
rect 22980 25644 22986 25656
rect 23017 25653 23029 25656
rect 23063 25653 23075 25687
rect 23017 25647 23075 25653
rect 23382 25644 23388 25696
rect 23440 25644 23446 25696
rect 31680 25684 31708 25792
rect 31772 25764 31800 25860
rect 31941 25857 31953 25860
rect 31987 25857 31999 25891
rect 31941 25851 31999 25857
rect 32309 25891 32367 25897
rect 32309 25857 32321 25891
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 31846 25780 31852 25832
rect 31904 25780 31910 25832
rect 32214 25780 32220 25832
rect 32272 25780 32278 25832
rect 31754 25712 31760 25764
rect 31812 25712 31818 25764
rect 31941 25687 31999 25693
rect 31941 25684 31953 25687
rect 31680 25656 31953 25684
rect 31941 25653 31953 25656
rect 31987 25684 31999 25687
rect 32324 25684 32352 25851
rect 31987 25656 32352 25684
rect 31987 25653 31999 25656
rect 31941 25647 31999 25653
rect 34514 25644 34520 25696
rect 34572 25644 34578 25696
rect 1104 25594 35248 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 35248 25594
rect 1104 25520 35248 25542
rect 13170 25480 13176 25492
rect 11164 25452 13176 25480
rect 8389 25415 8447 25421
rect 8389 25381 8401 25415
rect 8435 25412 8447 25415
rect 9674 25412 9680 25424
rect 8435 25384 9680 25412
rect 8435 25381 8447 25384
rect 8389 25375 8447 25381
rect 9674 25372 9680 25384
rect 9732 25412 9738 25424
rect 9732 25384 10272 25412
rect 9732 25372 9738 25384
rect 9858 25304 9864 25356
rect 9916 25304 9922 25356
rect 10244 25288 10272 25384
rect 9309 25279 9367 25285
rect 9309 25245 9321 25279
rect 9355 25276 9367 25279
rect 9398 25276 9404 25288
rect 9355 25248 9404 25276
rect 9355 25245 9367 25248
rect 9309 25239 9367 25245
rect 9398 25236 9404 25248
rect 9456 25236 9462 25288
rect 9490 25236 9496 25288
rect 9548 25276 9554 25288
rect 10045 25279 10103 25285
rect 10045 25276 10057 25279
rect 9548 25248 10057 25276
rect 9548 25236 9554 25248
rect 10045 25245 10057 25248
rect 10091 25245 10103 25279
rect 10045 25239 10103 25245
rect 10226 25236 10232 25288
rect 10284 25236 10290 25288
rect 10965 25279 11023 25285
rect 10876 25257 10934 25263
rect 10876 25223 10888 25257
rect 10922 25223 10934 25257
rect 10965 25245 10977 25279
rect 11011 25276 11023 25279
rect 11054 25276 11060 25288
rect 11011 25248 11060 25276
rect 11011 25245 11023 25248
rect 10965 25239 11023 25245
rect 11054 25236 11060 25248
rect 11112 25236 11118 25288
rect 11164 25285 11192 25452
rect 13170 25440 13176 25452
rect 13228 25440 13234 25492
rect 13354 25440 13360 25492
rect 13412 25480 13418 25492
rect 13633 25483 13691 25489
rect 13633 25480 13645 25483
rect 13412 25452 13645 25480
rect 13412 25440 13418 25452
rect 13633 25449 13645 25452
rect 13679 25480 13691 25483
rect 13722 25480 13728 25492
rect 13679 25452 13728 25480
rect 13679 25449 13691 25452
rect 13633 25443 13691 25449
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 14090 25440 14096 25492
rect 14148 25480 14154 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 14148 25452 14289 25480
rect 14148 25440 14154 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 14918 25440 14924 25492
rect 14976 25440 14982 25492
rect 15013 25483 15071 25489
rect 15013 25449 15025 25483
rect 15059 25480 15071 25483
rect 15838 25480 15844 25492
rect 15059 25452 15844 25480
rect 15059 25449 15071 25452
rect 15013 25443 15071 25449
rect 15838 25440 15844 25452
rect 15896 25440 15902 25492
rect 16574 25480 16580 25492
rect 15948 25452 16580 25480
rect 11698 25372 11704 25424
rect 11756 25412 11762 25424
rect 11756 25384 12434 25412
rect 11756 25372 11762 25384
rect 11333 25347 11391 25353
rect 11333 25344 11345 25347
rect 11256 25316 11345 25344
rect 11256 25285 11284 25316
rect 11333 25313 11345 25316
rect 11379 25313 11391 25347
rect 11716 25344 11744 25372
rect 11333 25307 11391 25313
rect 11624 25316 11744 25344
rect 11624 25285 11652 25316
rect 11882 25304 11888 25356
rect 11940 25344 11946 25356
rect 12406 25344 12434 25384
rect 12802 25372 12808 25424
rect 12860 25372 12866 25424
rect 12820 25344 12848 25372
rect 11940 25316 12296 25344
rect 12406 25316 12848 25344
rect 11940 25304 11946 25316
rect 11149 25279 11207 25285
rect 11149 25245 11161 25279
rect 11195 25245 11207 25279
rect 11149 25239 11207 25245
rect 11241 25279 11299 25285
rect 11241 25245 11253 25279
rect 11287 25245 11299 25279
rect 11241 25239 11299 25245
rect 11609 25279 11667 25285
rect 11609 25245 11621 25279
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 11698 25236 11704 25288
rect 11756 25236 11762 25288
rect 11793 25279 11851 25285
rect 11793 25245 11805 25279
rect 11839 25276 11851 25279
rect 11900 25276 11928 25304
rect 12268 25285 12296 25316
rect 11839 25248 11928 25276
rect 11839 25245 11851 25248
rect 11793 25239 11851 25245
rect 10876 25220 10934 25223
rect 9030 25168 9036 25220
rect 9088 25208 9094 25220
rect 9585 25211 9643 25217
rect 9585 25208 9597 25211
rect 9088 25180 9597 25208
rect 9088 25168 9094 25180
rect 9585 25177 9597 25180
rect 9631 25177 9643 25211
rect 9585 25171 9643 25177
rect 10410 25168 10416 25220
rect 10468 25208 10474 25220
rect 10870 25208 10876 25220
rect 10468 25180 10876 25208
rect 10468 25168 10474 25180
rect 10870 25168 10876 25180
rect 10928 25168 10934 25220
rect 11330 25168 11336 25220
rect 11388 25208 11394 25220
rect 11900 25208 11928 25248
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25245 12035 25279
rect 11977 25239 12035 25245
rect 12253 25279 12311 25285
rect 12253 25245 12265 25279
rect 12299 25245 12311 25279
rect 12253 25239 12311 25245
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25245 12403 25279
rect 12345 25239 12403 25245
rect 12529 25279 12587 25285
rect 12529 25245 12541 25279
rect 12575 25245 12587 25279
rect 12529 25239 12587 25245
rect 12621 25279 12679 25285
rect 12621 25245 12633 25279
rect 12667 25276 12679 25279
rect 12820 25276 12848 25316
rect 12667 25248 12848 25276
rect 12667 25245 12679 25248
rect 12621 25239 12679 25245
rect 11388 25180 11928 25208
rect 11992 25208 12020 25239
rect 12360 25208 12388 25239
rect 11992 25180 12388 25208
rect 12544 25208 12572 25239
rect 12986 25236 12992 25288
rect 13044 25236 13050 25288
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 13173 25279 13231 25285
rect 13173 25245 13185 25279
rect 13219 25276 13231 25279
rect 13262 25276 13268 25288
rect 13219 25248 13268 25276
rect 13219 25245 13231 25248
rect 13173 25239 13231 25245
rect 13004 25208 13032 25236
rect 12544 25180 13032 25208
rect 13096 25208 13124 25239
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 13372 25285 13400 25440
rect 13446 25372 13452 25424
rect 13504 25412 13510 25424
rect 13906 25412 13912 25424
rect 13504 25384 13912 25412
rect 13504 25372 13517 25384
rect 13906 25372 13912 25384
rect 13964 25412 13970 25424
rect 13964 25384 14136 25412
rect 13964 25372 13970 25384
rect 13489 25344 13517 25372
rect 13464 25316 13517 25344
rect 13648 25316 13860 25344
rect 13464 25285 13492 25316
rect 13357 25279 13415 25285
rect 13357 25245 13369 25279
rect 13403 25245 13415 25279
rect 13357 25239 13415 25245
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25245 13507 25279
rect 13449 25239 13507 25245
rect 13541 25279 13599 25285
rect 13541 25245 13553 25279
rect 13587 25276 13599 25279
rect 13648 25276 13676 25316
rect 13587 25248 13676 25276
rect 13725 25279 13783 25285
rect 13587 25245 13599 25248
rect 13541 25239 13599 25245
rect 13725 25245 13737 25279
rect 13771 25245 13783 25279
rect 13725 25239 13783 25245
rect 13630 25208 13636 25220
rect 13096 25180 13636 25208
rect 11388 25168 11394 25180
rect 12268 25152 12296 25180
rect 8757 25143 8815 25149
rect 8757 25109 8769 25143
rect 8803 25140 8815 25143
rect 8846 25140 8852 25152
rect 8803 25112 8852 25140
rect 8803 25109 8815 25112
rect 8757 25103 8815 25109
rect 8846 25100 8852 25112
rect 8904 25140 8910 25152
rect 10137 25143 10195 25149
rect 10137 25140 10149 25143
rect 8904 25112 10149 25140
rect 8904 25100 8910 25112
rect 10137 25109 10149 25112
rect 10183 25140 10195 25143
rect 10502 25140 10508 25152
rect 10183 25112 10508 25140
rect 10183 25109 10195 25112
rect 10137 25103 10195 25109
rect 10502 25100 10508 25112
rect 10560 25100 10566 25152
rect 10689 25143 10747 25149
rect 10689 25109 10701 25143
rect 10735 25140 10747 25143
rect 11238 25140 11244 25152
rect 10735 25112 11244 25140
rect 10735 25109 10747 25112
rect 10689 25103 10747 25109
rect 11238 25100 11244 25112
rect 11296 25100 11302 25152
rect 12066 25100 12072 25152
rect 12124 25100 12130 25152
rect 12250 25100 12256 25152
rect 12308 25100 12314 25152
rect 12342 25100 12348 25152
rect 12400 25140 12406 25152
rect 12544 25140 12572 25180
rect 12400 25112 12572 25140
rect 12400 25100 12406 25112
rect 12802 25100 12808 25152
rect 12860 25140 12866 25152
rect 12897 25143 12955 25149
rect 12897 25140 12909 25143
rect 12860 25112 12909 25140
rect 12860 25100 12866 25112
rect 12897 25109 12909 25112
rect 12943 25109 12955 25143
rect 12897 25103 12955 25109
rect 12986 25100 12992 25152
rect 13044 25140 13050 25152
rect 13096 25140 13124 25180
rect 13630 25168 13636 25180
rect 13688 25168 13694 25220
rect 13740 25152 13768 25239
rect 13832 25208 13860 25316
rect 14108 25288 14136 25384
rect 14936 25344 14964 25440
rect 15948 25412 15976 25452
rect 16574 25440 16580 25452
rect 16632 25440 16638 25492
rect 16669 25483 16727 25489
rect 16669 25449 16681 25483
rect 16715 25480 16727 25483
rect 17034 25480 17040 25492
rect 16715 25452 17040 25480
rect 16715 25449 16727 25452
rect 16669 25443 16727 25449
rect 17034 25440 17040 25452
rect 17092 25440 17098 25492
rect 23017 25483 23075 25489
rect 23017 25449 23029 25483
rect 23063 25480 23075 25483
rect 23658 25480 23664 25492
rect 23063 25452 23664 25480
rect 23063 25449 23075 25452
rect 23017 25443 23075 25449
rect 23658 25440 23664 25452
rect 23716 25440 23722 25492
rect 23750 25440 23756 25492
rect 23808 25440 23814 25492
rect 24854 25440 24860 25492
rect 24912 25440 24918 25492
rect 30558 25440 30564 25492
rect 30616 25440 30622 25492
rect 32033 25483 32091 25489
rect 32033 25449 32045 25483
rect 32079 25480 32091 25483
rect 32214 25480 32220 25492
rect 32079 25452 32220 25480
rect 32079 25449 32091 25452
rect 32033 25443 32091 25449
rect 32214 25440 32220 25452
rect 32272 25440 32278 25492
rect 15488 25384 15976 25412
rect 15151 25347 15209 25353
rect 15151 25344 15163 25347
rect 14936 25316 15163 25344
rect 15151 25313 15163 25316
rect 15197 25313 15209 25347
rect 15151 25307 15209 25313
rect 14090 25236 14096 25288
rect 14148 25236 14154 25288
rect 15286 25236 15292 25288
rect 15344 25236 15350 25288
rect 15488 25208 15516 25384
rect 16114 25372 16120 25424
rect 16172 25412 16178 25424
rect 16172 25384 16804 25412
rect 16172 25372 16178 25384
rect 15562 25304 15568 25356
rect 15620 25304 15626 25356
rect 16206 25304 16212 25356
rect 16264 25304 16270 25356
rect 16298 25304 16304 25356
rect 16356 25344 16362 25356
rect 16666 25344 16672 25356
rect 16356 25316 16672 25344
rect 16356 25304 16362 25316
rect 16666 25304 16672 25316
rect 16724 25304 16730 25356
rect 15746 25236 15752 25288
rect 15804 25276 15810 25288
rect 16117 25279 16175 25285
rect 15804 25248 15976 25276
rect 15804 25236 15810 25248
rect 13832 25180 15516 25208
rect 15657 25211 15715 25217
rect 13832 25152 13860 25180
rect 15657 25177 15669 25211
rect 15703 25208 15715 25211
rect 15948 25208 15976 25248
rect 16117 25245 16129 25279
rect 16163 25276 16175 25279
rect 16224 25276 16252 25304
rect 16776 25285 16804 25384
rect 20714 25372 20720 25424
rect 20772 25412 20778 25424
rect 21085 25415 21143 25421
rect 21085 25412 21097 25415
rect 20772 25384 21097 25412
rect 20772 25372 20778 25384
rect 16163 25248 16252 25276
rect 16577 25279 16635 25285
rect 16163 25245 16175 25248
rect 16117 25239 16175 25245
rect 16577 25245 16589 25279
rect 16623 25245 16635 25279
rect 16577 25239 16635 25245
rect 16761 25279 16819 25285
rect 16761 25245 16773 25279
rect 16807 25245 16819 25279
rect 16761 25239 16819 25245
rect 16592 25208 16620 25239
rect 15703 25180 15792 25208
rect 15948 25180 16620 25208
rect 20824 25208 20852 25384
rect 21085 25381 21097 25384
rect 21131 25381 21143 25415
rect 22646 25412 22652 25424
rect 21085 25375 21143 25381
rect 21376 25384 22652 25412
rect 20898 25236 20904 25288
rect 20956 25276 20962 25288
rect 21376 25285 21404 25384
rect 22646 25372 22652 25384
rect 22704 25372 22710 25424
rect 23290 25412 23296 25424
rect 22848 25384 23296 25412
rect 21818 25304 21824 25356
rect 21876 25304 21882 25356
rect 22557 25347 22615 25353
rect 22557 25344 22569 25347
rect 22066 25316 22569 25344
rect 21361 25279 21419 25285
rect 21361 25276 21373 25279
rect 20956 25248 21373 25276
rect 20956 25236 20962 25248
rect 21361 25245 21373 25248
rect 21407 25245 21419 25279
rect 21361 25239 21419 25245
rect 21637 25279 21695 25285
rect 21637 25245 21649 25279
rect 21683 25276 21695 25279
rect 21913 25279 21971 25285
rect 21913 25276 21925 25279
rect 21683 25248 21925 25276
rect 21683 25245 21695 25248
rect 21637 25239 21695 25245
rect 21913 25245 21925 25248
rect 21959 25245 21971 25279
rect 21913 25239 21971 25245
rect 22066 25208 22094 25316
rect 22557 25313 22569 25316
rect 22603 25344 22615 25347
rect 22848 25344 22876 25384
rect 23290 25372 23296 25384
rect 23348 25372 23354 25424
rect 22603 25316 22876 25344
rect 22940 25316 23428 25344
rect 22603 25313 22615 25316
rect 22557 25307 22615 25313
rect 22940 25288 22968 25316
rect 22922 25236 22928 25288
rect 22980 25236 22986 25288
rect 23198 25236 23204 25288
rect 23256 25236 23262 25288
rect 23400 25285 23428 25316
rect 24762 25304 24768 25356
rect 24820 25344 24826 25356
rect 24949 25347 25007 25353
rect 24949 25344 24961 25347
rect 24820 25316 24961 25344
rect 24820 25304 24826 25316
rect 24949 25313 24961 25316
rect 24995 25313 25007 25347
rect 24949 25307 25007 25313
rect 26142 25304 26148 25356
rect 26200 25304 26206 25356
rect 27338 25304 27344 25356
rect 27396 25344 27402 25356
rect 27525 25347 27583 25353
rect 27525 25344 27537 25347
rect 27396 25316 27537 25344
rect 27396 25304 27402 25316
rect 27525 25313 27537 25316
rect 27571 25313 27583 25347
rect 31941 25347 31999 25353
rect 31941 25344 31953 25347
rect 27525 25307 27583 25313
rect 31772 25316 31953 25344
rect 23385 25279 23443 25285
rect 23385 25245 23397 25279
rect 23431 25245 23443 25279
rect 23385 25239 23443 25245
rect 23658 25236 23664 25288
rect 23716 25236 23722 25288
rect 23937 25279 23995 25285
rect 23937 25245 23949 25279
rect 23983 25245 23995 25279
rect 23937 25239 23995 25245
rect 20824 25180 22094 25208
rect 22296 25180 23244 25208
rect 15703 25177 15715 25180
rect 15657 25171 15715 25177
rect 13044 25112 13124 25140
rect 13044 25100 13050 25112
rect 13722 25100 13728 25152
rect 13780 25100 13786 25152
rect 13814 25100 13820 25152
rect 13872 25100 13878 25152
rect 15764 25149 15792 25180
rect 15749 25143 15807 25149
rect 15749 25109 15761 25143
rect 15795 25109 15807 25143
rect 15749 25103 15807 25109
rect 16206 25100 16212 25152
rect 16264 25100 16270 25152
rect 20070 25100 20076 25152
rect 20128 25100 20134 25152
rect 20438 25100 20444 25152
rect 20496 25100 20502 25152
rect 20806 25100 20812 25152
rect 20864 25100 20870 25152
rect 21266 25100 21272 25152
rect 21324 25100 21330 25152
rect 21453 25143 21511 25149
rect 21453 25109 21465 25143
rect 21499 25140 21511 25143
rect 21726 25140 21732 25152
rect 21499 25112 21732 25140
rect 21499 25109 21511 25112
rect 21453 25103 21511 25109
rect 21726 25100 21732 25112
rect 21784 25100 21790 25152
rect 22296 25149 22324 25180
rect 22281 25143 22339 25149
rect 22281 25109 22293 25143
rect 22327 25109 22339 25143
rect 23216 25140 23244 25180
rect 23290 25168 23296 25220
rect 23348 25168 23354 25220
rect 23523 25211 23581 25217
rect 23523 25177 23535 25211
rect 23569 25208 23581 25211
rect 23952 25208 23980 25239
rect 24026 25236 24032 25288
rect 24084 25236 24090 25288
rect 24394 25236 24400 25288
rect 24452 25236 24458 25288
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25276 24731 25279
rect 24854 25276 24860 25288
rect 24719 25248 24860 25276
rect 24719 25245 24731 25248
rect 24673 25239 24731 25245
rect 24688 25208 24716 25239
rect 24854 25236 24860 25248
rect 24912 25236 24918 25288
rect 25774 25236 25780 25288
rect 25832 25236 25838 25288
rect 25958 25236 25964 25288
rect 26016 25236 26022 25288
rect 26160 25276 26188 25304
rect 31772 25288 31800 25316
rect 31941 25313 31953 25316
rect 31987 25313 31999 25347
rect 31941 25307 31999 25313
rect 32125 25347 32183 25353
rect 32125 25313 32137 25347
rect 32171 25344 32183 25347
rect 32306 25344 32312 25356
rect 32171 25316 32312 25344
rect 32171 25313 32183 25316
rect 32125 25307 32183 25313
rect 32306 25304 32312 25316
rect 32364 25344 32370 25356
rect 34057 25347 34115 25353
rect 32364 25316 32996 25344
rect 32364 25304 32370 25316
rect 32968 25288 32996 25316
rect 34057 25313 34069 25347
rect 34103 25313 34115 25347
rect 34057 25307 34115 25313
rect 27614 25276 27620 25288
rect 26160 25248 27620 25276
rect 27614 25236 27620 25248
rect 27672 25236 27678 25288
rect 27709 25279 27767 25285
rect 27709 25245 27721 25279
rect 27755 25276 27767 25279
rect 27798 25276 27804 25288
rect 27755 25248 27804 25276
rect 27755 25245 27767 25248
rect 27709 25239 27767 25245
rect 27798 25236 27804 25248
rect 27856 25236 27862 25288
rect 30469 25279 30527 25285
rect 30469 25245 30481 25279
rect 30515 25245 30527 25279
rect 30469 25239 30527 25245
rect 23569 25180 24716 25208
rect 23569 25177 23581 25180
rect 23523 25171 23581 25177
rect 24302 25140 24308 25152
rect 23216 25112 24308 25140
rect 22281 25103 22339 25109
rect 24302 25100 24308 25112
rect 24360 25140 24366 25152
rect 24489 25143 24547 25149
rect 24489 25140 24501 25143
rect 24360 25112 24501 25140
rect 24360 25100 24366 25112
rect 24489 25109 24501 25112
rect 24535 25109 24547 25143
rect 24489 25103 24547 25109
rect 27338 25100 27344 25152
rect 27396 25100 27402 25152
rect 30377 25143 30435 25149
rect 30377 25109 30389 25143
rect 30423 25140 30435 25143
rect 30484 25140 30512 25239
rect 31754 25236 31760 25288
rect 31812 25236 31818 25288
rect 31846 25236 31852 25288
rect 31904 25236 31910 25288
rect 32950 25236 32956 25288
rect 33008 25236 33014 25288
rect 31864 25208 31892 25236
rect 34072 25220 34100 25307
rect 34517 25279 34575 25285
rect 34517 25245 34529 25279
rect 34563 25276 34575 25279
rect 34882 25276 34888 25288
rect 34563 25248 34888 25276
rect 34563 25245 34575 25248
rect 34517 25239 34575 25245
rect 34882 25236 34888 25248
rect 34940 25236 34946 25288
rect 31864 25180 31984 25208
rect 31956 25152 31984 25180
rect 34054 25168 34060 25220
rect 34112 25168 34118 25220
rect 30650 25140 30656 25152
rect 30423 25112 30656 25140
rect 30423 25109 30435 25112
rect 30377 25103 30435 25109
rect 30650 25100 30656 25112
rect 30708 25100 30714 25152
rect 31938 25100 31944 25152
rect 31996 25100 32002 25152
rect 1104 25050 35236 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 35236 25050
rect 1104 24976 35236 24998
rect 9398 24896 9404 24948
rect 9456 24896 9462 24948
rect 11330 24896 11336 24948
rect 11388 24896 11394 24948
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 12342 24936 12348 24948
rect 11756 24908 12348 24936
rect 11756 24896 11762 24908
rect 12342 24896 12348 24908
rect 12400 24896 12406 24948
rect 15654 24896 15660 24948
rect 15712 24896 15718 24948
rect 15933 24939 15991 24945
rect 15933 24905 15945 24939
rect 15979 24936 15991 24939
rect 16206 24936 16212 24948
rect 15979 24908 16212 24936
rect 15979 24905 15991 24908
rect 15933 24899 15991 24905
rect 16206 24896 16212 24908
rect 16264 24896 16270 24948
rect 20806 24896 20812 24948
rect 20864 24936 20870 24948
rect 21361 24939 21419 24945
rect 21361 24936 21373 24939
rect 20864 24908 21373 24936
rect 20864 24896 20870 24908
rect 21361 24905 21373 24908
rect 21407 24905 21419 24939
rect 21361 24899 21419 24905
rect 21637 24939 21695 24945
rect 21637 24905 21649 24939
rect 21683 24936 21695 24939
rect 21818 24936 21824 24948
rect 21683 24908 21824 24936
rect 21683 24905 21695 24908
rect 21637 24899 21695 24905
rect 8846 24868 8852 24880
rect 8680 24840 8852 24868
rect 8021 24803 8079 24809
rect 8021 24769 8033 24803
rect 8067 24800 8079 24803
rect 8205 24803 8263 24809
rect 8205 24800 8217 24803
rect 8067 24772 8217 24800
rect 8067 24769 8079 24772
rect 8021 24763 8079 24769
rect 8205 24769 8217 24772
rect 8251 24800 8263 24803
rect 8570 24800 8576 24812
rect 8251 24772 8576 24800
rect 8251 24769 8263 24772
rect 8205 24763 8263 24769
rect 8570 24760 8576 24772
rect 8628 24760 8634 24812
rect 8680 24809 8708 24840
rect 8846 24828 8852 24840
rect 8904 24828 8910 24880
rect 9416 24868 9444 24896
rect 8956 24840 9168 24868
rect 9416 24840 9628 24868
rect 8665 24803 8723 24809
rect 8665 24769 8677 24803
rect 8711 24769 8723 24803
rect 8956 24800 8984 24840
rect 8665 24763 8723 24769
rect 8772 24772 8984 24800
rect 8772 24673 8800 24772
rect 9030 24760 9036 24812
rect 9088 24760 9094 24812
rect 9140 24800 9168 24840
rect 9214 24800 9220 24812
rect 9140 24772 9220 24800
rect 9214 24760 9220 24772
rect 9272 24800 9278 24812
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 9272 24772 9413 24800
rect 9272 24760 9278 24772
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 9600 24800 9628 24840
rect 10520 24840 11192 24868
rect 10520 24800 10548 24840
rect 11164 24809 11192 24840
rect 12434 24828 12440 24880
rect 12492 24868 12498 24880
rect 15672 24868 15700 24896
rect 20717 24871 20775 24877
rect 12492 24840 13860 24868
rect 15672 24840 16068 24868
rect 12492 24828 12498 24840
rect 9600 24772 10548 24800
rect 11149 24803 11207 24809
rect 9401 24763 9459 24769
rect 11149 24769 11161 24803
rect 11195 24800 11207 24803
rect 12069 24803 12127 24809
rect 12069 24800 12081 24803
rect 11195 24772 12081 24800
rect 11195 24769 11207 24772
rect 11149 24763 11207 24769
rect 12069 24769 12081 24772
rect 12115 24800 12127 24803
rect 13722 24800 13728 24812
rect 12115 24772 13728 24800
rect 12115 24769 12127 24772
rect 12069 24763 12127 24769
rect 13722 24760 13728 24772
rect 13780 24760 13786 24812
rect 13832 24744 13860 24840
rect 15654 24800 15660 24812
rect 15212 24772 15660 24800
rect 15212 24744 15240 24772
rect 15654 24760 15660 24772
rect 15712 24760 15718 24812
rect 15749 24803 15807 24809
rect 15749 24769 15761 24803
rect 15795 24800 15807 24803
rect 15930 24800 15936 24812
rect 15795 24772 15936 24800
rect 15795 24769 15807 24772
rect 15749 24763 15807 24769
rect 10965 24735 11023 24741
rect 10965 24732 10977 24735
rect 10244 24704 10977 24732
rect 8757 24667 8815 24673
rect 8757 24633 8769 24667
rect 8803 24633 8815 24667
rect 8757 24627 8815 24633
rect 8846 24624 8852 24676
rect 8904 24664 8910 24676
rect 10244 24664 10272 24704
rect 10965 24701 10977 24704
rect 11011 24701 11023 24735
rect 10965 24695 11023 24701
rect 13449 24735 13507 24741
rect 13449 24701 13461 24735
rect 13495 24732 13507 24735
rect 13814 24732 13820 24744
rect 13495 24704 13820 24732
rect 13495 24701 13507 24704
rect 13449 24695 13507 24701
rect 8904 24636 10272 24664
rect 8904 24624 8910 24636
rect 10689 24599 10747 24605
rect 10689 24565 10701 24599
rect 10735 24596 10747 24599
rect 10778 24596 10784 24608
rect 10735 24568 10784 24596
rect 10735 24565 10747 24568
rect 10689 24559 10747 24565
rect 10778 24556 10784 24568
rect 10836 24556 10842 24608
rect 10980 24596 11008 24695
rect 13814 24692 13820 24704
rect 13872 24692 13878 24744
rect 15194 24692 15200 24744
rect 15252 24692 15258 24744
rect 15764 24676 15792 24763
rect 15930 24760 15936 24772
rect 15988 24760 15994 24812
rect 16040 24809 16068 24840
rect 20717 24837 20729 24871
rect 20763 24868 20775 24871
rect 20990 24868 20996 24880
rect 20763 24840 20996 24868
rect 20763 24837 20775 24840
rect 20717 24831 20775 24837
rect 20990 24828 20996 24840
rect 21048 24828 21054 24880
rect 21082 24828 21088 24880
rect 21140 24868 21146 24880
rect 21269 24871 21327 24877
rect 21269 24868 21281 24871
rect 21140 24840 21281 24868
rect 21140 24828 21146 24840
rect 21269 24837 21281 24840
rect 21315 24837 21327 24871
rect 21376 24868 21404 24899
rect 21818 24896 21824 24908
rect 21876 24896 21882 24948
rect 22370 24896 22376 24948
rect 22428 24936 22434 24948
rect 22833 24939 22891 24945
rect 22833 24936 22845 24939
rect 22428 24908 22845 24936
rect 22428 24896 22434 24908
rect 22833 24905 22845 24908
rect 22879 24905 22891 24939
rect 22833 24899 22891 24905
rect 23198 24896 23204 24948
rect 23256 24936 23262 24948
rect 23293 24939 23351 24945
rect 23293 24936 23305 24939
rect 23256 24908 23305 24936
rect 23256 24896 23262 24908
rect 23293 24905 23305 24908
rect 23339 24905 23351 24939
rect 23293 24899 23351 24905
rect 23750 24896 23756 24948
rect 23808 24896 23814 24948
rect 24854 24896 24860 24948
rect 24912 24896 24918 24948
rect 25148 24908 25820 24936
rect 22462 24868 22468 24880
rect 21376 24840 22468 24868
rect 21269 24831 21327 24837
rect 22462 24828 22468 24840
rect 22520 24828 22526 24880
rect 22646 24828 22652 24880
rect 22704 24828 22710 24880
rect 22925 24871 22983 24877
rect 22925 24837 22937 24871
rect 22971 24868 22983 24871
rect 23768 24868 23796 24896
rect 22971 24840 23152 24868
rect 22971 24837 22983 24840
rect 22925 24831 22983 24837
rect 16025 24803 16083 24809
rect 16025 24769 16037 24803
rect 16071 24769 16083 24803
rect 16025 24763 16083 24769
rect 18322 24760 18328 24812
rect 18380 24800 18386 24812
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 18380 24772 19165 24800
rect 18380 24760 18386 24772
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19153 24763 19211 24769
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19978 24800 19984 24812
rect 19392 24772 19984 24800
rect 19392 24760 19398 24772
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20438 24760 20444 24812
rect 20496 24800 20502 24812
rect 21453 24803 21511 24809
rect 21453 24800 21465 24803
rect 20496 24772 21465 24800
rect 20496 24760 20502 24772
rect 21453 24769 21465 24772
rect 21499 24800 21511 24803
rect 23017 24803 23075 24809
rect 23017 24800 23029 24803
rect 21499 24772 23029 24800
rect 21499 24769 21511 24772
rect 21453 24763 21511 24769
rect 15838 24692 15844 24744
rect 15896 24692 15902 24744
rect 19058 24692 19064 24744
rect 19116 24692 19122 24744
rect 19521 24735 19579 24741
rect 19521 24701 19533 24735
rect 19567 24732 19579 24735
rect 19797 24735 19855 24741
rect 19797 24732 19809 24735
rect 19567 24704 19809 24732
rect 19567 24701 19579 24704
rect 19521 24695 19579 24701
rect 19797 24701 19809 24704
rect 19843 24701 19855 24735
rect 19797 24695 19855 24701
rect 22112 24676 22140 24772
rect 23017 24769 23029 24772
rect 23063 24769 23075 24803
rect 23017 24763 23075 24769
rect 11054 24624 11060 24676
rect 11112 24664 11118 24676
rect 13078 24664 13084 24676
rect 11112 24636 13084 24664
rect 11112 24624 11118 24636
rect 13078 24624 13084 24636
rect 13136 24624 13142 24676
rect 15378 24664 15384 24676
rect 13280 24636 15384 24664
rect 11793 24599 11851 24605
rect 11793 24596 11805 24599
rect 10980 24568 11805 24596
rect 11793 24565 11805 24568
rect 11839 24596 11851 24599
rect 12434 24596 12440 24608
rect 11839 24568 12440 24596
rect 11839 24565 11851 24568
rect 11793 24559 11851 24565
rect 12434 24556 12440 24568
rect 12492 24556 12498 24608
rect 12710 24556 12716 24608
rect 12768 24596 12774 24608
rect 13280 24596 13308 24636
rect 15378 24624 15384 24636
rect 15436 24624 15442 24676
rect 15746 24624 15752 24676
rect 15804 24624 15810 24676
rect 16390 24624 16396 24676
rect 16448 24624 16454 24676
rect 16482 24624 16488 24676
rect 16540 24664 16546 24676
rect 17954 24664 17960 24676
rect 16540 24636 17960 24664
rect 16540 24624 16546 24636
rect 17954 24624 17960 24636
rect 18012 24664 18018 24676
rect 21085 24667 21143 24673
rect 21085 24664 21097 24667
rect 18012 24636 21097 24664
rect 18012 24624 18018 24636
rect 21085 24633 21097 24636
rect 21131 24664 21143 24667
rect 21358 24664 21364 24676
rect 21131 24636 21364 24664
rect 21131 24633 21143 24636
rect 21085 24627 21143 24633
rect 21358 24624 21364 24636
rect 21416 24624 21422 24676
rect 22094 24624 22100 24676
rect 22152 24624 22158 24676
rect 12768 24568 13308 24596
rect 12768 24556 12774 24568
rect 13722 24556 13728 24608
rect 13780 24596 13786 24608
rect 13817 24599 13875 24605
rect 13817 24596 13829 24599
rect 13780 24568 13829 24596
rect 13780 24556 13786 24568
rect 13817 24565 13829 24568
rect 13863 24596 13875 24599
rect 16408 24596 16436 24624
rect 13863 24568 16436 24596
rect 13863 24565 13875 24568
rect 13817 24559 13875 24565
rect 22462 24556 22468 24608
rect 22520 24596 22526 24608
rect 23124 24596 23152 24840
rect 23492 24840 23796 24868
rect 24673 24871 24731 24877
rect 23492 24809 23520 24840
rect 24673 24837 24685 24871
rect 24719 24868 24731 24871
rect 25148 24868 25176 24908
rect 25792 24880 25820 24908
rect 29638 24896 29644 24948
rect 29696 24896 29702 24948
rect 34882 24896 34888 24948
rect 34940 24896 34946 24948
rect 24719 24840 25176 24868
rect 25240 24840 25452 24868
rect 24719 24837 24731 24840
rect 24673 24831 24731 24837
rect 23477 24803 23535 24809
rect 23477 24769 23489 24803
rect 23523 24769 23535 24803
rect 23477 24763 23535 24769
rect 23750 24760 23756 24812
rect 23808 24760 23814 24812
rect 23937 24803 23995 24809
rect 23937 24769 23949 24803
rect 23983 24800 23995 24803
rect 24026 24800 24032 24812
rect 23983 24772 24032 24800
rect 23983 24769 23995 24772
rect 23937 24763 23995 24769
rect 23201 24735 23259 24741
rect 23201 24701 23213 24735
rect 23247 24732 23259 24735
rect 23952 24732 23980 24763
rect 24026 24760 24032 24772
rect 24084 24760 24090 24812
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 23247 24704 23980 24732
rect 23247 24701 23259 24704
rect 23201 24695 23259 24701
rect 23658 24624 23664 24676
rect 23716 24664 23722 24676
rect 24228 24664 24256 24763
rect 24302 24760 24308 24812
rect 24360 24760 24366 24812
rect 24946 24760 24952 24812
rect 25004 24800 25010 24812
rect 25133 24803 25191 24809
rect 25133 24800 25145 24803
rect 25004 24772 25145 24800
rect 25004 24760 25010 24772
rect 25133 24769 25145 24772
rect 25179 24800 25191 24803
rect 25240 24800 25268 24840
rect 25179 24772 25268 24800
rect 25317 24803 25375 24809
rect 25179 24769 25191 24772
rect 25133 24763 25191 24769
rect 25317 24769 25329 24803
rect 25363 24769 25375 24803
rect 25424 24800 25452 24840
rect 25774 24828 25780 24880
rect 25832 24828 25838 24880
rect 31772 24840 32812 24868
rect 31772 24812 31800 24840
rect 25685 24803 25743 24809
rect 25685 24800 25697 24803
rect 25424 24772 25697 24800
rect 25317 24763 25375 24769
rect 25685 24769 25697 24772
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 25332 24732 25360 24763
rect 25866 24760 25872 24812
rect 25924 24800 25930 24812
rect 26237 24803 26295 24809
rect 26237 24800 26249 24803
rect 25924 24772 26249 24800
rect 25924 24760 25930 24772
rect 26237 24769 26249 24772
rect 26283 24769 26295 24803
rect 26237 24763 26295 24769
rect 26421 24803 26479 24809
rect 26421 24769 26433 24803
rect 26467 24769 26479 24803
rect 26421 24763 26479 24769
rect 25501 24735 25559 24741
rect 25501 24732 25513 24735
rect 23716 24636 24256 24664
rect 24596 24704 25513 24732
rect 23716 24624 23722 24636
rect 23198 24596 23204 24608
rect 22520 24568 23204 24596
rect 22520 24556 22526 24568
rect 23198 24556 23204 24568
rect 23256 24556 23262 24608
rect 24213 24599 24271 24605
rect 24213 24565 24225 24599
rect 24259 24596 24271 24599
rect 24596 24596 24624 24704
rect 25501 24701 25513 24704
rect 25547 24701 25559 24735
rect 25501 24695 25559 24701
rect 25958 24692 25964 24744
rect 26016 24732 26022 24744
rect 26436 24732 26464 24763
rect 31754 24760 31760 24812
rect 31812 24760 31818 24812
rect 31938 24760 31944 24812
rect 31996 24800 32002 24812
rect 32784 24809 32812 24840
rect 34146 24828 34152 24880
rect 34204 24828 34210 24880
rect 32309 24803 32367 24809
rect 32309 24800 32321 24803
rect 31996 24772 32321 24800
rect 31996 24760 32002 24772
rect 32309 24769 32321 24772
rect 32355 24769 32367 24803
rect 32309 24763 32367 24769
rect 32769 24803 32827 24809
rect 32769 24769 32781 24803
rect 32815 24769 32827 24803
rect 32769 24763 32827 24769
rect 32950 24760 32956 24812
rect 33008 24809 33014 24812
rect 33008 24800 33019 24809
rect 33008 24772 33053 24800
rect 33008 24763 33019 24772
rect 33008 24760 33014 24763
rect 26016 24704 26464 24732
rect 32401 24735 32459 24741
rect 26016 24692 26022 24704
rect 32401 24701 32413 24735
rect 32447 24732 32459 24735
rect 32861 24735 32919 24741
rect 32861 24732 32873 24735
rect 32447 24704 32873 24732
rect 32447 24701 32459 24704
rect 32401 24695 32459 24701
rect 32861 24701 32873 24704
rect 32907 24701 32919 24735
rect 32861 24695 32919 24701
rect 33042 24692 33048 24744
rect 33100 24732 33106 24744
rect 33137 24735 33195 24741
rect 33137 24732 33149 24735
rect 33100 24704 33149 24732
rect 33100 24692 33106 24704
rect 33137 24701 33149 24704
rect 33183 24701 33195 24735
rect 33413 24735 33471 24741
rect 33413 24732 33425 24735
rect 33137 24695 33195 24701
rect 33244 24704 33425 24732
rect 25133 24667 25191 24673
rect 25133 24633 25145 24667
rect 25179 24664 25191 24667
rect 25590 24664 25596 24676
rect 25179 24636 25596 24664
rect 25179 24633 25191 24636
rect 25133 24627 25191 24633
rect 24259 24568 24624 24596
rect 24673 24599 24731 24605
rect 24259 24565 24271 24568
rect 24213 24559 24271 24565
rect 24673 24565 24685 24599
rect 24719 24596 24731 24599
rect 25148 24596 25176 24627
rect 25590 24624 25596 24636
rect 25648 24664 25654 24676
rect 25976 24664 26004 24692
rect 25648 24636 26004 24664
rect 32677 24667 32735 24673
rect 25648 24624 25654 24636
rect 32677 24633 32689 24667
rect 32723 24664 32735 24667
rect 33244 24664 33272 24704
rect 33413 24701 33425 24704
rect 33459 24701 33471 24735
rect 33413 24695 33471 24701
rect 32723 24636 33272 24664
rect 32723 24633 32735 24636
rect 32677 24627 32735 24633
rect 24719 24568 25176 24596
rect 26605 24599 26663 24605
rect 24719 24565 24731 24568
rect 24673 24559 24731 24565
rect 26605 24565 26617 24599
rect 26651 24596 26663 24599
rect 27154 24596 27160 24608
rect 26651 24568 27160 24596
rect 26651 24565 26663 24568
rect 26605 24559 26663 24565
rect 27154 24556 27160 24568
rect 27212 24556 27218 24608
rect 1104 24506 35248 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 35248 24506
rect 1104 24432 35248 24454
rect 9214 24352 9220 24404
rect 9272 24352 9278 24404
rect 10505 24395 10563 24401
rect 10505 24361 10517 24395
rect 10551 24392 10563 24395
rect 11146 24392 11152 24404
rect 10551 24364 11152 24392
rect 10551 24361 10563 24364
rect 10505 24355 10563 24361
rect 11146 24352 11152 24364
rect 11204 24352 11210 24404
rect 11425 24395 11483 24401
rect 11425 24361 11437 24395
rect 11471 24392 11483 24395
rect 12710 24392 12716 24404
rect 11471 24364 12716 24392
rect 11471 24361 11483 24364
rect 11425 24355 11483 24361
rect 12710 24352 12716 24364
rect 12768 24352 12774 24404
rect 14093 24395 14151 24401
rect 12820 24364 13124 24392
rect 9232 24265 9260 24352
rect 11882 24324 11888 24336
rect 10612 24296 11888 24324
rect 9217 24259 9275 24265
rect 9217 24225 9229 24259
rect 9263 24225 9275 24259
rect 9217 24219 9275 24225
rect 10410 24216 10416 24268
rect 10468 24216 10474 24268
rect 934 24148 940 24200
rect 992 24188 998 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 992 24160 1409 24188
rect 992 24148 998 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 3053 24191 3111 24197
rect 3053 24157 3065 24191
rect 3099 24188 3111 24191
rect 3973 24191 4031 24197
rect 3973 24188 3985 24191
rect 3099 24160 3985 24188
rect 3099 24157 3111 24160
rect 3053 24151 3111 24157
rect 3973 24157 3985 24160
rect 4019 24188 4031 24191
rect 4062 24188 4068 24200
rect 4019 24160 4068 24188
rect 4019 24157 4031 24160
rect 3973 24151 4031 24157
rect 4062 24148 4068 24160
rect 4120 24148 4126 24200
rect 9030 24148 9036 24200
rect 9088 24188 9094 24200
rect 10612 24197 10640 24296
rect 11882 24284 11888 24296
rect 11940 24324 11946 24336
rect 12066 24324 12072 24336
rect 11940 24296 12072 24324
rect 11940 24284 11946 24296
rect 12066 24284 12072 24296
rect 12124 24284 12130 24336
rect 12161 24327 12219 24333
rect 12161 24293 12173 24327
rect 12207 24324 12219 24327
rect 12820 24324 12848 24364
rect 13096 24336 13124 24364
rect 14093 24361 14105 24395
rect 14139 24392 14151 24395
rect 15194 24392 15200 24404
rect 14139 24364 15200 24392
rect 14139 24361 14151 24364
rect 14093 24355 14151 24361
rect 15194 24352 15200 24364
rect 15252 24352 15258 24404
rect 15286 24352 15292 24404
rect 15344 24352 15350 24404
rect 15838 24352 15844 24404
rect 15896 24392 15902 24404
rect 16577 24395 16635 24401
rect 16577 24392 16589 24395
rect 15896 24364 16589 24392
rect 15896 24352 15902 24364
rect 16577 24361 16589 24364
rect 16623 24361 16635 24395
rect 16577 24355 16635 24361
rect 17037 24395 17095 24401
rect 17037 24361 17049 24395
rect 17083 24392 17095 24395
rect 17126 24392 17132 24404
rect 17083 24364 17132 24392
rect 17083 24361 17095 24364
rect 17037 24355 17095 24361
rect 17126 24352 17132 24364
rect 17184 24352 17190 24404
rect 17221 24395 17279 24401
rect 17221 24361 17233 24395
rect 17267 24392 17279 24395
rect 17267 24364 17816 24392
rect 17267 24361 17279 24364
rect 17221 24355 17279 24361
rect 12207 24296 12848 24324
rect 12897 24327 12955 24333
rect 12207 24293 12219 24296
rect 12161 24287 12219 24293
rect 12897 24293 12909 24327
rect 12943 24293 12955 24327
rect 12897 24287 12955 24293
rect 10686 24216 10692 24268
rect 10744 24256 10750 24268
rect 11517 24259 11575 24265
rect 11517 24256 11529 24259
rect 10744 24228 10916 24256
rect 10744 24216 10750 24228
rect 10888 24197 10916 24228
rect 10980 24228 11529 24256
rect 10980 24197 11008 24228
rect 11517 24225 11529 24228
rect 11563 24225 11575 24259
rect 12802 24256 12808 24268
rect 11517 24219 11575 24225
rect 12084 24228 12808 24256
rect 10597 24191 10655 24197
rect 9088 24160 9154 24188
rect 9088 24148 9094 24160
rect 10597 24157 10609 24191
rect 10643 24157 10655 24191
rect 10597 24151 10655 24157
rect 10873 24191 10931 24197
rect 10873 24157 10885 24191
rect 10919 24157 10931 24191
rect 10873 24151 10931 24157
rect 10965 24191 11023 24197
rect 10965 24157 10977 24191
rect 11011 24157 11023 24191
rect 10965 24151 11023 24157
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 11149 24191 11207 24197
rect 11149 24188 11161 24191
rect 11112 24160 11161 24188
rect 11112 24148 11118 24160
rect 11149 24157 11161 24160
rect 11195 24157 11207 24191
rect 11149 24151 11207 24157
rect 11238 24148 11244 24200
rect 11296 24148 11302 24200
rect 11793 24191 11851 24197
rect 11793 24157 11805 24191
rect 11839 24157 11851 24191
rect 11793 24151 11851 24157
rect 10045 24123 10103 24129
rect 10045 24089 10057 24123
rect 10091 24089 10103 24123
rect 10045 24083 10103 24089
rect 10321 24123 10379 24129
rect 10321 24089 10333 24123
rect 10367 24120 10379 24123
rect 10686 24120 10692 24132
rect 10367 24092 10692 24120
rect 10367 24089 10379 24092
rect 10321 24083 10379 24089
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24052 1639 24055
rect 2038 24052 2044 24064
rect 1627 24024 2044 24052
rect 1627 24021 1639 24024
rect 1581 24015 1639 24021
rect 2038 24012 2044 24024
rect 2096 24012 2102 24064
rect 2958 24012 2964 24064
rect 3016 24012 3022 24064
rect 3418 24012 3424 24064
rect 3476 24012 3482 24064
rect 6638 24012 6644 24064
rect 6696 24052 6702 24064
rect 8297 24055 8355 24061
rect 8297 24052 8309 24055
rect 6696 24024 8309 24052
rect 6696 24012 6702 24024
rect 8297 24021 8309 24024
rect 8343 24052 8355 24055
rect 8573 24055 8631 24061
rect 8573 24052 8585 24055
rect 8343 24024 8585 24052
rect 8343 24021 8355 24024
rect 8297 24015 8355 24021
rect 8573 24021 8585 24024
rect 8619 24021 8631 24055
rect 10060 24052 10088 24083
rect 10686 24080 10692 24092
rect 10744 24080 10750 24132
rect 10781 24123 10839 24129
rect 10781 24089 10793 24123
rect 10827 24120 10839 24123
rect 11808 24120 11836 24151
rect 11882 24148 11888 24200
rect 11940 24148 11946 24200
rect 12084 24154 12112 24228
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 12912 24256 12940 24287
rect 13078 24284 13084 24336
rect 13136 24284 13142 24336
rect 14553 24327 14611 24333
rect 14553 24293 14565 24327
rect 14599 24324 14611 24327
rect 15746 24324 15752 24336
rect 14599 24296 15752 24324
rect 14599 24293 14611 24296
rect 14553 24287 14611 24293
rect 15746 24284 15752 24296
rect 15804 24284 15810 24336
rect 16298 24284 16304 24336
rect 16356 24284 16362 24336
rect 17144 24324 17172 24352
rect 17144 24296 17264 24324
rect 13998 24256 14004 24268
rect 12912 24228 14004 24256
rect 13998 24216 14004 24228
rect 14056 24256 14062 24268
rect 14056 24228 14412 24256
rect 14056 24216 14062 24228
rect 11992 24126 12112 24154
rect 12253 24191 12311 24197
rect 12253 24157 12265 24191
rect 12299 24188 12311 24191
rect 12526 24188 12532 24200
rect 12299 24160 12532 24188
rect 12299 24157 12311 24160
rect 12253 24151 12311 24157
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 12621 24191 12679 24197
rect 12621 24157 12633 24191
rect 12667 24188 12679 24191
rect 12820 24188 12848 24216
rect 12667 24160 12848 24188
rect 12897 24191 12955 24197
rect 12667 24157 12679 24160
rect 12621 24151 12679 24157
rect 12897 24157 12909 24191
rect 12943 24188 12955 24191
rect 12989 24191 13047 24197
rect 12989 24188 13001 24191
rect 12943 24160 13001 24188
rect 12943 24157 12955 24160
rect 12897 24151 12955 24157
rect 12989 24157 13001 24160
rect 13035 24188 13047 24191
rect 13078 24188 13084 24200
rect 13035 24160 13084 24188
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13170 24148 13176 24200
rect 13228 24188 13234 24200
rect 14384 24197 14412 24228
rect 15286 24216 15292 24268
rect 15344 24256 15350 24268
rect 15657 24259 15715 24265
rect 15657 24256 15669 24259
rect 15344 24228 15669 24256
rect 15344 24216 15350 24228
rect 15657 24225 15669 24228
rect 15703 24256 15715 24259
rect 16316 24256 16344 24284
rect 15703 24228 16344 24256
rect 15703 24225 15715 24228
rect 15657 24219 15715 24225
rect 16390 24216 16396 24268
rect 16448 24256 16454 24268
rect 16448 24228 17172 24256
rect 16448 24216 16454 24228
rect 13474 24191 13532 24197
rect 13474 24188 13486 24191
rect 13228 24160 13486 24188
rect 13228 24148 13234 24160
rect 13474 24157 13486 24160
rect 13520 24157 13532 24191
rect 13474 24151 13532 24157
rect 14369 24191 14427 24197
rect 14369 24157 14381 24191
rect 14415 24188 14427 24191
rect 14461 24191 14519 24197
rect 14461 24188 14473 24191
rect 14415 24160 14473 24188
rect 14415 24157 14427 24160
rect 14369 24151 14427 24157
rect 14461 24157 14473 24160
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14550 24148 14556 24200
rect 14608 24188 14614 24200
rect 14645 24191 14703 24197
rect 14645 24188 14657 24191
rect 14608 24160 14657 24188
rect 14608 24148 14614 24160
rect 14645 24157 14657 24160
rect 14691 24157 14703 24191
rect 14645 24151 14703 24157
rect 15470 24148 15476 24200
rect 15528 24148 15534 24200
rect 15746 24148 15752 24200
rect 15804 24188 15810 24200
rect 17144 24197 17172 24228
rect 16485 24191 16543 24197
rect 16485 24188 16497 24191
rect 15804 24160 16497 24188
rect 15804 24148 15810 24160
rect 16485 24157 16497 24160
rect 16531 24157 16543 24191
rect 16485 24151 16543 24157
rect 17129 24191 17187 24197
rect 17129 24157 17141 24191
rect 17175 24157 17187 24191
rect 17236 24188 17264 24296
rect 17313 24191 17371 24197
rect 17313 24188 17325 24191
rect 17236 24160 17325 24188
rect 17129 24151 17187 24157
rect 17313 24157 17325 24160
rect 17359 24188 17371 24191
rect 17359 24160 17540 24188
rect 17788 24174 17816 24364
rect 22186 24352 22192 24404
rect 22244 24392 22250 24404
rect 22370 24392 22376 24404
rect 22244 24364 22376 24392
rect 22244 24352 22250 24364
rect 22370 24352 22376 24364
rect 22428 24392 22434 24404
rect 22557 24395 22615 24401
rect 22557 24392 22569 24395
rect 22428 24364 22569 24392
rect 22428 24352 22434 24364
rect 22557 24361 22569 24364
rect 22603 24392 22615 24395
rect 22830 24392 22836 24404
rect 22603 24364 22836 24392
rect 22603 24361 22615 24364
rect 22557 24355 22615 24361
rect 22830 24352 22836 24364
rect 22888 24352 22894 24404
rect 25866 24352 25872 24404
rect 25924 24352 25930 24404
rect 28074 24352 28080 24404
rect 28132 24392 28138 24404
rect 28169 24395 28227 24401
rect 28169 24392 28181 24395
rect 28132 24364 28181 24392
rect 28132 24352 28138 24364
rect 28169 24361 28181 24364
rect 28215 24361 28227 24395
rect 31573 24395 31631 24401
rect 28169 24355 28227 24361
rect 28276 24364 29408 24392
rect 20254 24324 20260 24336
rect 19306 24296 20260 24324
rect 18230 24216 18236 24268
rect 18288 24216 18294 24268
rect 17359 24157 17371 24160
rect 17313 24151 17371 24157
rect 11992 24120 12020 24126
rect 10827 24092 12020 24120
rect 10827 24089 10839 24092
rect 10781 24083 10839 24089
rect 12158 24080 12164 24132
rect 12216 24080 12222 24132
rect 12342 24080 12348 24132
rect 12400 24120 12406 24132
rect 13265 24123 13323 24129
rect 13265 24120 13277 24123
rect 12400 24092 13277 24120
rect 12400 24080 12406 24092
rect 13265 24089 13277 24092
rect 13311 24089 13323 24123
rect 13265 24083 13323 24089
rect 14093 24123 14151 24129
rect 14093 24089 14105 24123
rect 14139 24089 14151 24123
rect 16500 24120 16528 24151
rect 17405 24123 17463 24129
rect 17405 24120 17417 24123
rect 16500 24092 17417 24120
rect 14093 24083 14151 24089
rect 17405 24089 17417 24092
rect 17451 24089 17463 24123
rect 17512 24120 17540 24160
rect 19306 24120 19334 24296
rect 20254 24284 20260 24296
rect 20312 24324 20318 24336
rect 20625 24327 20683 24333
rect 20625 24324 20637 24327
rect 20312 24296 20637 24324
rect 20312 24284 20318 24296
rect 20625 24293 20637 24296
rect 20671 24324 20683 24327
rect 20993 24327 21051 24333
rect 20993 24324 21005 24327
rect 20671 24296 21005 24324
rect 20671 24293 20683 24296
rect 20625 24287 20683 24293
rect 20993 24293 21005 24296
rect 21039 24324 21051 24327
rect 21082 24324 21088 24336
rect 21039 24296 21088 24324
rect 21039 24293 21051 24296
rect 20993 24287 21051 24293
rect 21082 24284 21088 24296
rect 21140 24284 21146 24336
rect 21008 24228 25728 24256
rect 21008 24200 21036 24228
rect 20990 24148 20996 24200
rect 21048 24148 21054 24200
rect 21726 24148 21732 24200
rect 21784 24188 21790 24200
rect 22186 24188 22192 24200
rect 21784 24160 22192 24188
rect 21784 24148 21790 24160
rect 22186 24148 22192 24160
rect 22244 24148 22250 24200
rect 25590 24148 25596 24200
rect 25648 24148 25654 24200
rect 17512 24092 19334 24120
rect 17405 24083 17463 24089
rect 11974 24052 11980 24064
rect 10060 24024 11980 24052
rect 8573 24015 8631 24021
rect 11974 24012 11980 24024
rect 12032 24012 12038 24064
rect 12176 24052 12204 24080
rect 12713 24055 12771 24061
rect 12713 24052 12725 24055
rect 12176 24024 12725 24052
rect 12713 24021 12725 24024
rect 12759 24021 12771 24055
rect 12713 24015 12771 24021
rect 12802 24012 12808 24064
rect 12860 24052 12866 24064
rect 13357 24055 13415 24061
rect 13357 24052 13369 24055
rect 12860 24024 13369 24052
rect 12860 24012 12866 24024
rect 13357 24021 13369 24024
rect 13403 24021 13415 24055
rect 13357 24015 13415 24021
rect 13633 24055 13691 24061
rect 13633 24021 13645 24055
rect 13679 24052 13691 24055
rect 14108 24052 14136 24083
rect 21358 24080 21364 24132
rect 21416 24120 21422 24132
rect 25700 24120 25728 24228
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24188 25835 24191
rect 25884 24188 25912 24352
rect 27062 24284 27068 24336
rect 27120 24284 27126 24336
rect 27985 24327 28043 24333
rect 27985 24293 27997 24327
rect 28031 24324 28043 24327
rect 28276 24324 28304 24364
rect 28718 24324 28724 24336
rect 28031 24296 28304 24324
rect 28031 24293 28043 24296
rect 27985 24287 28043 24293
rect 27157 24259 27215 24265
rect 27157 24225 27169 24259
rect 27203 24256 27215 24259
rect 27338 24256 27344 24268
rect 27203 24228 27344 24256
rect 27203 24225 27215 24228
rect 27157 24219 27215 24225
rect 27338 24216 27344 24228
rect 27396 24216 27402 24268
rect 27614 24216 27620 24268
rect 27672 24256 27678 24268
rect 27672 24228 28212 24256
rect 27672 24216 27678 24228
rect 25823 24160 25912 24188
rect 26053 24191 26111 24197
rect 25823 24157 25835 24160
rect 25777 24151 25835 24157
rect 26053 24157 26065 24191
rect 26099 24157 26111 24191
rect 26053 24151 26111 24157
rect 26237 24191 26295 24197
rect 26237 24157 26249 24191
rect 26283 24188 26295 24191
rect 26329 24191 26387 24197
rect 26329 24188 26341 24191
rect 26283 24160 26341 24188
rect 26283 24157 26295 24160
rect 26237 24151 26295 24157
rect 26329 24157 26341 24160
rect 26375 24157 26387 24191
rect 26329 24151 26387 24157
rect 26697 24191 26755 24197
rect 26697 24157 26709 24191
rect 26743 24157 26755 24191
rect 26697 24151 26755 24157
rect 26068 24120 26096 24151
rect 21416 24092 22968 24120
rect 25700 24092 26096 24120
rect 26712 24120 26740 24151
rect 26970 24148 26976 24200
rect 27028 24148 27034 24200
rect 27430 24148 27436 24200
rect 27488 24148 27494 24200
rect 27632 24188 27660 24216
rect 27709 24191 27767 24197
rect 27709 24188 27721 24191
rect 27632 24160 27721 24188
rect 27709 24157 27721 24160
rect 27755 24157 27767 24191
rect 27709 24151 27767 24157
rect 27893 24191 27951 24197
rect 27893 24157 27905 24191
rect 27939 24157 27951 24191
rect 28077 24191 28135 24197
rect 28077 24188 28089 24191
rect 27893 24151 27951 24157
rect 28000 24160 28089 24188
rect 27249 24123 27307 24129
rect 27249 24120 27261 24123
rect 26712 24092 27261 24120
rect 21416 24080 21422 24092
rect 22940 24064 22968 24092
rect 13679 24024 14136 24052
rect 13679 24021 13691 24024
rect 13633 24015 13691 24021
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 14366 24012 14372 24064
rect 14424 24052 14430 24064
rect 20070 24052 20076 24064
rect 14424 24024 20076 24052
rect 14424 24012 14430 24024
rect 20070 24012 20076 24024
rect 20128 24052 20134 24064
rect 20165 24055 20223 24061
rect 20165 24052 20177 24055
rect 20128 24024 20177 24052
rect 20128 24012 20134 24024
rect 20165 24021 20177 24024
rect 20211 24052 20223 24055
rect 20438 24052 20444 24064
rect 20211 24024 20444 24052
rect 20211 24021 20223 24024
rect 20165 24015 20223 24021
rect 20438 24012 20444 24024
rect 20496 24012 20502 24064
rect 21729 24055 21787 24061
rect 21729 24021 21741 24055
rect 21775 24052 21787 24055
rect 22186 24052 22192 24064
rect 21775 24024 22192 24052
rect 21775 24021 21787 24024
rect 21729 24015 21787 24021
rect 22186 24012 22192 24024
rect 22244 24012 22250 24064
rect 22922 24012 22928 24064
rect 22980 24052 22986 24064
rect 23017 24055 23075 24061
rect 23017 24052 23029 24055
rect 22980 24024 23029 24052
rect 22980 24012 22986 24024
rect 23017 24021 23029 24024
rect 23063 24021 23075 24055
rect 23017 24015 23075 24021
rect 23382 24012 23388 24064
rect 23440 24012 23446 24064
rect 26068 24052 26096 24092
rect 27249 24089 27261 24092
rect 27295 24089 27307 24123
rect 27798 24120 27804 24132
rect 27249 24083 27307 24089
rect 27448 24092 27804 24120
rect 27448 24052 27476 24092
rect 27798 24080 27804 24092
rect 27856 24120 27862 24132
rect 27908 24120 27936 24151
rect 28000 24132 28028 24160
rect 28077 24157 28089 24160
rect 28123 24157 28135 24191
rect 28077 24151 28135 24157
rect 27856 24092 27936 24120
rect 27856 24080 27862 24092
rect 27982 24080 27988 24132
rect 28040 24080 28046 24132
rect 28184 24120 28212 24228
rect 28276 24188 28304 24296
rect 28460 24296 28724 24324
rect 28460 24197 28488 24296
rect 28718 24284 28724 24296
rect 28776 24284 28782 24336
rect 28537 24259 28595 24265
rect 28537 24225 28549 24259
rect 28583 24225 28595 24259
rect 28537 24219 28595 24225
rect 28353 24191 28411 24197
rect 28353 24188 28365 24191
rect 28276 24160 28365 24188
rect 28353 24157 28365 24160
rect 28399 24157 28411 24191
rect 28353 24151 28411 24157
rect 28445 24191 28503 24197
rect 28445 24157 28457 24191
rect 28491 24157 28503 24191
rect 28445 24151 28503 24157
rect 28460 24120 28488 24151
rect 28184 24092 28488 24120
rect 26068 24024 27476 24052
rect 27522 24012 27528 24064
rect 27580 24052 27586 24064
rect 27617 24055 27675 24061
rect 27617 24052 27629 24055
rect 27580 24024 27629 24052
rect 27580 24012 27586 24024
rect 27617 24021 27629 24024
rect 27663 24052 27675 24055
rect 28552 24052 28580 24219
rect 29086 24216 29092 24268
rect 29144 24216 29150 24268
rect 29380 24200 29408 24364
rect 31573 24361 31585 24395
rect 31619 24392 31631 24395
rect 31938 24392 31944 24404
rect 31619 24364 31944 24392
rect 31619 24361 31631 24364
rect 31573 24355 31631 24361
rect 31938 24352 31944 24364
rect 31996 24352 32002 24404
rect 34146 24352 34152 24404
rect 34204 24392 34210 24404
rect 34241 24395 34299 24401
rect 34241 24392 34253 24395
rect 34204 24364 34253 24392
rect 34204 24352 34210 24364
rect 34241 24361 34253 24364
rect 34287 24361 34299 24395
rect 34241 24355 34299 24361
rect 29638 24216 29644 24268
rect 29696 24256 29702 24268
rect 29825 24259 29883 24265
rect 29825 24256 29837 24259
rect 29696 24228 29837 24256
rect 29696 24216 29702 24228
rect 29825 24225 29837 24228
rect 29871 24225 29883 24259
rect 29825 24219 29883 24225
rect 28626 24148 28632 24200
rect 28684 24148 28690 24200
rect 28994 24148 29000 24200
rect 29052 24148 29058 24200
rect 29362 24148 29368 24200
rect 29420 24148 29426 24200
rect 34149 24191 34207 24197
rect 34149 24188 34161 24191
rect 34072 24160 34161 24188
rect 30101 24123 30159 24129
rect 30101 24120 30113 24123
rect 29380 24092 30113 24120
rect 28902 24052 28908 24064
rect 27663 24024 28908 24052
rect 27663 24021 27675 24024
rect 27617 24015 27675 24021
rect 28902 24012 28908 24024
rect 28960 24012 28966 24064
rect 29380 24061 29408 24092
rect 30101 24089 30113 24092
rect 30147 24089 30159 24123
rect 30101 24083 30159 24089
rect 30834 24080 30840 24132
rect 30892 24080 30898 24132
rect 34072 24064 34100 24160
rect 34149 24157 34161 24160
rect 34195 24188 34207 24191
rect 34514 24188 34520 24200
rect 34195 24160 34520 24188
rect 34195 24157 34207 24160
rect 34149 24151 34207 24157
rect 34514 24148 34520 24160
rect 34572 24148 34578 24200
rect 29365 24055 29423 24061
rect 29365 24021 29377 24055
rect 29411 24021 29423 24055
rect 29365 24015 29423 24021
rect 32674 24012 32680 24064
rect 32732 24052 32738 24064
rect 32953 24055 33011 24061
rect 32953 24052 32965 24055
rect 32732 24024 32965 24052
rect 32732 24012 32738 24024
rect 32953 24021 32965 24024
rect 32999 24052 33011 24055
rect 33042 24052 33048 24064
rect 32999 24024 33048 24052
rect 32999 24021 33011 24024
rect 32953 24015 33011 24021
rect 33042 24012 33048 24024
rect 33100 24012 33106 24064
rect 34054 24012 34060 24064
rect 34112 24012 34118 24064
rect 1104 23962 35236 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 35236 23962
rect 1104 23888 35236 23910
rect 11698 23808 11704 23860
rect 11756 23808 11762 23860
rect 11974 23808 11980 23860
rect 12032 23848 12038 23860
rect 12342 23848 12348 23860
rect 12032 23820 12348 23848
rect 12032 23808 12038 23820
rect 12342 23808 12348 23820
rect 12400 23808 12406 23860
rect 13170 23808 13176 23860
rect 13228 23808 13234 23860
rect 15289 23851 15347 23857
rect 15289 23817 15301 23851
rect 15335 23848 15347 23851
rect 15470 23848 15476 23860
rect 15335 23820 15476 23848
rect 15335 23817 15347 23820
rect 15289 23811 15347 23817
rect 15470 23808 15476 23820
rect 15528 23808 15534 23860
rect 15746 23808 15752 23860
rect 15804 23808 15810 23860
rect 15838 23808 15844 23860
rect 15896 23808 15902 23860
rect 17865 23851 17923 23857
rect 17865 23817 17877 23851
rect 17911 23848 17923 23851
rect 18230 23848 18236 23860
rect 17911 23820 18236 23848
rect 17911 23817 17923 23820
rect 17865 23811 17923 23817
rect 18230 23808 18236 23820
rect 18288 23808 18294 23860
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 21545 23851 21603 23857
rect 21545 23848 21557 23851
rect 20588 23820 21557 23848
rect 20588 23808 20594 23820
rect 21545 23817 21557 23820
rect 21591 23848 21603 23851
rect 21726 23848 21732 23860
rect 21591 23820 21732 23848
rect 21591 23817 21603 23820
rect 21545 23811 21603 23817
rect 21726 23808 21732 23820
rect 21784 23808 21790 23860
rect 22189 23851 22247 23857
rect 22189 23817 22201 23851
rect 22235 23817 22247 23851
rect 22189 23811 22247 23817
rect 22557 23851 22615 23857
rect 22557 23817 22569 23851
rect 22603 23848 22615 23851
rect 23658 23848 23664 23860
rect 22603 23820 23664 23848
rect 22603 23817 22615 23820
rect 22557 23811 22615 23817
rect 1854 23740 1860 23792
rect 1912 23740 1918 23792
rect 3694 23740 3700 23792
rect 3752 23740 3758 23792
rect 4706 23740 4712 23792
rect 4764 23740 4770 23792
rect 6638 23780 6644 23792
rect 6472 23752 6644 23780
rect 2958 23672 2964 23724
rect 3016 23672 3022 23724
rect 3418 23672 3424 23724
rect 3476 23672 3482 23724
rect 6472 23721 6500 23752
rect 6638 23740 6644 23752
rect 6696 23740 6702 23792
rect 8294 23780 8300 23792
rect 7958 23752 8300 23780
rect 8294 23740 8300 23752
rect 8352 23740 8358 23792
rect 9401 23783 9459 23789
rect 9401 23749 9413 23783
rect 9447 23780 9459 23783
rect 9447 23752 9996 23780
rect 9447 23749 9459 23752
rect 9401 23743 9459 23749
rect 9968 23721 9996 23752
rect 10962 23740 10968 23792
rect 11020 23780 11026 23792
rect 12621 23783 12679 23789
rect 12621 23780 12633 23783
rect 11020 23752 12633 23780
rect 11020 23740 11026 23752
rect 12621 23749 12633 23752
rect 12667 23749 12679 23783
rect 12621 23743 12679 23749
rect 5445 23715 5503 23721
rect 5445 23712 5457 23715
rect 5184 23684 5457 23712
rect 1394 23604 1400 23656
rect 1452 23644 1458 23656
rect 1581 23647 1639 23653
rect 1581 23644 1593 23647
rect 1452 23616 1593 23644
rect 1452 23604 1458 23616
rect 1581 23613 1593 23616
rect 1627 23613 1639 23647
rect 1581 23607 1639 23613
rect 5184 23520 5212 23684
rect 5445 23681 5457 23684
rect 5491 23681 5503 23715
rect 5445 23675 5503 23681
rect 6181 23715 6239 23721
rect 6181 23681 6193 23715
rect 6227 23712 6239 23715
rect 6457 23715 6515 23721
rect 6457 23712 6469 23715
rect 6227 23684 6469 23712
rect 6227 23681 6239 23684
rect 6181 23675 6239 23681
rect 6457 23681 6469 23684
rect 6503 23681 6515 23715
rect 8573 23715 8631 23721
rect 8573 23712 8585 23715
rect 6457 23675 6515 23681
rect 8220 23684 8585 23712
rect 5350 23604 5356 23656
rect 5408 23604 5414 23656
rect 8220 23653 8248 23684
rect 8573 23681 8585 23684
rect 8619 23681 8631 23715
rect 8573 23675 8631 23681
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23681 9827 23715
rect 9769 23675 9827 23681
rect 9953 23715 10011 23721
rect 9953 23681 9965 23715
rect 9999 23712 10011 23715
rect 10594 23712 10600 23724
rect 9999 23684 10600 23712
rect 9999 23681 10011 23684
rect 9953 23675 10011 23681
rect 6733 23647 6791 23653
rect 6733 23644 6745 23647
rect 6564 23616 6745 23644
rect 5813 23579 5871 23585
rect 5813 23545 5825 23579
rect 5859 23576 5871 23579
rect 6564 23576 6592 23616
rect 6733 23613 6745 23616
rect 6779 23613 6791 23647
rect 6733 23607 6791 23613
rect 8205 23647 8263 23653
rect 8205 23613 8217 23647
rect 8251 23613 8263 23647
rect 9784 23644 9812 23675
rect 10594 23672 10600 23684
rect 10652 23672 10658 23724
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 11164 23684 11529 23712
rect 11164 23644 11192 23684
rect 11517 23681 11529 23684
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 11701 23715 11759 23721
rect 11701 23681 11713 23715
rect 11747 23712 11759 23715
rect 11747 23684 12112 23712
rect 11747 23681 11759 23684
rect 11701 23675 11759 23681
rect 9784 23616 11192 23644
rect 8205 23607 8263 23613
rect 5859 23548 6592 23576
rect 5859 23545 5871 23548
rect 5813 23539 5871 23545
rect 3329 23511 3387 23517
rect 3329 23477 3341 23511
rect 3375 23508 3387 23511
rect 4798 23508 4804 23520
rect 3375 23480 4804 23508
rect 3375 23477 3387 23480
rect 3329 23471 3387 23477
rect 4798 23468 4804 23480
rect 4856 23468 4862 23520
rect 5166 23468 5172 23520
rect 5224 23468 5230 23520
rect 9769 23511 9827 23517
rect 9769 23477 9781 23511
rect 9815 23508 9827 23511
rect 10226 23508 10232 23520
rect 9815 23480 10232 23508
rect 9815 23477 9827 23480
rect 9769 23471 9827 23477
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 10413 23511 10471 23517
rect 10413 23477 10425 23511
rect 10459 23508 10471 23511
rect 10594 23508 10600 23520
rect 10459 23480 10600 23508
rect 10459 23477 10471 23480
rect 10413 23471 10471 23477
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 10778 23468 10784 23520
rect 10836 23508 10842 23520
rect 11164 23517 11192 23616
rect 12084 23517 12112 23684
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 12802 23712 12808 23724
rect 12584 23684 12808 23712
rect 12584 23672 12590 23684
rect 12802 23672 12808 23684
rect 12860 23672 12866 23724
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23712 12955 23715
rect 13188 23712 13216 23808
rect 14550 23780 14556 23792
rect 13740 23752 14556 23780
rect 13740 23721 13768 23752
rect 14550 23740 14556 23752
rect 14608 23740 14614 23792
rect 15764 23780 15792 23808
rect 15304 23752 15516 23780
rect 15304 23724 15332 23752
rect 13725 23715 13783 23721
rect 13725 23712 13737 23715
rect 12943 23684 13216 23712
rect 13556 23684 13737 23712
rect 12943 23681 12955 23684
rect 12897 23675 12955 23681
rect 13556 23644 13584 23684
rect 13725 23681 13737 23684
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 13817 23715 13875 23721
rect 13817 23681 13829 23715
rect 13863 23712 13875 23715
rect 14274 23712 14280 23724
rect 13863 23684 14280 23712
rect 13863 23681 13875 23684
rect 13817 23675 13875 23681
rect 13832 23644 13860 23675
rect 14274 23672 14280 23684
rect 14332 23672 14338 23724
rect 15286 23672 15292 23724
rect 15344 23672 15350 23724
rect 15378 23672 15384 23724
rect 15436 23672 15442 23724
rect 15488 23721 15516 23752
rect 15580 23752 15792 23780
rect 15856 23780 15884 23808
rect 17497 23783 17555 23789
rect 15856 23752 16896 23780
rect 15580 23721 15608 23752
rect 15473 23715 15531 23721
rect 15473 23681 15485 23715
rect 15519 23681 15531 23715
rect 15473 23675 15531 23681
rect 15565 23715 15623 23721
rect 15565 23681 15577 23715
rect 15611 23681 15623 23715
rect 15565 23675 15623 23681
rect 15746 23672 15752 23724
rect 15804 23672 15810 23724
rect 15841 23715 15899 23721
rect 15841 23681 15853 23715
rect 15887 23681 15899 23715
rect 16482 23712 16488 23724
rect 15841 23675 15899 23681
rect 15948 23684 16488 23712
rect 12176 23616 13584 23644
rect 13740 23616 13860 23644
rect 12176 23588 12204 23616
rect 12158 23536 12164 23588
rect 12216 23536 12222 23588
rect 12897 23579 12955 23585
rect 12897 23545 12909 23579
rect 12943 23576 12955 23579
rect 13740 23576 13768 23616
rect 13998 23604 14004 23656
rect 14056 23604 14062 23656
rect 15396 23644 15424 23672
rect 15856 23644 15884 23675
rect 15396 23616 15884 23644
rect 15948 23576 15976 23684
rect 16482 23672 16488 23684
rect 16540 23672 16546 23724
rect 16868 23721 16896 23752
rect 17497 23749 17509 23783
rect 17543 23780 17555 23783
rect 17954 23780 17960 23792
rect 17543 23752 17960 23780
rect 17543 23749 17555 23752
rect 17497 23743 17555 23749
rect 17954 23740 17960 23752
rect 18012 23740 18018 23792
rect 20349 23783 20407 23789
rect 20349 23749 20361 23783
rect 20395 23780 20407 23783
rect 20717 23783 20775 23789
rect 20717 23780 20729 23783
rect 20395 23752 20729 23780
rect 20395 23749 20407 23752
rect 20349 23743 20407 23749
rect 20717 23749 20729 23752
rect 20763 23749 20775 23783
rect 20717 23743 20775 23749
rect 20809 23783 20867 23789
rect 20809 23749 20821 23783
rect 20855 23780 20867 23783
rect 21082 23780 21088 23792
rect 20855 23752 21088 23780
rect 20855 23749 20867 23752
rect 20809 23743 20867 23749
rect 21082 23740 21088 23752
rect 21140 23740 21146 23792
rect 22204 23780 22232 23811
rect 23658 23808 23664 23820
rect 23716 23808 23722 23860
rect 24765 23851 24823 23857
rect 24765 23817 24777 23851
rect 24811 23848 24823 23851
rect 24811 23820 25176 23848
rect 24811 23817 24823 23820
rect 24765 23811 24823 23817
rect 23382 23780 23388 23792
rect 22204 23752 22600 23780
rect 16853 23715 16911 23721
rect 16853 23681 16865 23715
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17586 23672 17592 23724
rect 17644 23712 17650 23724
rect 17681 23715 17739 23721
rect 17681 23712 17693 23715
rect 17644 23684 17693 23712
rect 17644 23672 17650 23684
rect 17681 23681 17693 23684
rect 17727 23681 17739 23715
rect 17681 23675 17739 23681
rect 17865 23715 17923 23721
rect 17865 23681 17877 23715
rect 17911 23712 17923 23715
rect 17972 23712 18000 23740
rect 17911 23684 18000 23712
rect 17911 23681 17923 23684
rect 17865 23675 17923 23681
rect 16298 23604 16304 23656
rect 16356 23644 16362 23656
rect 16761 23647 16819 23653
rect 16761 23644 16773 23647
rect 16356 23616 16773 23644
rect 16356 23604 16362 23616
rect 16761 23613 16773 23616
rect 16807 23613 16819 23647
rect 17696 23644 17724 23675
rect 20254 23672 20260 23724
rect 20312 23672 20318 23724
rect 20441 23715 20499 23721
rect 20441 23681 20453 23715
rect 20487 23681 20499 23715
rect 20441 23675 20499 23681
rect 18141 23647 18199 23653
rect 18141 23644 18153 23647
rect 17696 23616 18153 23644
rect 16761 23607 16819 23613
rect 18141 23613 18153 23616
rect 18187 23613 18199 23647
rect 20456 23644 20484 23675
rect 20530 23672 20536 23724
rect 20588 23672 20594 23724
rect 20901 23715 20959 23721
rect 20901 23681 20913 23715
rect 20947 23712 20959 23715
rect 22094 23712 22100 23724
rect 20947 23684 22100 23712
rect 20947 23681 20959 23684
rect 20901 23675 20959 23681
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 22186 23672 22192 23724
rect 22244 23672 22250 23724
rect 22462 23672 22468 23724
rect 22520 23672 22526 23724
rect 18141 23607 18199 23613
rect 19904 23616 20484 23644
rect 12943 23548 13768 23576
rect 13832 23548 15976 23576
rect 12943 23545 12955 23548
rect 12897 23539 12955 23545
rect 11149 23511 11207 23517
rect 11149 23508 11161 23511
rect 10836 23480 11161 23508
rect 10836 23468 10842 23480
rect 11149 23477 11161 23480
rect 11195 23477 11207 23511
rect 11149 23471 11207 23477
rect 12069 23511 12127 23517
rect 12069 23477 12081 23511
rect 12115 23508 12127 23511
rect 12434 23508 12440 23520
rect 12115 23480 12440 23508
rect 12115 23477 12127 23480
rect 12069 23471 12127 23477
rect 12434 23468 12440 23480
rect 12492 23508 12498 23520
rect 13832 23508 13860 23548
rect 12492 23480 13860 23508
rect 13909 23511 13967 23517
rect 12492 23468 12498 23480
rect 13909 23477 13921 23511
rect 13955 23508 13967 23511
rect 15194 23508 15200 23520
rect 13955 23480 15200 23508
rect 13955 23477 13967 23480
rect 13909 23471 13967 23477
rect 15194 23468 15200 23480
rect 15252 23468 15258 23520
rect 17126 23468 17132 23520
rect 17184 23468 17190 23520
rect 19242 23468 19248 23520
rect 19300 23508 19306 23520
rect 19904 23517 19932 23616
rect 19889 23511 19947 23517
rect 19889 23508 19901 23511
rect 19300 23480 19901 23508
rect 19300 23468 19306 23480
rect 19889 23477 19901 23480
rect 19935 23477 19947 23511
rect 20456 23508 20484 23616
rect 21100 23616 21772 23644
rect 21100 23585 21128 23616
rect 21085 23579 21143 23585
rect 21085 23545 21097 23579
rect 21131 23545 21143 23579
rect 21744 23576 21772 23616
rect 21818 23604 21824 23656
rect 21876 23604 21882 23656
rect 22373 23647 22431 23653
rect 22373 23644 22385 23647
rect 22066 23616 22385 23644
rect 22066 23576 22094 23616
rect 22373 23613 22385 23616
rect 22419 23613 22431 23647
rect 22572 23644 22600 23752
rect 22756 23752 23388 23780
rect 22756 23724 22784 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 24949 23783 25007 23789
rect 24949 23749 24961 23783
rect 24995 23780 25007 23783
rect 25038 23780 25044 23792
rect 24995 23752 25044 23780
rect 24995 23749 25007 23752
rect 24949 23743 25007 23749
rect 22646 23672 22652 23724
rect 22704 23672 22710 23724
rect 22738 23672 22744 23724
rect 22796 23672 22802 23724
rect 22830 23672 22836 23724
rect 22888 23712 22894 23724
rect 22925 23715 22983 23721
rect 22925 23712 22937 23715
rect 22888 23684 22937 23712
rect 22888 23672 22894 23684
rect 22925 23681 22937 23684
rect 22971 23712 22983 23715
rect 23201 23715 23259 23721
rect 23201 23712 23213 23715
rect 22971 23684 23213 23712
rect 22971 23681 22983 23684
rect 22925 23675 22983 23681
rect 23201 23681 23213 23684
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 24486 23672 24492 23724
rect 24544 23712 24550 23724
rect 24581 23715 24639 23721
rect 24581 23712 24593 23715
rect 24544 23684 24593 23712
rect 24544 23672 24550 23684
rect 24581 23681 24593 23684
rect 24627 23681 24639 23715
rect 24581 23675 24639 23681
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23712 24915 23715
rect 24964 23712 24992 23743
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 25148 23789 25176 23820
rect 26970 23808 26976 23860
rect 27028 23808 27034 23860
rect 27154 23857 27160 23860
rect 27141 23851 27160 23857
rect 27141 23817 27153 23851
rect 27141 23811 27160 23817
rect 27154 23808 27160 23811
rect 27212 23808 27218 23860
rect 28626 23808 28632 23860
rect 28684 23808 28690 23860
rect 28718 23808 28724 23860
rect 28776 23808 28782 23860
rect 28902 23808 28908 23860
rect 28960 23808 28966 23860
rect 28994 23808 29000 23860
rect 29052 23808 29058 23860
rect 29086 23808 29092 23860
rect 29144 23848 29150 23860
rect 29365 23851 29423 23857
rect 29365 23848 29377 23851
rect 29144 23820 29377 23848
rect 29144 23808 29150 23820
rect 29365 23817 29377 23820
rect 29411 23817 29423 23851
rect 29365 23811 29423 23817
rect 30834 23808 30840 23860
rect 30892 23808 30898 23860
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23780 25191 23783
rect 25590 23780 25596 23792
rect 25179 23752 25596 23780
rect 25179 23749 25191 23752
rect 25133 23743 25191 23749
rect 25590 23740 25596 23752
rect 25648 23740 25654 23792
rect 27341 23783 27399 23789
rect 27341 23749 27353 23783
rect 27387 23780 27399 23783
rect 27430 23780 27436 23792
rect 27387 23752 27436 23780
rect 27387 23749 27399 23752
rect 27341 23743 27399 23749
rect 27430 23740 27436 23752
rect 27488 23780 27494 23792
rect 27525 23783 27583 23789
rect 27525 23780 27537 23783
rect 27488 23752 27537 23780
rect 27488 23740 27494 23752
rect 27525 23749 27537 23752
rect 27571 23749 27583 23783
rect 27525 23743 27583 23749
rect 27798 23740 27804 23792
rect 27856 23780 27862 23792
rect 28350 23780 28356 23792
rect 27856 23752 28356 23780
rect 27856 23740 27862 23752
rect 28350 23740 28356 23752
rect 28408 23740 28414 23792
rect 24903 23684 24992 23712
rect 27617 23715 27675 23721
rect 24903 23681 24915 23684
rect 24857 23675 24915 23681
rect 27617 23681 27629 23715
rect 27663 23681 27675 23715
rect 27617 23675 27675 23681
rect 28537 23715 28595 23721
rect 28537 23681 28549 23715
rect 28583 23681 28595 23715
rect 28537 23675 28595 23681
rect 27632 23644 27660 23675
rect 27982 23644 27988 23656
rect 22572 23616 27988 23644
rect 22373 23607 22431 23613
rect 27982 23604 27988 23616
rect 28040 23644 28046 23656
rect 28552 23644 28580 23675
rect 28040 23616 28580 23644
rect 28040 23604 28046 23616
rect 21744 23548 22094 23576
rect 21085 23539 21143 23545
rect 21266 23508 21272 23520
rect 20456 23480 21272 23508
rect 19889 23471 19947 23477
rect 21266 23468 21272 23480
rect 21324 23508 21330 23520
rect 22738 23508 22744 23520
rect 21324 23480 22744 23508
rect 21324 23468 21330 23480
rect 22738 23468 22744 23480
rect 22796 23468 22802 23520
rect 22833 23511 22891 23517
rect 22833 23477 22845 23511
rect 22879 23508 22891 23511
rect 23014 23508 23020 23520
rect 22879 23480 23020 23508
rect 22879 23477 22891 23480
rect 22833 23471 22891 23477
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 23198 23468 23204 23520
rect 23256 23508 23262 23520
rect 23569 23511 23627 23517
rect 23569 23508 23581 23511
rect 23256 23480 23581 23508
rect 23256 23468 23262 23480
rect 23569 23477 23581 23480
rect 23615 23477 23627 23511
rect 23569 23471 23627 23477
rect 24302 23468 24308 23520
rect 24360 23508 24366 23520
rect 24397 23511 24455 23517
rect 24397 23508 24409 23511
rect 24360 23480 24409 23508
rect 24360 23468 24366 23480
rect 24397 23477 24409 23480
rect 24443 23477 24455 23511
rect 24397 23471 24455 23477
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 25317 23511 25375 23517
rect 25317 23508 25329 23511
rect 24912 23480 25329 23508
rect 24912 23468 24918 23480
rect 25317 23477 25329 23480
rect 25363 23477 25375 23511
rect 25317 23471 25375 23477
rect 27157 23511 27215 23517
rect 27157 23477 27169 23511
rect 27203 23508 27215 23511
rect 27246 23508 27252 23520
rect 27203 23480 27252 23508
rect 27203 23477 27215 23480
rect 27157 23471 27215 23477
rect 27246 23468 27252 23480
rect 27304 23508 27310 23520
rect 27522 23508 27528 23520
rect 27304 23480 27528 23508
rect 27304 23468 27310 23480
rect 27522 23468 27528 23480
rect 27580 23468 27586 23520
rect 28552 23508 28580 23616
rect 28644 23576 28672 23808
rect 28736 23712 28764 23808
rect 28813 23715 28871 23721
rect 28813 23712 28825 23715
rect 28736 23684 28825 23712
rect 28813 23681 28825 23684
rect 28859 23681 28871 23715
rect 28920 23712 28948 23808
rect 29196 23752 29592 23780
rect 28997 23715 29055 23721
rect 28997 23712 29009 23715
rect 28920 23684 29009 23712
rect 28813 23675 28871 23681
rect 28997 23681 29009 23684
rect 29043 23681 29055 23715
rect 28997 23675 29055 23681
rect 29086 23672 29092 23724
rect 29144 23672 29150 23724
rect 28721 23647 28779 23653
rect 28721 23613 28733 23647
rect 28767 23644 28779 23647
rect 29196 23644 29224 23752
rect 29273 23715 29331 23721
rect 29273 23681 29285 23715
rect 29319 23681 29331 23715
rect 29273 23675 29331 23681
rect 28767 23616 29224 23644
rect 28767 23613 28779 23616
rect 28721 23607 28779 23613
rect 29089 23579 29147 23585
rect 29089 23576 29101 23579
rect 28644 23548 29101 23576
rect 29089 23545 29101 23548
rect 29135 23545 29147 23579
rect 29089 23539 29147 23545
rect 29288 23508 29316 23675
rect 29362 23672 29368 23724
rect 29420 23672 29426 23724
rect 29564 23721 29592 23752
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23681 29607 23715
rect 30745 23715 30803 23721
rect 30745 23712 30757 23715
rect 29549 23675 29607 23681
rect 30668 23684 30757 23712
rect 30668 23520 30696 23684
rect 30745 23681 30757 23684
rect 30791 23681 30803 23715
rect 30745 23675 30803 23681
rect 28552 23480 29316 23508
rect 30650 23468 30656 23520
rect 30708 23468 30714 23520
rect 1104 23418 35248 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 35248 23418
rect 1104 23344 35248 23366
rect 3418 23264 3424 23316
rect 3476 23264 3482 23316
rect 4525 23307 4583 23313
rect 4525 23273 4537 23307
rect 4571 23304 4583 23307
rect 4706 23304 4712 23316
rect 4571 23276 4712 23304
rect 4571 23273 4583 23276
rect 4525 23267 4583 23273
rect 4706 23264 4712 23276
rect 4764 23264 4770 23316
rect 8294 23264 8300 23316
rect 8352 23264 8358 23316
rect 8846 23264 8852 23316
rect 8904 23304 8910 23316
rect 13817 23307 13875 23313
rect 8904 23276 9168 23304
rect 8904 23264 8910 23276
rect 1670 23128 1676 23180
rect 1728 23128 1734 23180
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 1412 22964 1440 23060
rect 2222 22992 2228 23044
rect 2280 22992 2286 23044
rect 3436 23032 3464 23264
rect 4154 23196 4160 23248
rect 4212 23236 4218 23248
rect 4249 23239 4307 23245
rect 4249 23236 4261 23239
rect 4212 23208 4261 23236
rect 4212 23196 4218 23208
rect 4249 23205 4261 23208
rect 4295 23205 4307 23239
rect 4249 23199 4307 23205
rect 4264 23100 4292 23199
rect 5258 23128 5264 23180
rect 5316 23128 5322 23180
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23168 6423 23171
rect 6638 23168 6644 23180
rect 6411 23140 6644 23168
rect 6411 23137 6423 23140
rect 6365 23131 6423 23137
rect 6638 23128 6644 23140
rect 6696 23128 6702 23180
rect 9140 23177 9168 23276
rect 13817 23273 13829 23307
rect 13863 23304 13875 23307
rect 13906 23304 13912 23316
rect 13863 23276 13912 23304
rect 13863 23273 13875 23276
rect 13817 23267 13875 23273
rect 13906 23264 13912 23276
rect 13964 23304 13970 23316
rect 14366 23304 14372 23316
rect 13964 23276 14372 23304
rect 13964 23264 13970 23276
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 15105 23307 15163 23313
rect 15105 23273 15117 23307
rect 15151 23304 15163 23307
rect 15286 23304 15292 23316
rect 15151 23276 15292 23304
rect 15151 23273 15163 23276
rect 15105 23267 15163 23273
rect 15286 23264 15292 23276
rect 15344 23304 15350 23316
rect 15746 23304 15752 23316
rect 15344 23276 15752 23304
rect 15344 23264 15350 23276
rect 15746 23264 15752 23276
rect 15804 23264 15810 23316
rect 16209 23307 16267 23313
rect 16209 23273 16221 23307
rect 16255 23304 16267 23307
rect 19426 23304 19432 23316
rect 16255 23276 19432 23304
rect 16255 23273 16267 23276
rect 16209 23267 16267 23273
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 19705 23307 19763 23313
rect 19705 23273 19717 23307
rect 19751 23304 19763 23307
rect 19978 23304 19984 23316
rect 19751 23276 19984 23304
rect 19751 23273 19763 23276
rect 19705 23267 19763 23273
rect 19978 23264 19984 23276
rect 20036 23264 20042 23316
rect 20165 23307 20223 23313
rect 20165 23273 20177 23307
rect 20211 23304 20223 23307
rect 20254 23304 20260 23316
rect 20211 23276 20260 23304
rect 20211 23273 20223 23276
rect 20165 23267 20223 23273
rect 20254 23264 20260 23276
rect 20312 23264 20318 23316
rect 21818 23264 21824 23316
rect 21876 23304 21882 23316
rect 22005 23307 22063 23313
rect 22005 23304 22017 23307
rect 21876 23276 22017 23304
rect 21876 23264 21882 23276
rect 22005 23273 22017 23276
rect 22051 23273 22063 23307
rect 22005 23267 22063 23273
rect 22094 23264 22100 23316
rect 22152 23304 22158 23316
rect 22189 23307 22247 23313
rect 22189 23304 22201 23307
rect 22152 23276 22201 23304
rect 22152 23264 22158 23276
rect 22189 23273 22201 23276
rect 22235 23273 22247 23307
rect 22189 23267 22247 23273
rect 22281 23307 22339 23313
rect 22281 23273 22293 23307
rect 22327 23304 22339 23307
rect 22462 23304 22468 23316
rect 22327 23276 22468 23304
rect 22327 23273 22339 23276
rect 22281 23267 22339 23273
rect 15657 23239 15715 23245
rect 15657 23205 15669 23239
rect 15703 23236 15715 23239
rect 17589 23239 17647 23245
rect 15703 23208 17264 23236
rect 15703 23205 15715 23208
rect 15657 23199 15715 23205
rect 8113 23171 8171 23177
rect 8113 23137 8125 23171
rect 8159 23168 8171 23171
rect 9125 23171 9183 23177
rect 8159 23140 8984 23168
rect 8159 23137 8171 23140
rect 8113 23131 8171 23137
rect 4433 23103 4491 23109
rect 4433 23100 4445 23103
rect 4264 23072 4445 23100
rect 4433 23069 4445 23072
rect 4479 23069 4491 23103
rect 4433 23063 4491 23069
rect 4798 23060 4804 23112
rect 4856 23100 4862 23112
rect 5169 23103 5227 23109
rect 5169 23100 5181 23103
rect 4856 23072 5181 23100
rect 4856 23060 4862 23072
rect 5169 23069 5181 23072
rect 5215 23100 5227 23103
rect 5442 23100 5448 23112
rect 5215 23072 5448 23100
rect 5215 23069 5227 23072
rect 5169 23063 5227 23069
rect 5442 23060 5448 23072
rect 5500 23060 5506 23112
rect 8202 23060 8208 23112
rect 8260 23100 8266 23112
rect 8956 23109 8984 23140
rect 9125 23137 9137 23171
rect 9171 23137 9183 23171
rect 9125 23131 9183 23137
rect 15013 23171 15071 23177
rect 15013 23137 15025 23171
rect 15059 23168 15071 23171
rect 15378 23168 15384 23180
rect 15059 23140 15384 23168
rect 15059 23137 15071 23140
rect 15013 23131 15071 23137
rect 15378 23128 15384 23140
rect 15436 23168 15442 23180
rect 15841 23171 15899 23177
rect 15841 23168 15853 23171
rect 15436 23140 15853 23168
rect 15436 23128 15442 23140
rect 15841 23137 15853 23140
rect 15887 23137 15899 23171
rect 15841 23131 15899 23137
rect 17126 23128 17132 23180
rect 17184 23128 17190 23180
rect 8389 23103 8447 23109
rect 8389 23100 8401 23103
rect 8260 23072 8401 23100
rect 8260 23060 8266 23072
rect 8389 23069 8401 23072
rect 8435 23100 8447 23103
rect 8665 23103 8723 23109
rect 8665 23100 8677 23103
rect 8435 23072 8677 23100
rect 8435 23069 8447 23072
rect 8389 23063 8447 23069
rect 8665 23069 8677 23072
rect 8711 23069 8723 23103
rect 8665 23063 8723 23069
rect 8941 23103 8999 23109
rect 8941 23069 8953 23103
rect 8987 23069 8999 23103
rect 8941 23063 8999 23069
rect 10042 23060 10048 23112
rect 10100 23060 10106 23112
rect 10226 23060 10232 23112
rect 10284 23060 10290 23112
rect 15562 23109 15568 23112
rect 15532 23103 15568 23109
rect 15532 23069 15544 23103
rect 15620 23100 15626 23112
rect 17236 23109 17264 23208
rect 17589 23205 17601 23239
rect 17635 23236 17647 23239
rect 21085 23239 21143 23245
rect 17635 23208 18276 23236
rect 17635 23205 17647 23208
rect 17589 23199 17647 23205
rect 18248 23177 18276 23208
rect 21085 23205 21097 23239
rect 21131 23236 21143 23239
rect 22296 23236 22324 23267
rect 22462 23264 22468 23276
rect 22520 23264 22526 23316
rect 22557 23307 22615 23313
rect 22557 23273 22569 23307
rect 22603 23304 22615 23307
rect 22646 23304 22652 23316
rect 22603 23276 22652 23304
rect 22603 23273 22615 23276
rect 22557 23267 22615 23273
rect 22646 23264 22652 23276
rect 22704 23264 22710 23316
rect 23198 23264 23204 23316
rect 23256 23304 23262 23316
rect 23385 23307 23443 23313
rect 23385 23304 23397 23307
rect 23256 23276 23397 23304
rect 23256 23264 23262 23276
rect 23385 23273 23397 23276
rect 23431 23273 23443 23307
rect 23385 23267 23443 23273
rect 24394 23264 24400 23316
rect 24452 23304 24458 23316
rect 24489 23307 24547 23313
rect 24489 23304 24501 23307
rect 24452 23276 24501 23304
rect 24452 23264 24458 23276
rect 24489 23273 24501 23276
rect 24535 23273 24547 23307
rect 24489 23267 24547 23273
rect 24581 23307 24639 23313
rect 24581 23273 24593 23307
rect 24627 23304 24639 23307
rect 24854 23304 24860 23316
rect 24627 23276 24860 23304
rect 24627 23273 24639 23276
rect 24581 23267 24639 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 21131 23208 22324 23236
rect 23676 23208 25084 23236
rect 21131 23205 21143 23208
rect 21085 23199 21143 23205
rect 21468 23177 21496 23208
rect 18233 23171 18291 23177
rect 18233 23137 18245 23171
rect 18279 23137 18291 23171
rect 18233 23131 18291 23137
rect 20809 23171 20867 23177
rect 20809 23137 20821 23171
rect 20855 23168 20867 23171
rect 21453 23171 21511 23177
rect 20855 23140 21312 23168
rect 20855 23137 20867 23140
rect 20809 23131 20867 23137
rect 15933 23103 15991 23109
rect 15933 23100 15945 23103
rect 15620 23072 15945 23100
rect 15532 23063 15568 23069
rect 15562 23060 15568 23063
rect 15620 23060 15626 23072
rect 15933 23069 15945 23072
rect 15979 23069 15991 23103
rect 15933 23063 15991 23069
rect 17221 23103 17279 23109
rect 17221 23069 17233 23103
rect 17267 23069 17279 23103
rect 17221 23063 17279 23069
rect 11152 23044 11204 23050
rect 4706 23032 4712 23044
rect 3068 23004 3464 23032
rect 4172 23004 4712 23032
rect 2590 22964 2596 22976
rect 1412 22936 2596 22964
rect 2590 22924 2596 22936
rect 2648 22964 2654 22976
rect 3068 22964 3096 23004
rect 2648 22936 3096 22964
rect 3145 22967 3203 22973
rect 2648 22924 2654 22936
rect 3145 22933 3157 22967
rect 3191 22964 3203 22967
rect 4172 22964 4200 23004
rect 4706 22992 4712 23004
rect 4764 22992 4770 23044
rect 6641 23035 6699 23041
rect 6641 23032 6653 23035
rect 5552 23004 6653 23032
rect 5552 22973 5580 23004
rect 6641 23001 6653 23004
rect 6687 23001 6699 23035
rect 6641 22995 6699 23001
rect 7650 22992 7656 23044
rect 7708 22992 7714 23044
rect 15194 22992 15200 23044
rect 15252 22992 15258 23044
rect 11152 22986 11204 22992
rect 3191 22936 4200 22964
rect 5537 22967 5595 22973
rect 3191 22933 3203 22936
rect 3145 22927 3203 22933
rect 5537 22933 5549 22967
rect 5583 22933 5595 22967
rect 5537 22927 5595 22933
rect 12710 22924 12716 22976
rect 12768 22964 12774 22976
rect 13081 22967 13139 22973
rect 13081 22964 13093 22967
rect 12768 22936 13093 22964
rect 12768 22924 12774 22936
rect 13081 22933 13093 22936
rect 13127 22933 13139 22967
rect 13081 22927 13139 22933
rect 14366 22924 14372 22976
rect 14424 22924 14430 22976
rect 15212 22964 15240 22992
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 15212 22936 15485 22964
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 18248 22964 18276 23131
rect 18414 23060 18420 23112
rect 18472 23100 18478 23112
rect 18601 23103 18659 23109
rect 18472 23072 18552 23100
rect 18472 23060 18478 23072
rect 18524 23032 18552 23072
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 19521 23103 19579 23109
rect 19521 23100 19533 23103
rect 18647 23072 19533 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 19521 23069 19533 23072
rect 19567 23069 19579 23103
rect 19521 23063 19579 23069
rect 20717 23103 20775 23109
rect 20717 23069 20729 23103
rect 20763 23069 20775 23103
rect 20717 23063 20775 23069
rect 20901 23103 20959 23109
rect 20901 23069 20913 23103
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 18693 23035 18751 23041
rect 18693 23032 18705 23035
rect 18524 23004 18705 23032
rect 18693 23001 18705 23004
rect 18739 23001 18751 23035
rect 18693 22995 18751 23001
rect 18877 23035 18935 23041
rect 18877 23001 18889 23035
rect 18923 23001 18935 23035
rect 18877 22995 18935 23001
rect 19061 23035 19119 23041
rect 19061 23001 19073 23035
rect 19107 23032 19119 23035
rect 19245 23035 19303 23041
rect 19245 23032 19257 23035
rect 19107 23004 19257 23032
rect 19107 23001 19119 23004
rect 19061 22995 19119 23001
rect 19245 23001 19257 23004
rect 19291 23001 19303 23035
rect 19245 22995 19303 23001
rect 18598 22964 18604 22976
rect 18248 22936 18604 22964
rect 15473 22927 15531 22933
rect 18598 22924 18604 22936
rect 18656 22964 18662 22976
rect 18892 22964 18920 22995
rect 18656 22936 18920 22964
rect 18656 22924 18662 22936
rect 19334 22924 19340 22976
rect 19392 22924 19398 22976
rect 20625 22967 20683 22973
rect 20625 22933 20637 22967
rect 20671 22964 20683 22967
rect 20732 22964 20760 23063
rect 20916 23032 20944 23063
rect 20990 23060 20996 23112
rect 21048 23060 21054 23112
rect 21082 23060 21088 23112
rect 21140 23100 21146 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 21140 23072 21189 23100
rect 21140 23060 21146 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21284 23100 21312 23140
rect 21453 23137 21465 23171
rect 21499 23137 21511 23171
rect 23014 23168 23020 23180
rect 22112 23147 23020 23168
rect 21453 23131 21511 23137
rect 22097 23141 23020 23147
rect 21637 23103 21695 23109
rect 21637 23100 21649 23103
rect 21284 23072 21649 23100
rect 21177 23063 21235 23069
rect 21637 23069 21649 23072
rect 21683 23069 21695 23103
rect 22097 23107 22109 23141
rect 22143 23140 23020 23141
rect 22143 23107 22155 23140
rect 23014 23128 23020 23140
rect 23072 23128 23078 23180
rect 22097 23101 22155 23107
rect 22373 23103 22431 23109
rect 21637 23063 21695 23069
rect 22112 23032 22140 23101
rect 22373 23069 22385 23103
rect 22419 23069 22431 23103
rect 22373 23063 22431 23069
rect 22741 23103 22799 23109
rect 22741 23069 22753 23103
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 20916 23004 22140 23032
rect 21450 22964 21456 22976
rect 20671 22936 21456 22964
rect 20671 22933 20683 22936
rect 20625 22927 20683 22933
rect 21450 22924 21456 22936
rect 21508 22924 21514 22976
rect 21542 22924 21548 22976
rect 21600 22924 21606 22976
rect 22388 22964 22416 23063
rect 22756 23032 22784 23063
rect 22830 23060 22836 23112
rect 22888 23060 22894 23112
rect 23106 23060 23112 23112
rect 23164 23060 23170 23112
rect 23676 23100 23704 23208
rect 23753 23171 23811 23177
rect 23753 23137 23765 23171
rect 23799 23168 23811 23171
rect 24397 23171 24455 23177
rect 24397 23168 24409 23171
rect 23799 23140 24409 23168
rect 23799 23137 23811 23140
rect 23753 23131 23811 23137
rect 24397 23137 24409 23140
rect 24443 23137 24455 23171
rect 24397 23131 24455 23137
rect 23937 23103 23995 23109
rect 23937 23100 23949 23103
rect 23676 23072 23949 23100
rect 23937 23069 23949 23072
rect 23983 23100 23995 23103
rect 24026 23100 24032 23112
rect 23983 23072 24032 23100
rect 23983 23069 23995 23072
rect 23937 23063 23995 23069
rect 24026 23060 24032 23072
rect 24084 23060 24090 23112
rect 24213 23103 24271 23109
rect 24213 23069 24225 23103
rect 24259 23100 24271 23103
rect 24302 23100 24308 23112
rect 24259 23072 24308 23100
rect 24259 23069 24271 23072
rect 24213 23063 24271 23069
rect 24302 23060 24308 23072
rect 24360 23060 24366 23112
rect 24486 23060 24492 23112
rect 24544 23100 24550 23112
rect 24673 23103 24731 23109
rect 24673 23100 24685 23103
rect 24544 23072 24685 23100
rect 24544 23060 24550 23072
rect 24673 23069 24685 23072
rect 24719 23069 24731 23103
rect 24673 23063 24731 23069
rect 24762 23060 24768 23112
rect 24820 23060 24826 23112
rect 24854 23060 24860 23112
rect 24912 23060 24918 23112
rect 25056 23109 25084 23208
rect 25774 23128 25780 23180
rect 25832 23128 25838 23180
rect 34057 23171 34115 23177
rect 34057 23137 34069 23171
rect 34103 23168 34115 23171
rect 34103 23140 34652 23168
rect 34103 23137 34115 23140
rect 34057 23131 34115 23137
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23069 25099 23103
rect 25041 23063 25099 23069
rect 34517 23103 34575 23109
rect 34517 23069 34529 23103
rect 34563 23069 34575 23103
rect 34517 23063 34575 23069
rect 22756 23004 22876 23032
rect 22848 22976 22876 23004
rect 22922 22992 22928 23044
rect 22980 23032 22986 23044
rect 23201 23035 23259 23041
rect 23201 23032 23213 23035
rect 22980 23004 23213 23032
rect 22980 22992 22986 23004
rect 23201 23001 23213 23004
rect 23247 23001 23259 23035
rect 23201 22995 23259 23001
rect 24121 23035 24179 23041
rect 24121 23001 24133 23035
rect 24167 23032 24179 23035
rect 24780 23032 24808 23060
rect 24167 23004 24808 23032
rect 24167 23001 24179 23004
rect 24121 22995 24179 23001
rect 22462 22964 22468 22976
rect 22388 22936 22468 22964
rect 22462 22924 22468 22936
rect 22520 22964 22526 22976
rect 22738 22964 22744 22976
rect 22520 22936 22744 22964
rect 22520 22924 22526 22936
rect 22738 22924 22744 22936
rect 22796 22924 22802 22976
rect 22830 22924 22836 22976
rect 22888 22964 22894 22976
rect 23401 22967 23459 22973
rect 23401 22964 23413 22967
rect 22888 22936 23413 22964
rect 22888 22924 22894 22936
rect 23401 22933 23413 22936
rect 23447 22933 23459 22967
rect 23401 22927 23459 22933
rect 23569 22967 23627 22973
rect 23569 22933 23581 22967
rect 23615 22964 23627 22967
rect 24486 22964 24492 22976
rect 23615 22936 24492 22964
rect 23615 22933 23627 22936
rect 23569 22927 23627 22933
rect 24486 22924 24492 22936
rect 24544 22924 24550 22976
rect 34532 22964 34560 23063
rect 34624 23044 34652 23140
rect 34606 22992 34612 23044
rect 34664 22992 34670 23044
rect 34532 22936 35296 22964
rect 1104 22874 35236 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 35236 22874
rect 1104 22800 35236 22822
rect 2222 22720 2228 22772
rect 2280 22720 2286 22772
rect 7561 22763 7619 22769
rect 7561 22729 7573 22763
rect 7607 22760 7619 22763
rect 7650 22760 7656 22772
rect 7607 22732 7656 22760
rect 7607 22729 7619 22732
rect 7561 22723 7619 22729
rect 7650 22720 7656 22732
rect 7708 22720 7714 22772
rect 8113 22763 8171 22769
rect 8113 22729 8125 22763
rect 8159 22760 8171 22763
rect 8202 22760 8208 22772
rect 8159 22732 8208 22760
rect 8159 22729 8171 22732
rect 8113 22723 8171 22729
rect 2866 22652 2872 22704
rect 2924 22652 2930 22704
rect 3878 22652 3884 22704
rect 3936 22652 3942 22704
rect 2133 22627 2191 22633
rect 2133 22593 2145 22627
rect 2179 22593 2191 22627
rect 2133 22587 2191 22593
rect 7377 22627 7435 22633
rect 7377 22593 7389 22627
rect 7423 22624 7435 22627
rect 7653 22627 7711 22633
rect 7653 22624 7665 22627
rect 7423 22596 7665 22624
rect 7423 22593 7435 22596
rect 7377 22587 7435 22593
rect 7653 22593 7665 22596
rect 7699 22624 7711 22627
rect 8128 22624 8156 22723
rect 8202 22720 8208 22732
rect 8260 22720 8266 22772
rect 10965 22763 11023 22769
rect 10965 22729 10977 22763
rect 11011 22760 11023 22763
rect 12434 22760 12440 22772
rect 11011 22732 12440 22760
rect 11011 22729 11023 22732
rect 10965 22723 11023 22729
rect 7699 22596 8156 22624
rect 9033 22627 9091 22633
rect 7699 22593 7711 22596
rect 7653 22587 7711 22593
rect 9033 22593 9045 22627
rect 9079 22624 9091 22627
rect 9674 22624 9680 22636
rect 9079 22596 9680 22624
rect 9079 22593 9091 22596
rect 9033 22587 9091 22593
rect 2041 22423 2099 22429
rect 2041 22389 2053 22423
rect 2087 22420 2099 22423
rect 2148 22420 2176 22587
rect 9674 22584 9680 22596
rect 9732 22624 9738 22636
rect 9861 22627 9919 22633
rect 9861 22624 9873 22627
rect 9732 22596 9873 22624
rect 9732 22584 9738 22596
rect 9861 22593 9873 22596
rect 9907 22593 9919 22627
rect 9861 22587 9919 22593
rect 10137 22627 10195 22633
rect 10137 22593 10149 22627
rect 10183 22624 10195 22627
rect 10318 22624 10324 22636
rect 10183 22596 10324 22624
rect 10183 22593 10195 22596
rect 10137 22587 10195 22593
rect 2590 22516 2596 22568
rect 2648 22556 2654 22568
rect 4341 22559 4399 22565
rect 2648 22528 3924 22556
rect 2648 22516 2654 22528
rect 2682 22420 2688 22432
rect 2087 22392 2688 22420
rect 2087 22389 2099 22392
rect 2041 22383 2099 22389
rect 2682 22380 2688 22392
rect 2740 22380 2746 22432
rect 3896 22420 3924 22528
rect 4341 22525 4353 22559
rect 4387 22556 4399 22559
rect 4798 22556 4804 22568
rect 4387 22528 4804 22556
rect 4387 22525 4399 22528
rect 4341 22519 4399 22525
rect 4798 22516 4804 22528
rect 4856 22516 4862 22568
rect 9876 22556 9904 22587
rect 10318 22584 10324 22596
rect 10376 22624 10382 22636
rect 10980 22624 11008 22723
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 14090 22760 14096 22772
rect 13832 22732 14096 22760
rect 12452 22692 12480 22720
rect 13541 22695 13599 22701
rect 12452 22664 12848 22692
rect 12710 22624 12716 22636
rect 10376 22596 11008 22624
rect 11992 22596 12716 22624
rect 10376 22584 10382 22596
rect 11882 22556 11888 22568
rect 9876 22528 11888 22556
rect 11882 22516 11888 22528
rect 11940 22516 11946 22568
rect 9953 22491 10011 22497
rect 9953 22457 9965 22491
rect 9999 22488 10011 22491
rect 10042 22488 10048 22500
rect 9999 22460 10048 22488
rect 9999 22457 10011 22460
rect 9953 22451 10011 22457
rect 10042 22448 10048 22460
rect 10100 22448 10106 22500
rect 10778 22488 10784 22500
rect 10520 22460 10784 22488
rect 4709 22423 4767 22429
rect 4709 22420 4721 22423
rect 3896 22392 4721 22420
rect 4709 22389 4721 22392
rect 4755 22420 4767 22423
rect 4890 22420 4896 22432
rect 4755 22392 4896 22420
rect 4755 22389 4767 22392
rect 4709 22383 4767 22389
rect 4890 22380 4896 22392
rect 4948 22420 4954 22432
rect 6638 22420 6644 22432
rect 4948 22392 6644 22420
rect 4948 22380 4954 22392
rect 6638 22380 6644 22392
rect 6696 22380 6702 22432
rect 8665 22423 8723 22429
rect 8665 22389 8677 22423
rect 8711 22420 8723 22423
rect 9306 22420 9312 22432
rect 8711 22392 9312 22420
rect 8711 22389 8723 22392
rect 8665 22383 8723 22389
rect 9306 22380 9312 22392
rect 9364 22380 9370 22432
rect 9401 22423 9459 22429
rect 9401 22389 9413 22423
rect 9447 22420 9459 22423
rect 9490 22420 9496 22432
rect 9447 22392 9496 22420
rect 9447 22389 9459 22392
rect 9401 22383 9459 22389
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 9766 22380 9772 22432
rect 9824 22420 9830 22432
rect 10520 22420 10548 22460
rect 10778 22448 10784 22460
rect 10836 22488 10842 22500
rect 11992 22497 12020 22596
rect 12710 22584 12716 22596
rect 12768 22584 12774 22636
rect 12820 22633 12848 22664
rect 13541 22661 13553 22695
rect 13587 22661 13599 22695
rect 13541 22655 13599 22661
rect 13633 22695 13691 22701
rect 13633 22661 13645 22695
rect 13679 22692 13691 22695
rect 13832 22692 13860 22732
rect 14090 22720 14096 22732
rect 14148 22760 14154 22772
rect 14274 22760 14280 22772
rect 14148 22732 14280 22760
rect 14148 22720 14154 22732
rect 14274 22720 14280 22732
rect 14332 22720 14338 22772
rect 14458 22720 14464 22772
rect 14516 22760 14522 22772
rect 15105 22763 15163 22769
rect 15105 22760 15117 22763
rect 14516 22732 15117 22760
rect 14516 22720 14522 22732
rect 15105 22729 15117 22732
rect 15151 22729 15163 22763
rect 15105 22723 15163 22729
rect 15381 22763 15439 22769
rect 15381 22729 15393 22763
rect 15427 22760 15439 22763
rect 15562 22760 15568 22772
rect 15427 22732 15568 22760
rect 15427 22729 15439 22732
rect 15381 22723 15439 22729
rect 13679 22664 13860 22692
rect 13679 22661 13691 22664
rect 13633 22655 13691 22661
rect 12805 22627 12863 22633
rect 12805 22593 12817 22627
rect 12851 22593 12863 22627
rect 12805 22587 12863 22593
rect 13446 22584 13452 22636
rect 13504 22584 13510 22636
rect 12728 22556 12756 22584
rect 13553 22556 13581 22655
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 13740 22614 13829 22624
rect 12728 22528 13581 22556
rect 13648 22596 13829 22614
rect 13648 22586 13768 22596
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 11977 22491 12035 22497
rect 11977 22488 11989 22491
rect 10836 22460 11989 22488
rect 10836 22448 10842 22460
rect 11977 22457 11989 22460
rect 12023 22457 12035 22491
rect 11977 22451 12035 22457
rect 12529 22491 12587 22497
rect 12529 22457 12541 22491
rect 12575 22488 12587 22491
rect 12986 22488 12992 22500
rect 12575 22460 12992 22488
rect 12575 22457 12587 22460
rect 12529 22451 12587 22457
rect 12986 22448 12992 22460
rect 13044 22488 13050 22500
rect 13648 22488 13676 22586
rect 13906 22584 13912 22636
rect 13964 22584 13970 22636
rect 14093 22627 14151 22633
rect 14093 22593 14105 22627
rect 14139 22593 14151 22627
rect 15120 22624 15148 22723
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 15841 22763 15899 22769
rect 15841 22729 15853 22763
rect 15887 22760 15899 22763
rect 17586 22760 17592 22772
rect 15887 22732 17592 22760
rect 15887 22729 15899 22732
rect 15841 22723 15899 22729
rect 15289 22627 15347 22633
rect 15289 22624 15301 22627
rect 15120 22596 15301 22624
rect 14093 22587 14151 22593
rect 15289 22593 15301 22596
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 15473 22627 15531 22633
rect 15473 22593 15485 22627
rect 15519 22624 15531 22627
rect 15856 22624 15884 22723
rect 17586 22720 17592 22732
rect 17644 22720 17650 22772
rect 18598 22720 18604 22772
rect 18656 22720 18662 22772
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 20993 22763 21051 22769
rect 20993 22760 21005 22763
rect 20956 22732 21005 22760
rect 20956 22720 20962 22732
rect 20993 22729 21005 22732
rect 21039 22729 21051 22763
rect 20993 22723 21051 22729
rect 21174 22720 21180 22772
rect 21232 22720 21238 22772
rect 21542 22720 21548 22772
rect 21600 22760 21606 22772
rect 21821 22763 21879 22769
rect 21821 22760 21833 22763
rect 21600 22732 21833 22760
rect 21600 22720 21606 22732
rect 21821 22729 21833 22732
rect 21867 22729 21879 22763
rect 22649 22763 22707 22769
rect 22649 22760 22661 22763
rect 21821 22723 21879 22729
rect 22480 22732 22661 22760
rect 18616 22633 18644 22720
rect 21192 22692 21220 22720
rect 22480 22701 22508 22732
rect 22649 22729 22661 22732
rect 22695 22760 22707 22763
rect 22830 22760 22836 22772
rect 22695 22732 22836 22760
rect 22695 22729 22707 22732
rect 22649 22723 22707 22729
rect 22830 22720 22836 22732
rect 22888 22720 22894 22772
rect 23014 22720 23020 22772
rect 23072 22760 23078 22772
rect 23493 22763 23551 22769
rect 23493 22760 23505 22763
rect 23072 22732 23505 22760
rect 23072 22720 23078 22732
rect 23493 22729 23505 22732
rect 23539 22729 23551 22763
rect 23493 22723 23551 22729
rect 24486 22720 24492 22772
rect 24544 22720 24550 22772
rect 24854 22720 24860 22772
rect 24912 22760 24918 22772
rect 24949 22763 25007 22769
rect 24949 22760 24961 22763
rect 24912 22732 24961 22760
rect 24912 22720 24918 22732
rect 24949 22729 24961 22732
rect 24995 22729 25007 22763
rect 24949 22723 25007 22729
rect 29638 22720 29644 22772
rect 29696 22760 29702 22772
rect 29917 22763 29975 22769
rect 29917 22760 29929 22763
rect 29696 22732 29929 22760
rect 29696 22720 29702 22732
rect 29917 22729 29929 22732
rect 29963 22729 29975 22763
rect 29917 22723 29975 22729
rect 32677 22763 32735 22769
rect 32677 22729 32689 22763
rect 32723 22729 32735 22763
rect 32677 22723 32735 22729
rect 34885 22763 34943 22769
rect 34885 22729 34897 22763
rect 34931 22760 34943 22763
rect 35268 22760 35296 22936
rect 34931 22732 35296 22760
rect 34931 22729 34943 22732
rect 34885 22723 34943 22729
rect 22465 22695 22523 22701
rect 21192 22664 22324 22692
rect 15519 22596 15884 22624
rect 18601 22627 18659 22633
rect 15519 22593 15531 22596
rect 15473 22587 15531 22593
rect 18601 22593 18613 22627
rect 18647 22593 18659 22627
rect 18601 22587 18659 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22624 20775 22627
rect 20990 22624 20996 22636
rect 20763 22596 20996 22624
rect 20763 22593 20775 22596
rect 20717 22587 20775 22593
rect 14108 22556 14136 22587
rect 14182 22556 14188 22568
rect 14108 22528 14188 22556
rect 14182 22516 14188 22528
rect 14240 22556 14246 22568
rect 14366 22556 14372 22568
rect 14240 22528 14372 22556
rect 14240 22516 14246 22528
rect 14366 22516 14372 22528
rect 14424 22556 14430 22568
rect 15488 22556 15516 22587
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22624 22155 22627
rect 22186 22624 22192 22636
rect 22143 22596 22192 22624
rect 22143 22593 22155 22596
rect 22097 22587 22155 22593
rect 14424 22528 15516 22556
rect 14424 22516 14430 22528
rect 18046 22516 18052 22568
rect 18104 22556 18110 22568
rect 18414 22556 18420 22568
rect 18104 22528 18420 22556
rect 18104 22516 18110 22528
rect 18414 22516 18420 22528
rect 18472 22556 18478 22568
rect 18509 22559 18567 22565
rect 18509 22556 18521 22559
rect 18472 22528 18521 22556
rect 18472 22516 18478 22528
rect 18509 22525 18521 22528
rect 18555 22525 18567 22559
rect 18509 22519 18567 22525
rect 21726 22516 21732 22568
rect 21784 22556 21790 22568
rect 22005 22559 22063 22565
rect 22005 22556 22017 22559
rect 21784 22528 22017 22556
rect 21784 22516 21790 22528
rect 22005 22525 22017 22528
rect 22051 22525 22063 22559
rect 22005 22519 22063 22525
rect 14553 22491 14611 22497
rect 14553 22488 14565 22491
rect 13044 22460 13676 22488
rect 13923 22460 14565 22488
rect 13044 22448 13050 22460
rect 9824 22392 10548 22420
rect 9824 22380 9830 22392
rect 10594 22380 10600 22432
rect 10652 22420 10658 22432
rect 11054 22420 11060 22432
rect 10652 22392 11060 22420
rect 10652 22380 10658 22392
rect 11054 22380 11060 22392
rect 11112 22380 11118 22432
rect 13262 22380 13268 22432
rect 13320 22380 13326 22432
rect 13446 22380 13452 22432
rect 13504 22420 13510 22432
rect 13923 22420 13951 22460
rect 14553 22457 14565 22460
rect 14599 22457 14611 22491
rect 14553 22451 14611 22457
rect 18969 22491 19027 22497
rect 18969 22457 18981 22491
rect 19015 22488 19027 22491
rect 19518 22488 19524 22500
rect 19015 22460 19524 22488
rect 19015 22457 19027 22460
rect 18969 22451 19027 22457
rect 19518 22448 19524 22460
rect 19576 22448 19582 22500
rect 21450 22448 21456 22500
rect 21508 22488 21514 22500
rect 21545 22491 21603 22497
rect 21545 22488 21557 22491
rect 21508 22460 21557 22488
rect 21508 22448 21514 22460
rect 21545 22457 21557 22460
rect 21591 22488 21603 22491
rect 22112 22488 22140 22587
rect 22186 22584 22192 22596
rect 22244 22584 22250 22636
rect 22296 22624 22324 22664
rect 22465 22661 22477 22695
rect 22511 22661 22523 22695
rect 22465 22655 22523 22661
rect 23290 22652 23296 22704
rect 23348 22692 23354 22704
rect 23937 22695 23995 22701
rect 23937 22692 23949 22695
rect 23348 22664 23949 22692
rect 23348 22652 23354 22664
rect 23937 22661 23949 22664
rect 23983 22661 23995 22695
rect 23937 22655 23995 22661
rect 22554 22624 22560 22636
rect 22296 22596 22560 22624
rect 22554 22584 22560 22596
rect 22612 22584 22618 22636
rect 22741 22627 22799 22633
rect 22741 22593 22753 22627
rect 22787 22593 22799 22627
rect 22741 22587 22799 22593
rect 22370 22516 22376 22568
rect 22428 22516 22434 22568
rect 22756 22488 22784 22587
rect 22830 22516 22836 22568
rect 22888 22556 22894 22568
rect 23308 22556 23336 22652
rect 24504 22624 24532 22720
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 24504 22596 24593 22624
rect 24581 22593 24593 22596
rect 24627 22593 24639 22627
rect 24581 22587 24639 22593
rect 26234 22584 26240 22636
rect 26292 22624 26298 22636
rect 27709 22627 27767 22633
rect 27709 22624 27721 22627
rect 26292 22596 27721 22624
rect 26292 22584 26298 22596
rect 27709 22593 27721 22596
rect 27755 22624 27767 22627
rect 28442 22624 28448 22636
rect 27755 22596 28448 22624
rect 27755 22593 27767 22596
rect 27709 22587 27767 22593
rect 28442 22584 28448 22596
rect 28500 22584 28506 22636
rect 29932 22624 29960 22723
rect 30926 22652 30932 22704
rect 30984 22652 30990 22704
rect 32692 22692 32720 22723
rect 33413 22695 33471 22701
rect 33413 22692 33425 22695
rect 32692 22664 33425 22692
rect 33413 22661 33425 22664
rect 33459 22661 33471 22695
rect 33413 22655 33471 22661
rect 34146 22652 34152 22704
rect 34204 22652 34210 22704
rect 30101 22627 30159 22633
rect 30101 22624 30113 22627
rect 29932 22596 30113 22624
rect 30101 22593 30113 22596
rect 30147 22593 30159 22627
rect 32030 22624 32036 22636
rect 30101 22587 30159 22593
rect 31864 22596 32036 22624
rect 24489 22559 24547 22565
rect 24489 22556 24501 22559
rect 22888 22528 23336 22556
rect 23676 22528 24501 22556
rect 22888 22516 22894 22528
rect 23676 22497 23704 22528
rect 24489 22525 24501 22528
rect 24535 22556 24547 22559
rect 25038 22556 25044 22568
rect 24535 22528 25044 22556
rect 24535 22525 24547 22528
rect 24489 22519 24547 22525
rect 25038 22516 25044 22528
rect 25096 22516 25102 22568
rect 27614 22516 27620 22568
rect 27672 22556 27678 22568
rect 27985 22559 28043 22565
rect 27985 22556 27997 22559
rect 27672 22528 27997 22556
rect 27672 22516 27678 22528
rect 27985 22525 27997 22528
rect 28031 22525 28043 22559
rect 27985 22519 28043 22525
rect 30374 22516 30380 22568
rect 30432 22516 30438 22568
rect 31864 22565 31892 22596
rect 32030 22584 32036 22596
rect 32088 22624 32094 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 32088 22596 32321 22624
rect 32088 22584 32094 22596
rect 32309 22593 32321 22596
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 32490 22584 32496 22636
rect 32548 22624 32554 22636
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 32548 22596 32781 22624
rect 32548 22584 32554 22596
rect 32769 22593 32781 22596
rect 32815 22593 32827 22627
rect 32769 22587 32827 22593
rect 32950 22584 32956 22636
rect 33008 22584 33014 22636
rect 31849 22559 31907 22565
rect 31849 22525 31861 22559
rect 31895 22525 31907 22559
rect 31849 22519 31907 22525
rect 32401 22559 32459 22565
rect 32401 22525 32413 22559
rect 32447 22556 32459 22559
rect 32861 22559 32919 22565
rect 32861 22556 32873 22559
rect 32447 22528 32873 22556
rect 32447 22525 32459 22528
rect 32401 22519 32459 22525
rect 32861 22525 32873 22528
rect 32907 22525 32919 22559
rect 32861 22519 32919 22525
rect 23661 22491 23719 22497
rect 21591 22460 23152 22488
rect 21591 22457 21603 22460
rect 21545 22451 21603 22457
rect 23124 22432 23152 22460
rect 23661 22457 23673 22491
rect 23707 22457 23719 22491
rect 23661 22451 23719 22457
rect 32582 22448 32588 22500
rect 32640 22488 32646 22500
rect 32968 22488 32996 22584
rect 33137 22559 33195 22565
rect 33137 22525 33149 22559
rect 33183 22525 33195 22559
rect 33137 22519 33195 22525
rect 32640 22460 32996 22488
rect 32640 22448 32646 22460
rect 13504 22392 13951 22420
rect 13504 22380 13510 22392
rect 14274 22380 14280 22432
rect 14332 22380 14338 22432
rect 23106 22380 23112 22432
rect 23164 22380 23170 22432
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 23477 22423 23535 22429
rect 23477 22420 23489 22423
rect 23440 22392 23489 22420
rect 23440 22380 23446 22392
rect 23477 22389 23489 22392
rect 23523 22389 23535 22423
rect 23477 22383 23535 22389
rect 27522 22380 27528 22432
rect 27580 22380 27586 22432
rect 27890 22380 27896 22432
rect 27948 22380 27954 22432
rect 32674 22380 32680 22432
rect 32732 22420 32738 22432
rect 33152 22420 33180 22519
rect 32732 22392 33180 22420
rect 32732 22380 32738 22392
rect 1104 22330 35248 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 35248 22330
rect 1104 22256 35248 22278
rect 3878 22176 3884 22228
rect 3936 22176 3942 22228
rect 4801 22219 4859 22225
rect 4801 22185 4813 22219
rect 4847 22216 4859 22219
rect 4890 22216 4896 22228
rect 4847 22188 4896 22216
rect 4847 22185 4859 22188
rect 4801 22179 4859 22185
rect 4890 22176 4896 22188
rect 4948 22176 4954 22228
rect 5169 22219 5227 22225
rect 5169 22185 5181 22219
rect 5215 22216 5227 22219
rect 5258 22216 5264 22228
rect 5215 22188 5264 22216
rect 5215 22185 5227 22188
rect 5169 22179 5227 22185
rect 5258 22176 5264 22188
rect 5316 22176 5322 22228
rect 5442 22176 5448 22228
rect 5500 22216 5506 22228
rect 5813 22219 5871 22225
rect 5813 22216 5825 22219
rect 5500 22188 5825 22216
rect 5500 22176 5506 22188
rect 5813 22185 5825 22188
rect 5859 22185 5871 22219
rect 5813 22179 5871 22185
rect 10413 22219 10471 22225
rect 10413 22185 10425 22219
rect 10459 22216 10471 22219
rect 13998 22216 14004 22228
rect 10459 22188 14004 22216
rect 10459 22185 10471 22188
rect 10413 22179 10471 22185
rect 13998 22176 14004 22188
rect 14056 22216 14062 22228
rect 15105 22219 15163 22225
rect 14056 22188 15056 22216
rect 14056 22176 14062 22188
rect 5077 22151 5135 22157
rect 5077 22117 5089 22151
rect 5123 22148 5135 22151
rect 8757 22151 8815 22157
rect 5123 22120 5856 22148
rect 5123 22117 5135 22120
rect 5077 22111 5135 22117
rect 5261 22083 5319 22089
rect 5261 22049 5273 22083
rect 5307 22080 5319 22083
rect 5442 22080 5448 22092
rect 5307 22052 5448 22080
rect 5307 22049 5319 22052
rect 5261 22043 5319 22049
rect 5442 22040 5448 22052
rect 5500 22088 5506 22092
rect 5500 22080 5580 22088
rect 5500 22060 5672 22080
rect 5500 22040 5506 22060
rect 5552 22052 5672 22060
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 992 21984 1409 22012
rect 992 21972 998 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 1397 21975 1455 21981
rect 2700 21984 3985 22012
rect 2700 21888 2728 21984
rect 3973 21981 3985 21984
rect 4019 22012 4031 22015
rect 4062 22012 4068 22024
rect 4019 21984 4068 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 4062 21972 4068 21984
rect 4120 22012 4126 22024
rect 4249 22015 4307 22021
rect 4249 22012 4261 22015
rect 4120 21984 4261 22012
rect 4120 21972 4126 21984
rect 4249 21981 4261 21984
rect 4295 21981 4307 22015
rect 4985 22015 5043 22021
rect 4985 22012 4997 22015
rect 4249 21975 4307 21981
rect 4632 21984 4997 22012
rect 4632 21888 4660 21984
rect 4985 21981 4997 21984
rect 5031 21981 5043 22015
rect 4985 21975 5043 21981
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 5644 22021 5672 22052
rect 5537 22015 5595 22021
rect 5537 22012 5549 22015
rect 5460 21984 5549 22012
rect 1578 21836 1584 21888
rect 1636 21836 1642 21888
rect 2682 21836 2688 21888
rect 2740 21836 2746 21888
rect 4614 21836 4620 21888
rect 4672 21836 4678 21888
rect 5166 21836 5172 21888
rect 5224 21876 5230 21888
rect 5460 21876 5488 21984
rect 5537 21981 5549 21984
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 21981 5687 22015
rect 5629 21975 5687 21981
rect 5718 21972 5724 22024
rect 5776 22012 5782 22024
rect 5828 22021 5856 22120
rect 8757 22117 8769 22151
rect 8803 22148 8815 22151
rect 10781 22151 10839 22157
rect 8803 22120 9904 22148
rect 8803 22117 8815 22120
rect 8757 22111 8815 22117
rect 9766 22080 9772 22092
rect 9508 22052 9772 22080
rect 5813 22015 5871 22021
rect 5813 22012 5825 22015
rect 5776 21984 5825 22012
rect 5776 21972 5782 21984
rect 5813 21981 5825 21984
rect 5859 21981 5871 22015
rect 5813 21975 5871 21981
rect 5902 21972 5908 22024
rect 5960 21972 5966 22024
rect 7745 22015 7803 22021
rect 7745 22012 7757 22015
rect 7668 21984 7757 22012
rect 7668 21888 7696 21984
rect 7745 21981 7757 21984
rect 7791 22012 7803 22015
rect 8018 22012 8024 22024
rect 7791 21984 8024 22012
rect 7791 21981 7803 21984
rect 7745 21975 7803 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9401 22015 9459 22021
rect 9171 21984 9352 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9324 21956 9352 21984
rect 9401 21981 9413 22015
rect 9447 22012 9459 22015
rect 9508 22012 9536 22052
rect 9766 22040 9772 22052
rect 9824 22040 9830 22092
rect 9447 21984 9536 22012
rect 9447 21981 9459 21984
rect 9401 21975 9459 21981
rect 9674 21972 9680 22024
rect 9732 21972 9738 22024
rect 9306 21904 9312 21956
rect 9364 21904 9370 21956
rect 6181 21879 6239 21885
rect 6181 21876 6193 21879
rect 5224 21848 6193 21876
rect 5224 21836 5230 21848
rect 6181 21845 6193 21848
rect 6227 21845 6239 21879
rect 6181 21839 6239 21845
rect 7650 21836 7656 21888
rect 7708 21836 7714 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 7837 21879 7895 21885
rect 7837 21876 7849 21879
rect 7800 21848 7849 21876
rect 7800 21836 7806 21848
rect 7837 21845 7849 21848
rect 7883 21845 7895 21879
rect 7837 21839 7895 21845
rect 8018 21836 8024 21888
rect 8076 21876 8082 21888
rect 8113 21879 8171 21885
rect 8113 21876 8125 21879
rect 8076 21848 8125 21876
rect 8076 21836 8082 21848
rect 8113 21845 8125 21848
rect 8159 21845 8171 21879
rect 8113 21839 8171 21845
rect 9217 21879 9275 21885
rect 9217 21845 9229 21879
rect 9263 21876 9275 21879
rect 9490 21876 9496 21888
rect 9263 21848 9496 21876
rect 9263 21845 9275 21848
rect 9217 21839 9275 21845
rect 9490 21836 9496 21848
rect 9548 21836 9554 21888
rect 9582 21836 9588 21888
rect 9640 21836 9646 21888
rect 9784 21876 9812 22040
rect 9876 22021 9904 22120
rect 10781 22117 10793 22151
rect 10827 22148 10839 22151
rect 10962 22148 10968 22160
rect 10827 22120 10968 22148
rect 10827 22117 10839 22120
rect 10781 22111 10839 22117
rect 10962 22108 10968 22120
rect 11020 22108 11026 22160
rect 13081 22151 13139 22157
rect 13081 22117 13093 22151
rect 13127 22148 13139 22151
rect 14642 22148 14648 22160
rect 13127 22120 14648 22148
rect 13127 22117 13139 22120
rect 13081 22111 13139 22117
rect 14642 22108 14648 22120
rect 14700 22108 14706 22160
rect 10137 22083 10195 22089
rect 10137 22049 10149 22083
rect 10183 22080 10195 22083
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 10183 22052 10701 22080
rect 10183 22049 10195 22052
rect 10137 22043 10195 22049
rect 10689 22049 10701 22052
rect 10735 22080 10747 22083
rect 10735 22052 11560 22080
rect 10735 22049 10747 22052
rect 10689 22043 10747 22049
rect 9861 22015 9919 22021
rect 9861 21981 9873 22015
rect 9907 21981 9919 22015
rect 9861 21975 9919 21981
rect 9876 21944 9904 21975
rect 10226 21972 10232 22024
rect 10284 21972 10290 22024
rect 10870 21972 10876 22024
rect 10928 21972 10934 22024
rect 11532 22021 11560 22052
rect 11790 22040 11796 22092
rect 11848 22040 11854 22092
rect 12526 22080 12532 22092
rect 11992 22052 12532 22080
rect 11149 22015 11207 22021
rect 11149 21981 11161 22015
rect 11195 21981 11207 22015
rect 11149 21975 11207 21981
rect 11517 22015 11575 22021
rect 11517 21981 11529 22015
rect 11563 22012 11575 22015
rect 11808 22012 11836 22040
rect 11563 21984 11836 22012
rect 11563 21981 11575 21984
rect 11517 21975 11575 21981
rect 11164 21944 11192 21975
rect 11882 21972 11888 22024
rect 11940 21972 11946 22024
rect 11992 22021 12020 22052
rect 12526 22040 12532 22052
rect 12584 22080 12590 22092
rect 13262 22080 13268 22092
rect 12584 22052 13268 22080
rect 12584 22040 12590 22052
rect 13262 22040 13268 22052
rect 13320 22040 13326 22092
rect 15028 22080 15056 22188
rect 15105 22185 15117 22219
rect 15151 22216 15163 22219
rect 15286 22216 15292 22228
rect 15151 22188 15292 22216
rect 15151 22185 15163 22188
rect 15105 22179 15163 22185
rect 15286 22176 15292 22188
rect 15344 22176 15350 22228
rect 20898 22176 20904 22228
rect 20956 22216 20962 22228
rect 23017 22219 23075 22225
rect 23017 22216 23029 22219
rect 20956 22188 23029 22216
rect 20956 22176 20962 22188
rect 23017 22185 23029 22188
rect 23063 22216 23075 22219
rect 23382 22216 23388 22228
rect 23063 22188 23388 22216
rect 23063 22185 23075 22188
rect 23017 22179 23075 22185
rect 23382 22176 23388 22188
rect 23440 22176 23446 22228
rect 30374 22176 30380 22228
rect 30432 22176 30438 22228
rect 30926 22176 30932 22228
rect 30984 22176 30990 22228
rect 34146 22176 34152 22228
rect 34204 22216 34210 22228
rect 34241 22219 34299 22225
rect 34241 22216 34253 22219
rect 34204 22188 34253 22216
rect 34204 22176 34210 22188
rect 34241 22185 34253 22188
rect 34287 22185 34299 22219
rect 34241 22179 34299 22185
rect 18046 22108 18052 22160
rect 18104 22108 18110 22160
rect 26234 22148 26240 22160
rect 20548 22120 26240 22148
rect 13464 22052 14596 22080
rect 15028 22052 15424 22080
rect 11977 22015 12035 22021
rect 11977 21981 11989 22015
rect 12023 21981 12035 22015
rect 11977 21975 12035 21981
rect 12437 22015 12495 22021
rect 12437 21981 12449 22015
rect 12483 21981 12495 22015
rect 12437 21975 12495 21981
rect 11992 21944 12020 21975
rect 12452 21944 12480 21975
rect 12710 21972 12716 22024
rect 12768 21972 12774 22024
rect 12802 21972 12808 22024
rect 12860 21972 12866 22024
rect 9876 21916 11100 21944
rect 11164 21916 12020 21944
rect 12406 21916 12480 21944
rect 12728 21944 12756 21972
rect 13464 21953 13492 22052
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13553 21984 14105 22012
rect 13449 21947 13507 21953
rect 13449 21944 13461 21947
rect 12728 21916 13461 21944
rect 11072 21888 11100 21916
rect 10134 21876 10140 21888
rect 9784 21848 10140 21876
rect 10134 21836 10140 21848
rect 10192 21836 10198 21888
rect 11054 21836 11060 21888
rect 11112 21876 11118 21888
rect 11698 21876 11704 21888
rect 11112 21848 11704 21876
rect 11112 21836 11118 21848
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 11790 21836 11796 21888
rect 11848 21876 11854 21888
rect 12406 21876 12434 21916
rect 13449 21913 13461 21916
rect 13495 21913 13507 21947
rect 13449 21907 13507 21913
rect 11848 21848 12434 21876
rect 11848 21836 11854 21848
rect 12618 21836 12624 21888
rect 12676 21876 12682 21888
rect 13553 21876 13581 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14185 22015 14243 22021
rect 14185 21981 14197 22015
rect 14231 22012 14243 22015
rect 14274 22012 14280 22024
rect 14231 21984 14280 22012
rect 14231 21981 14243 21984
rect 14185 21975 14243 21981
rect 14274 21972 14280 21984
rect 14332 21972 14338 22024
rect 14568 22021 14596 22052
rect 14553 22015 14611 22021
rect 14553 21981 14565 22015
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 15010 21972 15016 22024
rect 15068 22012 15074 22024
rect 15396 22021 15424 22052
rect 17586 22040 17592 22092
rect 17644 22040 17650 22092
rect 19334 22040 19340 22092
rect 19392 22080 19398 22092
rect 20548 22089 20576 22120
rect 26234 22108 26240 22120
rect 26292 22108 26298 22160
rect 26326 22108 26332 22160
rect 26384 22108 26390 22160
rect 26804 22120 27844 22148
rect 20533 22083 20591 22089
rect 19392 22052 19932 22080
rect 19392 22040 19398 22052
rect 15105 22015 15163 22021
rect 15105 22012 15117 22015
rect 15068 21984 15117 22012
rect 15068 21972 15074 21984
rect 15105 21981 15117 21984
rect 15151 21981 15163 22015
rect 15105 21975 15163 21981
rect 15381 22015 15439 22021
rect 15381 21981 15393 22015
rect 15427 22012 15439 22015
rect 15654 22012 15660 22024
rect 15427 21984 15660 22012
rect 15427 21981 15439 21984
rect 15381 21975 15439 21981
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 17678 21972 17684 22024
rect 17736 21972 17742 22024
rect 19518 21972 19524 22024
rect 19576 21972 19582 22024
rect 19904 22021 19932 22052
rect 20533 22049 20545 22083
rect 20579 22049 20591 22083
rect 20533 22043 20591 22049
rect 21726 22040 21732 22092
rect 21784 22040 21790 22092
rect 22465 22083 22523 22089
rect 22465 22049 22477 22083
rect 22511 22080 22523 22083
rect 22554 22080 22560 22092
rect 22511 22052 22560 22080
rect 22511 22049 22523 22052
rect 22465 22043 22523 22049
rect 22554 22040 22560 22052
rect 22612 22040 22618 22092
rect 25961 22083 26019 22089
rect 25961 22049 25973 22083
rect 26007 22080 26019 22083
rect 26050 22080 26056 22092
rect 26007 22052 26056 22080
rect 26007 22049 26019 22052
rect 25961 22043 26019 22049
rect 26050 22040 26056 22052
rect 26108 22040 26114 22092
rect 26602 22080 26608 22092
rect 26436 22052 26608 22080
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 22012 19947 22015
rect 20070 22012 20076 22024
rect 19935 21984 20076 22012
rect 19935 21981 19947 21984
rect 19889 21975 19947 21981
rect 20070 21972 20076 21984
rect 20128 21972 20134 22024
rect 26436 22021 26464 22052
rect 26602 22040 26608 22052
rect 26660 22040 26666 22092
rect 21177 22015 21235 22021
rect 21177 21981 21189 22015
rect 21223 22012 21235 22015
rect 21269 22015 21327 22021
rect 21269 22012 21281 22015
rect 21223 21984 21281 22012
rect 21223 21981 21235 21984
rect 21177 21975 21235 21981
rect 21269 21981 21281 21984
rect 21315 22012 21327 22015
rect 26421 22015 26479 22021
rect 21315 21984 22508 22012
rect 21315 21981 21327 21984
rect 21269 21975 21327 21981
rect 22480 21956 22508 21984
rect 26421 21981 26433 22015
rect 26467 21981 26479 22015
rect 26697 22015 26755 22021
rect 26697 22012 26709 22015
rect 26421 21975 26479 21981
rect 26528 21984 26709 22012
rect 13814 21904 13820 21956
rect 13872 21944 13878 21956
rect 13909 21947 13967 21953
rect 13909 21944 13921 21947
rect 13872 21916 13921 21944
rect 13872 21904 13878 21916
rect 13909 21913 13921 21916
rect 13955 21944 13967 21947
rect 14366 21944 14372 21956
rect 13955 21916 14372 21944
rect 13955 21913 13967 21916
rect 13909 21907 13967 21913
rect 14366 21904 14372 21916
rect 14424 21904 14430 21956
rect 14461 21947 14519 21953
rect 14461 21913 14473 21947
rect 14507 21944 14519 21947
rect 21361 21947 21419 21953
rect 21361 21944 21373 21947
rect 14507 21916 21373 21944
rect 14507 21913 14519 21916
rect 14461 21907 14519 21913
rect 21361 21913 21373 21916
rect 21407 21944 21419 21947
rect 22186 21944 22192 21956
rect 21407 21916 22192 21944
rect 21407 21913 21419 21916
rect 21361 21907 21419 21913
rect 22186 21904 22192 21916
rect 22244 21904 22250 21956
rect 22462 21904 22468 21956
rect 22520 21904 22526 21956
rect 26528 21888 26556 21984
rect 26697 21981 26709 21984
rect 26743 22012 26755 22015
rect 26804 22012 26832 22120
rect 27246 22040 27252 22092
rect 27304 22080 27310 22092
rect 27525 22083 27583 22089
rect 27525 22080 27537 22083
rect 27304 22052 27537 22080
rect 27304 22040 27310 22052
rect 27525 22049 27537 22052
rect 27571 22049 27583 22083
rect 27525 22043 27583 22049
rect 27816 22024 27844 22120
rect 27890 22108 27896 22160
rect 27948 22108 27954 22160
rect 27908 22080 27936 22108
rect 28353 22083 28411 22089
rect 28353 22080 28365 22083
rect 27908 22052 28120 22080
rect 26743 21984 26832 22012
rect 26743 21981 26755 21984
rect 26697 21975 26755 21981
rect 26878 21972 26884 22024
rect 26936 21972 26942 22024
rect 27338 21972 27344 22024
rect 27396 21972 27402 22024
rect 27706 21972 27712 22024
rect 27764 21972 27770 22024
rect 27798 21972 27804 22024
rect 27856 21972 27862 22024
rect 28092 22021 28120 22052
rect 28276 22052 28365 22080
rect 27893 22015 27951 22021
rect 27893 21981 27905 22015
rect 27939 21981 27951 22015
rect 27893 21975 27951 21981
rect 28077 22015 28135 22021
rect 28077 21981 28089 22015
rect 28123 21981 28135 22015
rect 28077 21975 28135 21981
rect 28169 22015 28227 22021
rect 28169 21981 28181 22015
rect 28215 21981 28227 22015
rect 28169 21975 28227 21981
rect 26786 21904 26792 21956
rect 26844 21944 26850 21956
rect 27019 21947 27077 21953
rect 27019 21944 27031 21947
rect 26844 21916 27031 21944
rect 26844 21904 26850 21916
rect 27019 21913 27031 21916
rect 27065 21913 27077 21947
rect 27019 21907 27077 21913
rect 27154 21904 27160 21956
rect 27212 21904 27218 21956
rect 27249 21947 27307 21953
rect 27249 21913 27261 21947
rect 27295 21944 27307 21947
rect 27617 21947 27675 21953
rect 27617 21944 27629 21947
rect 27295 21916 27629 21944
rect 27295 21913 27307 21916
rect 27249 21907 27307 21913
rect 27617 21913 27629 21916
rect 27663 21913 27675 21947
rect 27724 21944 27752 21972
rect 27908 21944 27936 21975
rect 27724 21916 27936 21944
rect 27617 21907 27675 21913
rect 27982 21904 27988 21956
rect 28040 21944 28046 21956
rect 28184 21944 28212 21975
rect 28040 21916 28212 21944
rect 28040 21904 28046 21916
rect 12676 21848 13581 21876
rect 12676 21836 12682 21848
rect 14090 21836 14096 21888
rect 14148 21876 14154 21888
rect 14737 21879 14795 21885
rect 14737 21876 14749 21879
rect 14148 21848 14749 21876
rect 14148 21836 14154 21848
rect 14737 21845 14749 21848
rect 14783 21845 14795 21879
rect 14737 21839 14795 21845
rect 15286 21836 15292 21888
rect 15344 21836 15350 21888
rect 26510 21836 26516 21888
rect 26568 21836 26574 21888
rect 26602 21836 26608 21888
rect 26660 21836 26666 21888
rect 26878 21836 26884 21888
rect 26936 21876 26942 21888
rect 27522 21876 27528 21888
rect 26936 21848 27528 21876
rect 26936 21836 26942 21848
rect 27522 21836 27528 21848
rect 27580 21876 27586 21888
rect 28276 21876 28304 22052
rect 28353 22049 28365 22052
rect 28399 22049 28411 22083
rect 28353 22043 28411 22049
rect 28813 22083 28871 22089
rect 28813 22049 28825 22083
rect 28859 22049 28871 22083
rect 28813 22043 28871 22049
rect 28442 21972 28448 22024
rect 28500 21972 28506 22024
rect 28828 21888 28856 22043
rect 31754 22040 31760 22092
rect 31812 22080 31818 22092
rect 31849 22083 31907 22089
rect 31849 22080 31861 22083
rect 31812 22052 31861 22080
rect 31812 22040 31818 22052
rect 31849 22049 31861 22052
rect 31895 22049 31907 22083
rect 31849 22043 31907 22049
rect 30101 22015 30159 22021
rect 30101 21981 30113 22015
rect 30147 22012 30159 22015
rect 30193 22015 30251 22021
rect 30193 22012 30205 22015
rect 30147 21984 30205 22012
rect 30147 21981 30159 21984
rect 30101 21975 30159 21981
rect 30193 21981 30205 21984
rect 30239 21981 30251 22015
rect 30837 22015 30895 22021
rect 30837 22012 30849 22015
rect 30193 21975 30251 21981
rect 30668 21984 30849 22012
rect 29086 21904 29092 21956
rect 29144 21944 29150 21956
rect 29733 21947 29791 21953
rect 29733 21944 29745 21947
rect 29144 21916 29745 21944
rect 29144 21904 29150 21916
rect 29733 21913 29745 21916
rect 29779 21913 29791 21947
rect 29733 21907 29791 21913
rect 29914 21904 29920 21956
rect 29972 21904 29978 21956
rect 30668 21888 30696 21984
rect 30837 21981 30849 21984
rect 30883 21981 30895 22015
rect 30837 21975 30895 21981
rect 32030 21972 32036 22024
rect 32088 21972 32094 22024
rect 34054 21972 34060 22024
rect 34112 22012 34118 22024
rect 34149 22015 34207 22021
rect 34149 22012 34161 22015
rect 34112 21984 34161 22012
rect 34112 21972 34118 21984
rect 34149 21981 34161 21984
rect 34195 21981 34207 22015
rect 34149 21975 34207 21981
rect 32217 21947 32275 21953
rect 32217 21913 32229 21947
rect 32263 21944 32275 21947
rect 32490 21944 32496 21956
rect 32263 21916 32496 21944
rect 32263 21913 32275 21916
rect 32217 21907 32275 21913
rect 32490 21904 32496 21916
rect 32548 21904 32554 21956
rect 27580 21848 28304 21876
rect 27580 21836 27586 21848
rect 28810 21836 28816 21888
rect 28868 21836 28874 21888
rect 30650 21836 30656 21888
rect 30708 21836 30714 21888
rect 32674 21836 32680 21888
rect 32732 21876 32738 21888
rect 32953 21879 33011 21885
rect 32953 21876 32965 21879
rect 32732 21848 32965 21876
rect 32732 21836 32738 21848
rect 32953 21845 32965 21848
rect 32999 21845 33011 21879
rect 32953 21839 33011 21845
rect 34057 21879 34115 21885
rect 34057 21845 34069 21879
rect 34103 21876 34115 21879
rect 34164 21876 34192 21975
rect 34422 21876 34428 21888
rect 34103 21848 34428 21876
rect 34103 21845 34115 21848
rect 34057 21839 34115 21845
rect 34422 21836 34428 21848
rect 34480 21836 34486 21888
rect 1104 21786 35236 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 35236 21786
rect 1104 21712 35236 21734
rect 1578 21632 1584 21684
rect 1636 21632 1642 21684
rect 4614 21632 4620 21684
rect 4672 21672 4678 21684
rect 5902 21672 5908 21684
rect 4672 21644 5908 21672
rect 4672 21632 4678 21644
rect 1596 21604 1624 21632
rect 3145 21607 3203 21613
rect 3145 21604 3157 21607
rect 1596 21576 3157 21604
rect 3145 21573 3157 21576
rect 3191 21573 3203 21607
rect 4801 21607 4859 21613
rect 4801 21604 4813 21607
rect 4370 21576 4813 21604
rect 3145 21567 3203 21573
rect 4801 21573 4813 21576
rect 4847 21573 4859 21607
rect 4801 21567 4859 21573
rect 4982 21564 4988 21616
rect 5040 21564 5046 21616
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 2682 21536 2688 21548
rect 2179 21508 2688 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2682 21496 2688 21508
rect 2740 21496 2746 21548
rect 4890 21496 4896 21548
rect 4948 21496 4954 21548
rect 5166 21496 5172 21548
rect 5224 21496 5230 21548
rect 5258 21496 5264 21548
rect 5316 21496 5322 21548
rect 5350 21496 5356 21548
rect 5408 21496 5414 21548
rect 5460 21536 5488 21644
rect 5902 21632 5908 21644
rect 5960 21632 5966 21684
rect 9306 21632 9312 21684
rect 9364 21672 9370 21684
rect 10502 21672 10508 21684
rect 9364 21644 10508 21672
rect 9364 21632 9370 21644
rect 10502 21632 10508 21644
rect 10560 21632 10566 21684
rect 10965 21675 11023 21681
rect 10965 21641 10977 21675
rect 11011 21672 11023 21675
rect 11790 21672 11796 21684
rect 11011 21644 11796 21672
rect 11011 21641 11023 21644
rect 10965 21635 11023 21641
rect 11790 21632 11796 21644
rect 11848 21632 11854 21684
rect 11882 21632 11888 21684
rect 11940 21632 11946 21684
rect 12066 21632 12072 21684
rect 12124 21632 12130 21684
rect 12158 21632 12164 21684
rect 12216 21632 12222 21684
rect 12710 21632 12716 21684
rect 12768 21672 12774 21684
rect 13541 21675 13599 21681
rect 13541 21672 13553 21675
rect 12768 21644 13553 21672
rect 12768 21632 12774 21644
rect 13541 21641 13553 21644
rect 13587 21672 13599 21675
rect 13814 21672 13820 21684
rect 13587 21644 13820 21672
rect 13587 21641 13599 21644
rect 13541 21635 13599 21641
rect 13814 21632 13820 21644
rect 13872 21672 13878 21684
rect 14458 21672 14464 21684
rect 13872 21644 14464 21672
rect 13872 21632 13878 21644
rect 14458 21632 14464 21644
rect 14516 21632 14522 21684
rect 14642 21632 14648 21684
rect 14700 21632 14706 21684
rect 17586 21632 17592 21684
rect 17644 21632 17650 21684
rect 19242 21632 19248 21684
rect 19300 21672 19306 21684
rect 21726 21672 21732 21684
rect 19300 21644 21732 21672
rect 19300 21632 19306 21644
rect 21726 21632 21732 21644
rect 21784 21672 21790 21684
rect 21784 21644 22094 21672
rect 21784 21632 21790 21644
rect 5810 21564 5816 21616
rect 5868 21604 5874 21616
rect 5868 21576 6592 21604
rect 5868 21564 5874 21576
rect 5537 21539 5595 21545
rect 5537 21536 5549 21539
rect 5460 21508 5549 21536
rect 5537 21505 5549 21508
rect 5583 21505 5595 21539
rect 5537 21499 5595 21505
rect 5718 21496 5724 21548
rect 5776 21536 5782 21548
rect 6564 21545 6592 21576
rect 8018 21564 8024 21616
rect 8076 21564 8082 21616
rect 5997 21539 6055 21545
rect 5997 21536 6009 21539
rect 5776 21508 6009 21536
rect 5776 21496 5782 21508
rect 5997 21505 6009 21508
rect 6043 21505 6055 21539
rect 5997 21499 6055 21505
rect 6181 21539 6239 21545
rect 6181 21505 6193 21539
rect 6227 21505 6239 21539
rect 6181 21499 6239 21505
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6549 21539 6607 21545
rect 6549 21505 6561 21539
rect 6595 21505 6607 21539
rect 6549 21499 6607 21505
rect 1394 21428 1400 21480
rect 1452 21468 1458 21480
rect 2590 21468 2596 21480
rect 1452 21440 2596 21468
rect 1452 21428 1458 21440
rect 2590 21428 2596 21440
rect 2648 21468 2654 21480
rect 2869 21471 2927 21477
rect 2869 21468 2881 21471
rect 2648 21440 2881 21468
rect 2648 21428 2654 21440
rect 2869 21437 2881 21440
rect 2915 21468 2927 21471
rect 3142 21468 3148 21480
rect 2915 21440 3148 21468
rect 2915 21437 2927 21440
rect 2869 21431 2927 21437
rect 3142 21428 3148 21440
rect 3200 21428 3206 21480
rect 4985 21471 5043 21477
rect 4985 21437 4997 21471
rect 5031 21437 5043 21471
rect 4985 21431 5043 21437
rect 5000 21344 5028 21431
rect 5074 21360 5080 21412
rect 5132 21400 5138 21412
rect 5368 21400 5396 21496
rect 5445 21471 5503 21477
rect 5445 21437 5457 21471
rect 5491 21468 5503 21471
rect 6089 21471 6147 21477
rect 6089 21468 6101 21471
rect 5491 21440 6101 21468
rect 5491 21437 5503 21440
rect 5445 21431 5503 21437
rect 6089 21437 6101 21440
rect 6135 21437 6147 21471
rect 6089 21431 6147 21437
rect 6196 21400 6224 21499
rect 6380 21412 6408 21499
rect 8846 21496 8852 21548
rect 8904 21496 8910 21548
rect 9953 21539 10011 21545
rect 9953 21536 9965 21539
rect 9416 21508 9965 21536
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 6822 21468 6828 21480
rect 6512 21440 6828 21468
rect 6512 21428 6518 21440
rect 6822 21428 6828 21440
rect 6880 21468 6886 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6880 21440 7021 21468
rect 6880 21428 6886 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7285 21471 7343 21477
rect 7285 21468 7297 21471
rect 7009 21431 7067 21437
rect 7116 21440 7297 21468
rect 5132 21372 6224 21400
rect 5132 21360 5138 21372
rect 6362 21360 6368 21412
rect 6420 21360 6426 21412
rect 6638 21360 6644 21412
rect 6696 21400 6702 21412
rect 7116 21400 7144 21440
rect 7285 21437 7297 21440
rect 7331 21437 7343 21471
rect 7285 21431 7343 21437
rect 8757 21471 8815 21477
rect 8757 21437 8769 21471
rect 8803 21468 8815 21471
rect 9416 21468 9444 21508
rect 9953 21505 9965 21508
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 10226 21496 10232 21548
rect 10284 21536 10290 21548
rect 10781 21539 10839 21545
rect 10781 21536 10793 21539
rect 10284 21508 10793 21536
rect 10284 21496 10290 21508
rect 10781 21505 10793 21508
rect 10827 21505 10839 21539
rect 10781 21499 10839 21505
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 8803 21440 9444 21468
rect 8803 21437 8815 21440
rect 8757 21431 8815 21437
rect 9490 21428 9496 21480
rect 9548 21428 9554 21480
rect 10137 21471 10195 21477
rect 10137 21437 10149 21471
rect 10183 21468 10195 21471
rect 10318 21468 10324 21480
rect 10183 21440 10324 21468
rect 10183 21437 10195 21440
rect 10137 21431 10195 21437
rect 10318 21428 10324 21440
rect 10376 21428 10382 21480
rect 6696 21372 7144 21400
rect 6696 21360 6702 21372
rect 10980 21344 11008 21499
rect 11054 21496 11060 21548
rect 11112 21536 11118 21548
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 11112 21508 11529 21536
rect 11112 21496 11118 21508
rect 11517 21505 11529 21508
rect 11563 21505 11575 21539
rect 11517 21499 11575 21505
rect 11701 21539 11759 21545
rect 11701 21505 11713 21539
rect 11747 21536 11759 21539
rect 11808 21536 11836 21632
rect 11900 21545 11928 21632
rect 12084 21604 12112 21632
rect 13173 21607 13231 21613
rect 13173 21604 13185 21607
rect 12084 21576 13185 21604
rect 13173 21573 13185 21576
rect 13219 21604 13231 21607
rect 13630 21604 13636 21616
rect 13219 21576 13636 21604
rect 13219 21573 13231 21576
rect 13173 21567 13231 21573
rect 13630 21564 13636 21576
rect 13688 21564 13694 21616
rect 13998 21564 14004 21616
rect 14056 21604 14062 21616
rect 14553 21607 14611 21613
rect 14553 21604 14565 21607
rect 14056 21576 14565 21604
rect 14056 21564 14062 21576
rect 14553 21573 14565 21576
rect 14599 21573 14611 21607
rect 14553 21567 14611 21573
rect 15488 21576 17172 21604
rect 11747 21508 11836 21536
rect 11885 21539 11943 21545
rect 11747 21505 11759 21508
rect 11701 21499 11759 21505
rect 11885 21505 11897 21539
rect 11931 21505 11943 21539
rect 11885 21499 11943 21505
rect 11532 21400 11560 21499
rect 11974 21496 11980 21548
rect 12032 21496 12038 21548
rect 13078 21496 13084 21548
rect 13136 21536 13142 21548
rect 14829 21539 14887 21545
rect 14829 21536 14841 21539
rect 13136 21508 14841 21536
rect 13136 21496 13142 21508
rect 14829 21505 14841 21508
rect 14875 21536 14887 21539
rect 15010 21536 15016 21548
rect 14875 21508 15016 21536
rect 14875 21505 14887 21508
rect 14829 21499 14887 21505
rect 15010 21496 15016 21508
rect 15068 21536 15074 21548
rect 15197 21539 15255 21545
rect 15197 21536 15209 21539
rect 15068 21508 15209 21536
rect 15068 21496 15074 21508
rect 15197 21505 15209 21508
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 15286 21496 15292 21548
rect 15344 21536 15350 21548
rect 15381 21539 15439 21545
rect 15381 21536 15393 21539
rect 15344 21508 15393 21536
rect 15344 21496 15350 21508
rect 15381 21505 15393 21508
rect 15427 21505 15439 21539
rect 15381 21499 15439 21505
rect 11793 21471 11851 21477
rect 11793 21437 11805 21471
rect 11839 21468 11851 21471
rect 12526 21468 12532 21480
rect 11839 21440 12532 21468
rect 11839 21437 11851 21440
rect 11793 21431 11851 21437
rect 12526 21428 12532 21440
rect 12584 21428 12590 21480
rect 14642 21428 14648 21480
rect 14700 21468 14706 21480
rect 15396 21468 15424 21499
rect 14700 21440 15424 21468
rect 14700 21428 14706 21440
rect 12802 21400 12808 21412
rect 11532 21372 12808 21400
rect 12802 21360 12808 21372
rect 12860 21360 12866 21412
rect 2222 21292 2228 21344
rect 2280 21292 2286 21344
rect 2682 21292 2688 21344
rect 2740 21332 2746 21344
rect 2866 21332 2872 21344
rect 2740 21304 2872 21332
rect 2740 21292 2746 21304
rect 2866 21292 2872 21304
rect 2924 21292 2930 21344
rect 4982 21292 4988 21344
rect 5040 21292 5046 21344
rect 5813 21335 5871 21341
rect 5813 21301 5825 21335
rect 5859 21332 5871 21335
rect 6546 21332 6552 21344
rect 5859 21304 6552 21332
rect 5859 21301 5871 21304
rect 5813 21295 5871 21301
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 6730 21292 6736 21344
rect 6788 21292 6794 21344
rect 10962 21292 10968 21344
rect 11020 21332 11026 21344
rect 11974 21332 11980 21344
rect 11020 21304 11980 21332
rect 11020 21292 11026 21304
rect 11974 21292 11980 21304
rect 12032 21292 12038 21344
rect 12621 21335 12679 21341
rect 12621 21301 12633 21335
rect 12667 21332 12679 21335
rect 12894 21332 12900 21344
rect 12667 21304 12900 21332
rect 12667 21301 12679 21304
rect 12621 21295 12679 21301
rect 12894 21292 12900 21304
rect 12952 21292 12958 21344
rect 15013 21335 15071 21341
rect 15013 21301 15025 21335
rect 15059 21332 15071 21335
rect 15488 21332 15516 21576
rect 15654 21496 15660 21548
rect 15712 21496 15718 21548
rect 16666 21496 16672 21548
rect 16724 21536 16730 21548
rect 16853 21539 16911 21545
rect 16853 21536 16865 21539
rect 16724 21508 16865 21536
rect 16724 21496 16730 21508
rect 16853 21505 16865 21508
rect 16899 21505 16911 21539
rect 16853 21499 16911 21505
rect 15565 21471 15623 21477
rect 15565 21437 15577 21471
rect 15611 21468 15623 21471
rect 15611 21440 16896 21468
rect 15611 21437 15623 21440
rect 15565 21431 15623 21437
rect 15059 21304 15516 21332
rect 16868 21332 16896 21440
rect 16942 21428 16948 21480
rect 17000 21428 17006 21480
rect 17144 21400 17172 21576
rect 17221 21471 17279 21477
rect 17221 21437 17233 21471
rect 17267 21468 17279 21471
rect 17604 21468 17632 21632
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21536 19395 21539
rect 20622 21536 20628 21548
rect 19383 21508 20628 21536
rect 19383 21505 19395 21508
rect 19337 21499 19395 21505
rect 17267 21440 17632 21468
rect 17267 21437 17279 21440
rect 17221 21431 17279 21437
rect 19352 21400 19380 21499
rect 20622 21496 20628 21508
rect 20680 21496 20686 21548
rect 19426 21428 19432 21480
rect 19484 21428 19490 21480
rect 22066 21468 22094 21644
rect 22554 21632 22560 21684
rect 22612 21632 22618 21684
rect 23109 21675 23167 21681
rect 23109 21641 23121 21675
rect 23155 21672 23167 21675
rect 23566 21672 23572 21684
rect 23155 21644 23572 21672
rect 23155 21641 23167 21644
rect 23109 21635 23167 21641
rect 23566 21632 23572 21644
rect 23624 21632 23630 21684
rect 26786 21632 26792 21684
rect 26844 21632 26850 21684
rect 27154 21632 27160 21684
rect 27212 21632 27218 21684
rect 27706 21672 27712 21684
rect 27264 21644 27712 21672
rect 22572 21604 22600 21632
rect 22830 21604 22836 21616
rect 22572 21576 22836 21604
rect 22830 21564 22836 21576
rect 22888 21604 22894 21616
rect 23385 21607 23443 21613
rect 23385 21604 23397 21607
rect 22888 21576 23397 21604
rect 22888 21564 22894 21576
rect 23124 21545 23152 21576
rect 23385 21573 23397 21576
rect 23431 21573 23443 21607
rect 26602 21604 26608 21616
rect 23385 21567 23443 21573
rect 26436 21576 26608 21604
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 23109 21539 23167 21545
rect 23109 21505 23121 21539
rect 23155 21536 23167 21539
rect 23155 21508 23189 21536
rect 23155 21505 23167 21508
rect 23109 21499 23167 21505
rect 22649 21471 22707 21477
rect 22649 21468 22661 21471
rect 22066 21440 22661 21468
rect 22649 21437 22661 21440
rect 22695 21468 22707 21471
rect 22940 21468 22968 21499
rect 22695 21440 23336 21468
rect 22695 21437 22707 21440
rect 22649 21431 22707 21437
rect 17144 21372 19380 21400
rect 19702 21360 19708 21412
rect 19760 21360 19766 21412
rect 23308 21344 23336 21440
rect 26326 21428 26332 21480
rect 26384 21428 26390 21480
rect 26436 21477 26464 21576
rect 26602 21564 26608 21576
rect 26660 21604 26666 21616
rect 27264 21604 27292 21644
rect 27706 21632 27712 21644
rect 27764 21672 27770 21684
rect 27801 21675 27859 21681
rect 27801 21672 27813 21675
rect 27764 21644 27813 21672
rect 27764 21632 27770 21644
rect 27801 21641 27813 21644
rect 27847 21641 27859 21675
rect 27801 21635 27859 21641
rect 27890 21632 27896 21684
rect 27948 21672 27954 21684
rect 27985 21675 28043 21681
rect 27985 21672 27997 21675
rect 27948 21644 27997 21672
rect 27948 21632 27954 21644
rect 27985 21641 27997 21644
rect 28031 21641 28043 21675
rect 27985 21635 28043 21641
rect 29086 21632 29092 21684
rect 29144 21632 29150 21684
rect 29358 21675 29416 21681
rect 29358 21641 29370 21675
rect 29404 21672 29416 21675
rect 29914 21672 29920 21684
rect 29404 21644 29920 21672
rect 29404 21641 29416 21644
rect 29358 21635 29416 21641
rect 29914 21632 29920 21644
rect 29972 21632 29978 21684
rect 28353 21607 28411 21613
rect 28353 21604 28365 21607
rect 26660 21576 27292 21604
rect 27540 21576 28365 21604
rect 26660 21564 26666 21576
rect 27540 21548 27568 21576
rect 28353 21573 28365 21576
rect 28399 21573 28411 21607
rect 28353 21567 28411 21573
rect 28718 21564 28724 21616
rect 28776 21564 28782 21616
rect 28810 21564 28816 21616
rect 28868 21604 28874 21616
rect 28937 21607 28995 21613
rect 28937 21604 28949 21607
rect 28868 21576 28949 21604
rect 28868 21564 28874 21576
rect 28937 21573 28949 21576
rect 28983 21604 28995 21607
rect 29457 21607 29515 21613
rect 29457 21604 29469 21607
rect 28983 21576 29469 21604
rect 28983 21573 28995 21576
rect 28937 21567 28995 21573
rect 29457 21573 29469 21576
rect 29503 21573 29515 21607
rect 29457 21567 29515 21573
rect 26510 21496 26516 21548
rect 26568 21496 26574 21548
rect 26786 21496 26792 21548
rect 26844 21496 26850 21548
rect 27522 21496 27528 21548
rect 27580 21496 27586 21548
rect 27798 21496 27804 21548
rect 27856 21536 27862 21548
rect 27893 21539 27951 21545
rect 27893 21536 27905 21539
rect 27856 21508 27905 21536
rect 27856 21496 27862 21508
rect 27893 21505 27905 21508
rect 27939 21505 27951 21539
rect 27893 21499 27951 21505
rect 28166 21496 28172 21548
rect 28224 21496 28230 21548
rect 29181 21539 29239 21545
rect 29181 21536 29193 21539
rect 28920 21508 29193 21536
rect 26421 21471 26479 21477
rect 26421 21437 26433 21471
rect 26467 21437 26479 21471
rect 26421 21431 26479 21437
rect 26605 21471 26663 21477
rect 26605 21437 26617 21471
rect 26651 21437 26663 21471
rect 26605 21431 26663 21437
rect 26620 21400 26648 21431
rect 26694 21400 26700 21412
rect 26620 21372 26700 21400
rect 26694 21360 26700 21372
rect 26752 21360 26758 21412
rect 26804 21400 26832 21496
rect 28920 21400 28948 21508
rect 29181 21505 29193 21508
rect 29227 21505 29239 21539
rect 29181 21499 29239 21505
rect 29273 21539 29331 21545
rect 29273 21505 29285 21539
rect 29319 21505 29331 21539
rect 29273 21499 29331 21505
rect 28994 21428 29000 21480
rect 29052 21468 29058 21480
rect 29288 21468 29316 21499
rect 29052 21440 29316 21468
rect 29052 21428 29058 21440
rect 26804 21372 28948 21400
rect 20714 21332 20720 21344
rect 16868 21304 20720 21332
rect 15059 21301 15071 21304
rect 15013 21295 15071 21301
rect 20714 21292 20720 21304
rect 20772 21292 20778 21344
rect 21818 21292 21824 21344
rect 21876 21332 21882 21344
rect 23106 21332 23112 21344
rect 21876 21304 23112 21332
rect 21876 21292 21882 21304
rect 23106 21292 23112 21304
rect 23164 21292 23170 21344
rect 23290 21292 23296 21344
rect 23348 21292 23354 21344
rect 26418 21292 26424 21344
rect 26476 21332 26482 21344
rect 27433 21335 27491 21341
rect 27433 21332 27445 21335
rect 26476 21304 27445 21332
rect 26476 21292 26482 21304
rect 27433 21301 27445 21304
rect 27479 21301 27491 21335
rect 27433 21295 27491 21301
rect 27522 21292 27528 21344
rect 27580 21292 27586 21344
rect 27614 21292 27620 21344
rect 27672 21292 27678 21344
rect 28920 21341 28948 21372
rect 28905 21335 28963 21341
rect 28905 21301 28917 21335
rect 28951 21301 28963 21335
rect 28905 21295 28963 21301
rect 1104 21242 35248 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 35248 21242
rect 1104 21168 35248 21190
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 3421 21131 3479 21137
rect 3421 21128 3433 21131
rect 3200 21100 3433 21128
rect 3200 21088 3206 21100
rect 3421 21097 3433 21100
rect 3467 21097 3479 21131
rect 3421 21091 3479 21097
rect 4890 21088 4896 21140
rect 4948 21128 4954 21140
rect 4985 21131 5043 21137
rect 4985 21128 4997 21131
rect 4948 21100 4997 21128
rect 4948 21088 4954 21100
rect 4985 21097 4997 21100
rect 5031 21128 5043 21131
rect 5350 21128 5356 21140
rect 5031 21100 5356 21128
rect 5031 21097 5043 21100
rect 4985 21091 5043 21097
rect 5350 21088 5356 21100
rect 5408 21088 5414 21140
rect 6638 21088 6644 21140
rect 6696 21088 6702 21140
rect 6730 21088 6736 21140
rect 6788 21088 6794 21140
rect 8481 21131 8539 21137
rect 8481 21097 8493 21131
rect 8527 21128 8539 21131
rect 8846 21128 8852 21140
rect 8527 21100 8852 21128
rect 8527 21097 8539 21100
rect 8481 21091 8539 21097
rect 8846 21088 8852 21100
rect 8904 21088 8910 21140
rect 10229 21131 10287 21137
rect 10229 21097 10241 21131
rect 10275 21128 10287 21131
rect 10318 21128 10324 21140
rect 10275 21100 10324 21128
rect 10275 21097 10287 21100
rect 10229 21091 10287 21097
rect 10318 21088 10324 21100
rect 10376 21128 10382 21140
rect 10505 21131 10563 21137
rect 10505 21128 10517 21131
rect 10376 21100 10517 21128
rect 10376 21088 10382 21100
rect 10505 21097 10517 21100
rect 10551 21097 10563 21131
rect 10505 21091 10563 21097
rect 10781 21131 10839 21137
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 10870 21128 10876 21140
rect 10827 21100 10876 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 1670 20952 1676 21004
rect 1728 20952 1734 21004
rect 4798 20952 4804 21004
rect 4856 20992 4862 21004
rect 6362 20992 6368 21004
rect 4856 20964 6368 20992
rect 4856 20952 4862 20964
rect 6362 20952 6368 20964
rect 6420 20952 6426 21004
rect 6748 20992 6776 21088
rect 6472 20964 6776 20992
rect 1394 20884 1400 20936
rect 1452 20884 1458 20936
rect 6472 20933 6500 20964
rect 6457 20927 6515 20933
rect 6457 20893 6469 20927
rect 6503 20893 6515 20927
rect 6457 20887 6515 20893
rect 6546 20884 6552 20936
rect 6604 20884 6610 20936
rect 6730 20884 6736 20936
rect 6788 20884 6794 20936
rect 10520 20924 10548 21091
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 11882 21088 11888 21140
rect 11940 21088 11946 21140
rect 11974 21088 11980 21140
rect 12032 21128 12038 21140
rect 12434 21128 12440 21140
rect 12032 21100 12440 21128
rect 12032 21088 12038 21100
rect 12434 21088 12440 21100
rect 12492 21128 12498 21140
rect 12618 21128 12624 21140
rect 12492 21100 12624 21128
rect 12492 21088 12498 21100
rect 12618 21088 12624 21100
rect 12676 21088 12682 21140
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 13817 21131 13875 21137
rect 13817 21128 13829 21131
rect 13188 21100 13829 21128
rect 11701 21063 11759 21069
rect 11701 21029 11713 21063
rect 11747 21060 11759 21063
rect 11900 21060 11928 21088
rect 11747 21032 11928 21060
rect 11747 21029 11759 21032
rect 11701 21023 11759 21029
rect 10781 20995 10839 21001
rect 10781 20961 10793 20995
rect 10827 20992 10839 20995
rect 10962 20992 10968 21004
rect 10827 20964 10968 20992
rect 10827 20961 10839 20964
rect 10781 20955 10839 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 11072 20964 11560 20992
rect 10873 20927 10931 20933
rect 10873 20924 10885 20927
rect 10520 20896 10885 20924
rect 10873 20893 10885 20896
rect 10919 20924 10931 20927
rect 11072 20924 11100 20964
rect 10919 20896 11100 20924
rect 11149 20927 11207 20933
rect 10919 20893 10931 20896
rect 10873 20887 10931 20893
rect 11149 20893 11161 20927
rect 11195 20924 11207 20927
rect 11241 20927 11299 20933
rect 11241 20924 11253 20927
rect 11195 20896 11253 20924
rect 11195 20893 11207 20896
rect 11149 20887 11207 20893
rect 11241 20893 11253 20896
rect 11287 20924 11299 20927
rect 11330 20924 11336 20936
rect 11287 20896 11336 20924
rect 11287 20893 11299 20896
rect 11241 20887 11299 20893
rect 11330 20884 11336 20896
rect 11388 20884 11394 20936
rect 11425 20927 11483 20933
rect 11425 20893 11437 20927
rect 11471 20893 11483 20927
rect 11532 20924 11560 20964
rect 12710 20952 12716 21004
rect 12768 20952 12774 21004
rect 12894 20952 12900 21004
rect 12952 20992 12958 21004
rect 13188 20992 13216 21100
rect 13817 21097 13829 21100
rect 13863 21128 13875 21131
rect 13906 21128 13912 21140
rect 13863 21100 13912 21128
rect 13863 21097 13875 21100
rect 13817 21091 13875 21097
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 14277 21131 14335 21137
rect 14277 21097 14289 21131
rect 14323 21097 14335 21131
rect 20438 21128 20444 21140
rect 14277 21091 14335 21097
rect 19812 21100 20444 21128
rect 14292 21060 14320 21091
rect 17862 21060 17868 21072
rect 12952 20964 13216 20992
rect 13464 21032 14320 21060
rect 17328 21032 17868 21060
rect 12952 20952 12958 20964
rect 11793 20927 11851 20933
rect 11793 20924 11805 20927
rect 11532 20896 11805 20924
rect 11425 20887 11483 20893
rect 11793 20893 11805 20896
rect 11839 20893 11851 20927
rect 11793 20887 11851 20893
rect 2222 20816 2228 20868
rect 2280 20816 2286 20868
rect 6564 20856 6592 20884
rect 7009 20859 7067 20865
rect 7009 20856 7021 20859
rect 6564 20828 7021 20856
rect 7009 20825 7021 20828
rect 7055 20825 7067 20859
rect 7009 20819 7067 20825
rect 7742 20816 7748 20868
rect 7800 20816 7806 20868
rect 11440 20856 11468 20887
rect 11882 20884 11888 20936
rect 11940 20924 11946 20936
rect 12728 20924 12756 20952
rect 11940 20896 12756 20924
rect 11940 20884 11946 20896
rect 13262 20884 13268 20936
rect 13320 20884 13326 20936
rect 13464 20933 13492 21032
rect 13630 20952 13636 21004
rect 13688 20952 13694 21004
rect 13814 20952 13820 21004
rect 13872 20952 13878 21004
rect 13449 20927 13507 20933
rect 13449 20893 13461 20927
rect 13495 20893 13507 20927
rect 13449 20887 13507 20893
rect 13541 20927 13599 20933
rect 13541 20893 13553 20927
rect 13587 20893 13599 20927
rect 13832 20924 13860 20952
rect 13909 20927 13967 20933
rect 13909 20924 13921 20927
rect 13832 20896 13921 20924
rect 13541 20887 13599 20893
rect 13909 20893 13921 20896
rect 13955 20893 13967 20927
rect 13909 20887 13967 20893
rect 11348 20828 11836 20856
rect 3145 20791 3203 20797
rect 3145 20757 3157 20791
rect 3191 20788 3203 20791
rect 5258 20788 5264 20800
rect 3191 20760 5264 20788
rect 3191 20757 3203 20760
rect 3145 20751 3203 20757
rect 5258 20748 5264 20760
rect 5316 20748 5322 20800
rect 6730 20748 6736 20800
rect 6788 20788 6794 20800
rect 8938 20788 8944 20800
rect 6788 20760 8944 20788
rect 6788 20748 6794 20760
rect 8938 20748 8944 20760
rect 8996 20788 9002 20800
rect 9125 20791 9183 20797
rect 9125 20788 9137 20791
rect 8996 20760 9137 20788
rect 8996 20748 9002 20760
rect 9125 20757 9137 20760
rect 9171 20757 9183 20791
rect 9125 20751 9183 20757
rect 11057 20791 11115 20797
rect 11057 20757 11069 20791
rect 11103 20788 11115 20791
rect 11348 20788 11376 20828
rect 11808 20800 11836 20828
rect 11974 20816 11980 20868
rect 12032 20856 12038 20868
rect 12250 20856 12256 20868
rect 12032 20828 12256 20856
rect 12032 20816 12038 20828
rect 12250 20816 12256 20828
rect 12308 20856 12314 20868
rect 13464 20856 13492 20887
rect 12308 20828 13492 20856
rect 13556 20856 13584 20887
rect 16666 20884 16672 20936
rect 16724 20884 16730 20936
rect 16853 20927 16911 20933
rect 16853 20893 16865 20927
rect 16899 20924 16911 20927
rect 16899 20896 16988 20924
rect 16899 20893 16911 20896
rect 16853 20887 16911 20893
rect 13633 20859 13691 20865
rect 13633 20856 13645 20859
rect 13556 20828 13645 20856
rect 12308 20816 12314 20828
rect 13633 20825 13645 20828
rect 13679 20856 13691 20859
rect 14245 20859 14303 20865
rect 14245 20856 14257 20859
rect 13679 20828 14257 20856
rect 13679 20825 13691 20828
rect 13633 20819 13691 20825
rect 14245 20825 14257 20828
rect 14291 20825 14303 20859
rect 14245 20819 14303 20825
rect 14366 20816 14372 20868
rect 14424 20856 14430 20868
rect 14461 20859 14519 20865
rect 14461 20856 14473 20859
rect 14424 20828 14473 20856
rect 14424 20816 14430 20828
rect 14461 20825 14473 20828
rect 14507 20825 14519 20859
rect 14461 20819 14519 20825
rect 16960 20800 16988 20896
rect 17126 20884 17132 20936
rect 17184 20884 17190 20936
rect 17328 20933 17356 21032
rect 17862 21020 17868 21032
rect 17920 21020 17926 21072
rect 17773 20995 17831 21001
rect 17773 20961 17785 20995
rect 17819 20992 17831 20995
rect 18417 20995 18475 21001
rect 18417 20992 18429 20995
rect 17819 20964 18429 20992
rect 17819 20961 17831 20964
rect 17773 20955 17831 20961
rect 18417 20961 18429 20964
rect 18463 20961 18475 20995
rect 18417 20955 18475 20961
rect 17313 20927 17371 20933
rect 17313 20893 17325 20927
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17405 20927 17463 20933
rect 17405 20893 17417 20927
rect 17451 20893 17463 20927
rect 17405 20887 17463 20893
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 17586 20924 17592 20936
rect 17543 20896 17592 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 17037 20859 17095 20865
rect 17037 20825 17049 20859
rect 17083 20856 17095 20859
rect 17420 20856 17448 20887
rect 17586 20884 17592 20896
rect 17644 20884 17650 20936
rect 17865 20927 17923 20933
rect 17865 20893 17877 20927
rect 17911 20893 17923 20927
rect 17865 20887 17923 20893
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 17880 20856 17908 20887
rect 17083 20828 17908 20856
rect 17083 20825 17095 20828
rect 17037 20819 17095 20825
rect 11103 20760 11376 20788
rect 11103 20757 11115 20760
rect 11057 20751 11115 20757
rect 11790 20748 11796 20800
rect 11848 20748 11854 20800
rect 12526 20748 12532 20800
rect 12584 20748 12590 20800
rect 13814 20748 13820 20800
rect 13872 20788 13878 20800
rect 14093 20791 14151 20797
rect 14093 20788 14105 20791
rect 13872 20760 14105 20788
rect 13872 20748 13878 20760
rect 14093 20757 14105 20760
rect 14139 20757 14151 20791
rect 14093 20751 14151 20757
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17862 20748 17868 20800
rect 17920 20788 17926 20800
rect 18064 20788 18092 20887
rect 19702 20884 19708 20936
rect 19760 20924 19766 20936
rect 19812 20933 19840 21100
rect 20438 21088 20444 21100
rect 20496 21128 20502 21140
rect 20625 21131 20683 21137
rect 20625 21128 20637 21131
rect 20496 21100 20637 21128
rect 20496 21088 20502 21100
rect 20625 21097 20637 21100
rect 20671 21097 20683 21131
rect 20625 21091 20683 21097
rect 21818 21088 21824 21140
rect 21876 21088 21882 21140
rect 22373 21131 22431 21137
rect 22373 21097 22385 21131
rect 22419 21128 22431 21131
rect 22419 21100 23428 21128
rect 22419 21097 22431 21100
rect 22373 21091 22431 21097
rect 20070 21020 20076 21072
rect 20128 21020 20134 21072
rect 22925 21063 22983 21069
rect 22925 21060 22937 21063
rect 22112 21032 22937 21060
rect 22112 21001 22140 21032
rect 22925 21029 22937 21032
rect 22971 21029 22983 21063
rect 22925 21023 22983 21029
rect 22097 20995 22155 21001
rect 20272 20964 20668 20992
rect 20272 20936 20300 20964
rect 19797 20927 19855 20933
rect 19797 20924 19809 20927
rect 19760 20896 19809 20924
rect 19760 20884 19766 20896
rect 19797 20893 19809 20896
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20924 20223 20927
rect 20254 20924 20260 20936
rect 20211 20896 20260 20924
rect 20211 20893 20223 20896
rect 20165 20887 20223 20893
rect 20254 20884 20260 20896
rect 20312 20884 20318 20936
rect 20640 20933 20668 20964
rect 22097 20961 22109 20995
rect 22143 20961 22155 20995
rect 22649 20995 22707 21001
rect 22649 20992 22661 20995
rect 22097 20955 22155 20961
rect 22388 20964 22661 20992
rect 20533 20927 20591 20933
rect 20533 20893 20545 20927
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 20717 20927 20775 20933
rect 20717 20893 20729 20927
rect 20763 20893 20775 20927
rect 20717 20887 20775 20893
rect 22175 20927 22233 20933
rect 22175 20893 22187 20927
rect 22221 20924 22233 20927
rect 22388 20924 22416 20964
rect 22649 20961 22661 20964
rect 22695 20961 22707 20995
rect 23106 20992 23112 21004
rect 22649 20955 22707 20961
rect 22756 20964 23112 20992
rect 22221 20896 22416 20924
rect 22221 20893 22233 20896
rect 22175 20887 22233 20893
rect 20548 20856 20576 20887
rect 20732 20856 20760 20887
rect 22554 20884 22560 20936
rect 22612 20935 22618 20936
rect 22612 20926 22623 20935
rect 22756 20933 22784 20964
rect 23106 20952 23112 20964
rect 23164 20992 23170 21004
rect 23400 21001 23428 21100
rect 23566 21088 23572 21140
rect 23624 21088 23630 21140
rect 24026 21088 24032 21140
rect 24084 21128 24090 21140
rect 24213 21131 24271 21137
rect 24213 21128 24225 21131
rect 24084 21100 24225 21128
rect 24084 21088 24090 21100
rect 24213 21097 24225 21100
rect 24259 21097 24271 21131
rect 24213 21091 24271 21097
rect 24857 21131 24915 21137
rect 24857 21097 24869 21131
rect 24903 21128 24915 21131
rect 24946 21128 24952 21140
rect 24903 21100 24952 21128
rect 24903 21097 24915 21100
rect 24857 21091 24915 21097
rect 24946 21088 24952 21100
rect 25004 21088 25010 21140
rect 26237 21131 26295 21137
rect 26237 21097 26249 21131
rect 26283 21128 26295 21131
rect 26326 21128 26332 21140
rect 26283 21100 26332 21128
rect 26283 21097 26295 21100
rect 26237 21091 26295 21097
rect 26326 21088 26332 21100
rect 26384 21088 26390 21140
rect 26694 21088 26700 21140
rect 26752 21128 26758 21140
rect 27614 21128 27620 21140
rect 26752 21100 27620 21128
rect 26752 21088 26758 21100
rect 27614 21088 27620 21100
rect 27672 21088 27678 21140
rect 25314 21060 25320 21072
rect 23584 21032 25320 21060
rect 23385 20995 23443 21001
rect 23164 20964 23336 20992
rect 23164 20952 23170 20964
rect 22741 20927 22799 20933
rect 22612 20898 22655 20926
rect 22612 20889 22623 20898
rect 22741 20893 22753 20927
rect 22787 20893 22799 20927
rect 22612 20884 22618 20889
rect 22741 20887 22799 20893
rect 22830 20884 22836 20936
rect 22888 20884 22894 20936
rect 23017 20927 23075 20933
rect 23017 20893 23029 20927
rect 23063 20924 23075 20927
rect 23198 20924 23204 20936
rect 23063 20896 23204 20924
rect 23063 20893 23075 20896
rect 23017 20887 23075 20893
rect 20180 20828 20760 20856
rect 21008 20828 21864 20856
rect 20180 20800 20208 20828
rect 17920 20760 18092 20788
rect 17920 20748 17926 20760
rect 18322 20748 18328 20800
rect 18380 20748 18386 20800
rect 20162 20748 20168 20800
rect 20220 20748 20226 20800
rect 21008 20797 21036 20828
rect 20993 20791 21051 20797
rect 20993 20757 21005 20791
rect 21039 20757 21051 20791
rect 21836 20788 21864 20828
rect 22922 20816 22928 20868
rect 22980 20856 22986 20868
rect 23032 20856 23060 20887
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 23308 20924 23336 20964
rect 23385 20961 23397 20995
rect 23431 20992 23443 20995
rect 23474 20992 23480 21004
rect 23431 20964 23480 20992
rect 23431 20961 23443 20964
rect 23385 20955 23443 20961
rect 23474 20952 23480 20964
rect 23532 20952 23538 21004
rect 23584 20924 23612 21032
rect 25314 21020 25320 21032
rect 25372 21020 25378 21072
rect 23753 20995 23811 21001
rect 23753 20961 23765 20995
rect 23799 20992 23811 20995
rect 23799 20964 24164 20992
rect 23799 20961 23811 20964
rect 23753 20955 23811 20961
rect 24136 20936 24164 20964
rect 24486 20952 24492 21004
rect 24544 20952 24550 21004
rect 26053 20995 26111 21001
rect 26053 20992 26065 20995
rect 24872 20964 26065 20992
rect 24872 20936 24900 20964
rect 26053 20961 26065 20964
rect 26099 20992 26111 20995
rect 34057 20995 34115 21001
rect 26099 20964 26556 20992
rect 26099 20961 26111 20964
rect 26053 20955 26111 20961
rect 23308 20896 23612 20924
rect 23658 20884 23664 20936
rect 23716 20884 23722 20936
rect 23842 20884 23848 20936
rect 23900 20884 23906 20936
rect 23969 20927 24027 20933
rect 23969 20924 23981 20927
rect 23952 20893 23981 20924
rect 24015 20893 24027 20927
rect 23952 20887 24027 20893
rect 22980 20828 23060 20856
rect 23385 20859 23443 20865
rect 22980 20816 22986 20828
rect 23385 20825 23397 20859
rect 23431 20856 23443 20859
rect 23750 20856 23756 20868
rect 23431 20828 23756 20856
rect 23431 20825 23443 20828
rect 23385 20819 23443 20825
rect 23750 20816 23756 20828
rect 23808 20856 23814 20868
rect 23952 20856 23980 20887
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24581 20927 24639 20933
rect 24581 20924 24593 20927
rect 24176 20896 24593 20924
rect 24176 20884 24182 20896
rect 24581 20893 24593 20896
rect 24627 20893 24639 20927
rect 24581 20887 24639 20893
rect 24854 20884 24860 20936
rect 24912 20884 24918 20936
rect 25774 20884 25780 20936
rect 25832 20884 25838 20936
rect 25866 20884 25872 20936
rect 25924 20884 25930 20936
rect 26528 20933 26556 20964
rect 34057 20961 34069 20995
rect 34103 20961 34115 20995
rect 34057 20955 34115 20961
rect 25961 20927 26019 20933
rect 25961 20893 25973 20927
rect 26007 20893 26019 20927
rect 25961 20887 26019 20893
rect 26329 20927 26387 20933
rect 26329 20893 26341 20927
rect 26375 20893 26387 20927
rect 26329 20887 26387 20893
rect 26513 20927 26571 20933
rect 26513 20893 26525 20927
rect 26559 20893 26571 20927
rect 26513 20887 26571 20893
rect 25976 20856 26004 20887
rect 26344 20856 26372 20887
rect 34072 20868 34100 20955
rect 34514 20884 34520 20936
rect 34572 20884 34578 20936
rect 23808 20828 23980 20856
rect 25424 20828 26372 20856
rect 23808 20816 23814 20828
rect 25424 20788 25452 20828
rect 34054 20816 34060 20868
rect 34112 20816 34118 20868
rect 21836 20760 25452 20788
rect 20993 20751 21051 20757
rect 25498 20748 25504 20800
rect 25556 20748 25562 20800
rect 25866 20748 25872 20800
rect 25924 20788 25930 20800
rect 26418 20788 26424 20800
rect 25924 20760 26424 20788
rect 25924 20748 25930 20760
rect 26418 20748 26424 20760
rect 26476 20788 26482 20800
rect 27890 20788 27896 20800
rect 26476 20760 27896 20788
rect 26476 20748 26482 20760
rect 27890 20748 27896 20760
rect 27948 20748 27954 20800
rect 1104 20698 35236 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 35236 20698
rect 1104 20624 35236 20646
rect 9490 20544 9496 20596
rect 9548 20584 9554 20596
rect 11333 20587 11391 20593
rect 9548 20556 9674 20584
rect 9548 20544 9554 20556
rect 9646 20516 9674 20556
rect 11333 20553 11345 20587
rect 11379 20584 11391 20587
rect 11698 20584 11704 20596
rect 11379 20556 11704 20584
rect 11379 20553 11391 20556
rect 11333 20547 11391 20553
rect 11698 20544 11704 20556
rect 11756 20544 11762 20596
rect 13906 20544 13912 20596
rect 13964 20544 13970 20596
rect 14001 20587 14059 20593
rect 14001 20553 14013 20587
rect 14047 20584 14059 20587
rect 14182 20584 14188 20596
rect 14047 20556 14188 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 14182 20544 14188 20556
rect 14240 20544 14246 20596
rect 16684 20556 16988 20584
rect 10686 20516 10692 20528
rect 9646 20488 10692 20516
rect 10686 20476 10692 20488
rect 10744 20516 10750 20528
rect 10965 20519 11023 20525
rect 10965 20516 10977 20519
rect 10744 20488 10977 20516
rect 10744 20476 10750 20488
rect 10965 20485 10977 20488
rect 11011 20516 11023 20519
rect 11514 20516 11520 20528
rect 11011 20488 11520 20516
rect 11011 20485 11023 20488
rect 10965 20479 11023 20485
rect 11514 20476 11520 20488
rect 11572 20476 11578 20528
rect 11790 20476 11796 20528
rect 11848 20476 11854 20528
rect 12268 20488 13216 20516
rect 12268 20460 12296 20488
rect 13188 20460 13216 20488
rect 13262 20476 13268 20528
rect 13320 20516 13326 20528
rect 13449 20519 13507 20525
rect 13449 20516 13461 20519
rect 13320 20488 13461 20516
rect 13320 20476 13326 20488
rect 13449 20485 13461 20488
rect 13495 20516 13507 20519
rect 14366 20516 14372 20528
rect 13495 20488 14372 20516
rect 13495 20485 13507 20488
rect 13449 20479 13507 20485
rect 14366 20476 14372 20488
rect 14424 20476 14430 20528
rect 15102 20476 15108 20528
rect 15160 20516 15166 20528
rect 16684 20525 16712 20556
rect 16485 20519 16543 20525
rect 16485 20516 16497 20519
rect 15160 20488 16497 20516
rect 15160 20476 15166 20488
rect 16485 20485 16497 20488
rect 16531 20516 16543 20519
rect 16669 20519 16727 20525
rect 16669 20516 16681 20519
rect 16531 20488 16681 20516
rect 16531 20485 16543 20488
rect 16485 20479 16543 20485
rect 16669 20485 16681 20488
rect 16715 20485 16727 20519
rect 16669 20479 16727 20485
rect 16850 20476 16856 20528
rect 16908 20476 16914 20528
rect 16960 20516 16988 20556
rect 17126 20544 17132 20596
rect 17184 20584 17190 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17184 20556 17601 20584
rect 17184 20544 17190 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17589 20547 17647 20553
rect 17678 20544 17684 20596
rect 17736 20584 17742 20596
rect 22465 20587 22523 20593
rect 17736 20556 22094 20584
rect 17736 20544 17742 20556
rect 17696 20516 17724 20544
rect 16960 20488 17724 20516
rect 22066 20516 22094 20556
rect 22465 20553 22477 20587
rect 22511 20584 22523 20587
rect 22554 20584 22560 20596
rect 22511 20556 22560 20584
rect 22511 20553 22523 20556
rect 22465 20547 22523 20553
rect 22554 20544 22560 20556
rect 22612 20544 22618 20596
rect 22738 20544 22744 20596
rect 22796 20544 22802 20596
rect 22830 20544 22836 20596
rect 22888 20584 22894 20596
rect 23109 20587 23167 20593
rect 23109 20584 23121 20587
rect 22888 20556 23121 20584
rect 22888 20544 22894 20556
rect 23109 20553 23121 20556
rect 23155 20553 23167 20587
rect 23109 20547 23167 20553
rect 23474 20544 23480 20596
rect 23532 20544 23538 20596
rect 23569 20587 23627 20593
rect 23569 20553 23581 20587
rect 23615 20553 23627 20587
rect 23569 20547 23627 20553
rect 22756 20516 22784 20544
rect 22066 20488 22784 20516
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 3053 20451 3111 20457
rect 3053 20448 3065 20451
rect 2271 20420 3065 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 3053 20417 3065 20420
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 3068 20312 3096 20411
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 12066 20448 12072 20460
rect 11112 20420 12072 20448
rect 11112 20408 11118 20420
rect 12066 20408 12072 20420
rect 12124 20408 12130 20460
rect 12250 20408 12256 20460
rect 12308 20408 12314 20460
rect 12526 20408 12532 20460
rect 12584 20408 12590 20460
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 13906 20448 13912 20460
rect 13228 20420 13912 20448
rect 13228 20408 13234 20420
rect 13906 20408 13912 20420
rect 13964 20408 13970 20460
rect 14182 20408 14188 20460
rect 14240 20408 14246 20460
rect 14274 20408 14280 20460
rect 14332 20408 14338 20460
rect 14458 20408 14464 20460
rect 14516 20408 14522 20460
rect 15289 20451 15347 20457
rect 15289 20417 15301 20451
rect 15335 20448 15347 20451
rect 15470 20448 15476 20460
rect 15335 20420 15476 20448
rect 15335 20417 15347 20420
rect 15289 20411 15347 20417
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 16942 20408 16948 20460
rect 17000 20448 17006 20460
rect 17221 20451 17279 20457
rect 17221 20448 17233 20451
rect 17000 20420 17233 20448
rect 17000 20408 17006 20420
rect 17221 20417 17233 20420
rect 17267 20417 17279 20451
rect 17221 20411 17279 20417
rect 17405 20451 17463 20457
rect 17405 20417 17417 20451
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 23492 20448 23520 20544
rect 23584 20516 23612 20547
rect 24486 20544 24492 20596
rect 24544 20544 24550 20596
rect 25314 20544 25320 20596
rect 25372 20584 25378 20596
rect 25372 20556 26004 20584
rect 25372 20544 25378 20556
rect 23842 20516 23848 20528
rect 23584 20488 23848 20516
rect 23842 20476 23848 20488
rect 23900 20516 23906 20528
rect 24029 20519 24087 20525
rect 24029 20516 24041 20519
rect 23900 20488 24041 20516
rect 23900 20476 23906 20488
rect 24029 20485 24041 20488
rect 24075 20485 24087 20519
rect 24029 20479 24087 20485
rect 25608 20488 25820 20516
rect 23569 20451 23627 20457
rect 23569 20448 23581 20451
rect 23492 20420 23581 20448
rect 20165 20411 20223 20417
rect 23569 20417 23581 20420
rect 23615 20417 23627 20451
rect 23569 20411 23627 20417
rect 11517 20383 11575 20389
rect 11517 20380 11529 20383
rect 10244 20352 11529 20380
rect 3329 20315 3387 20321
rect 3329 20312 3341 20315
rect 2884 20284 3341 20312
rect 2884 20256 2912 20284
rect 3329 20281 3341 20284
rect 3375 20281 3387 20315
rect 3329 20275 3387 20281
rect 10244 20256 10272 20352
rect 11517 20349 11529 20352
rect 11563 20380 11575 20383
rect 12158 20380 12164 20392
rect 11563 20352 12164 20380
rect 11563 20349 11575 20352
rect 11517 20343 11575 20349
rect 12158 20340 12164 20352
rect 12216 20340 12222 20392
rect 12544 20380 12572 20408
rect 14200 20380 14228 20408
rect 12544 20352 14228 20380
rect 14292 20380 14320 20408
rect 14737 20383 14795 20389
rect 14737 20380 14749 20383
rect 14292 20352 14749 20380
rect 2314 20204 2320 20256
rect 2372 20204 2378 20256
rect 2777 20247 2835 20253
rect 2777 20213 2789 20247
rect 2823 20244 2835 20247
rect 2866 20244 2872 20256
rect 2823 20216 2872 20244
rect 2823 20213 2835 20216
rect 2777 20207 2835 20213
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 2961 20247 3019 20253
rect 2961 20213 2973 20247
rect 3007 20244 3019 20247
rect 3050 20244 3056 20256
rect 3007 20216 3056 20244
rect 3007 20213 3019 20216
rect 2961 20207 3019 20213
rect 3050 20204 3056 20216
rect 3108 20204 3114 20256
rect 8665 20247 8723 20253
rect 8665 20213 8677 20247
rect 8711 20244 8723 20247
rect 8938 20244 8944 20256
rect 8711 20216 8944 20244
rect 8711 20213 8723 20216
rect 8665 20207 8723 20213
rect 8938 20204 8944 20216
rect 8996 20204 9002 20256
rect 9490 20204 9496 20256
rect 9548 20244 9554 20256
rect 9769 20247 9827 20253
rect 9769 20244 9781 20247
rect 9548 20216 9781 20244
rect 9548 20204 9554 20216
rect 9769 20213 9781 20216
rect 9815 20213 9827 20247
rect 9769 20207 9827 20213
rect 10226 20204 10232 20256
rect 10284 20204 10290 20256
rect 10502 20204 10508 20256
rect 10560 20244 10566 20256
rect 10597 20247 10655 20253
rect 10597 20244 10609 20247
rect 10560 20216 10609 20244
rect 10560 20204 10566 20216
rect 10597 20213 10609 20216
rect 10643 20244 10655 20247
rect 11238 20244 11244 20256
rect 10643 20216 11244 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 11238 20204 11244 20216
rect 11296 20204 11302 20256
rect 12710 20204 12716 20256
rect 12768 20204 12774 20256
rect 13081 20247 13139 20253
rect 13081 20213 13093 20247
rect 13127 20244 13139 20247
rect 13188 20244 13216 20352
rect 14737 20349 14749 20352
rect 14783 20349 14795 20383
rect 14737 20343 14795 20349
rect 15378 20340 15384 20392
rect 15436 20340 15442 20392
rect 15657 20383 15715 20389
rect 15657 20349 15669 20383
rect 15703 20380 15715 20383
rect 16666 20380 16672 20392
rect 15703 20352 16672 20380
rect 15703 20349 15715 20352
rect 15657 20343 15715 20349
rect 16666 20340 16672 20352
rect 16724 20380 16730 20392
rect 17420 20380 17448 20411
rect 16724 20352 17448 20380
rect 16724 20340 16730 20352
rect 20181 20324 20209 20411
rect 23658 20408 23664 20460
rect 23716 20448 23722 20460
rect 23716 20420 23888 20448
rect 23716 20408 23722 20420
rect 20438 20340 20444 20392
rect 20496 20340 20502 20392
rect 23750 20340 23756 20392
rect 23808 20340 23814 20392
rect 23860 20389 23888 20420
rect 23845 20383 23903 20389
rect 23845 20349 23857 20383
rect 23891 20380 23903 20383
rect 25608 20380 25636 20488
rect 25792 20460 25820 20488
rect 25976 20460 26004 20556
rect 28718 20544 28724 20596
rect 28776 20584 28782 20596
rect 28905 20587 28963 20593
rect 28905 20584 28917 20587
rect 28776 20556 28917 20584
rect 28776 20544 28782 20556
rect 28905 20553 28917 20556
rect 28951 20553 28963 20587
rect 28905 20547 28963 20553
rect 28276 20488 28580 20516
rect 25685 20451 25743 20457
rect 25685 20417 25697 20451
rect 25731 20417 25743 20451
rect 25685 20411 25743 20417
rect 23891 20352 25636 20380
rect 23891 20349 23903 20352
rect 23845 20343 23903 20349
rect 13449 20315 13507 20321
rect 13449 20281 13461 20315
rect 13495 20312 13507 20315
rect 13630 20312 13636 20324
rect 13495 20284 13636 20312
rect 13495 20281 13507 20284
rect 13449 20275 13507 20281
rect 13630 20272 13636 20284
rect 13688 20272 13694 20324
rect 17037 20315 17095 20321
rect 17037 20281 17049 20315
rect 17083 20312 17095 20315
rect 17402 20312 17408 20324
rect 17083 20284 17408 20312
rect 17083 20281 17095 20284
rect 17037 20275 17095 20281
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 20162 20272 20168 20324
rect 20220 20272 20226 20324
rect 20349 20315 20407 20321
rect 20349 20281 20361 20315
rect 20395 20312 20407 20315
rect 20395 20284 23520 20312
rect 20395 20281 20407 20284
rect 20349 20275 20407 20281
rect 13127 20216 13216 20244
rect 13127 20213 13139 20216
rect 13081 20207 13139 20213
rect 14182 20204 14188 20256
rect 14240 20204 14246 20256
rect 14918 20204 14924 20256
rect 14976 20244 14982 20256
rect 16853 20247 16911 20253
rect 16853 20244 16865 20247
rect 14976 20216 16865 20244
rect 14976 20204 14982 20216
rect 16853 20213 16865 20216
rect 16899 20244 16911 20247
rect 17770 20244 17776 20256
rect 16899 20216 17776 20244
rect 16899 20213 16911 20216
rect 16853 20207 16911 20213
rect 17770 20204 17776 20216
rect 17828 20204 17834 20256
rect 20254 20204 20260 20256
rect 20312 20204 20318 20256
rect 22830 20204 22836 20256
rect 22888 20204 22894 20256
rect 23492 20244 23520 20284
rect 23566 20272 23572 20324
rect 23624 20312 23630 20324
rect 23661 20315 23719 20321
rect 23661 20312 23673 20315
rect 23624 20284 23673 20312
rect 23624 20272 23630 20284
rect 23661 20281 23673 20284
rect 23707 20281 23719 20315
rect 23768 20312 23796 20340
rect 24305 20315 24363 20321
rect 24305 20312 24317 20315
rect 23768 20284 24317 20312
rect 23661 20275 23719 20281
rect 24305 20281 24317 20284
rect 24351 20281 24363 20315
rect 25700 20312 25728 20411
rect 25774 20408 25780 20460
rect 25832 20408 25838 20460
rect 25958 20408 25964 20460
rect 26016 20408 26022 20460
rect 27893 20451 27951 20457
rect 27893 20448 27905 20451
rect 26344 20420 27905 20448
rect 25792 20380 25820 20408
rect 26344 20380 26372 20420
rect 27893 20417 27905 20420
rect 27939 20448 27951 20451
rect 28166 20448 28172 20460
rect 27939 20420 28172 20448
rect 27939 20417 27951 20420
rect 27893 20411 27951 20417
rect 28166 20408 28172 20420
rect 28224 20408 28230 20460
rect 25792 20352 26372 20380
rect 26237 20315 26295 20321
rect 26237 20312 26249 20315
rect 24305 20275 24363 20281
rect 25608 20284 26249 20312
rect 25608 20256 25636 20284
rect 26237 20281 26249 20284
rect 26283 20281 26295 20315
rect 26237 20275 26295 20281
rect 24854 20244 24860 20256
rect 23492 20216 24860 20244
rect 24854 20204 24860 20216
rect 24912 20204 24918 20256
rect 25590 20204 25596 20256
rect 25648 20204 25654 20256
rect 25869 20247 25927 20253
rect 25869 20213 25881 20247
rect 25915 20244 25927 20247
rect 26344 20244 26372 20352
rect 27614 20340 27620 20392
rect 27672 20380 27678 20392
rect 27985 20383 28043 20389
rect 27985 20380 27997 20383
rect 27672 20352 27997 20380
rect 27672 20340 27678 20352
rect 27985 20349 27997 20352
rect 28031 20380 28043 20383
rect 28276 20380 28304 20488
rect 28445 20451 28503 20457
rect 28445 20417 28457 20451
rect 28491 20417 28503 20451
rect 28445 20411 28503 20417
rect 28031 20352 28304 20380
rect 28031 20349 28043 20352
rect 27985 20343 28043 20349
rect 28460 20256 28488 20411
rect 25915 20216 26372 20244
rect 25915 20213 25927 20216
rect 25869 20207 25927 20213
rect 28166 20204 28172 20256
rect 28224 20204 28230 20256
rect 28442 20204 28448 20256
rect 28500 20204 28506 20256
rect 28552 20253 28580 20488
rect 28537 20247 28595 20253
rect 28537 20213 28549 20247
rect 28583 20213 28595 20247
rect 28537 20207 28595 20213
rect 1104 20154 35248 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 35248 20154
rect 1104 20080 35248 20102
rect 4706 20000 4712 20052
rect 4764 20000 4770 20052
rect 10686 20000 10692 20052
rect 10744 20000 10750 20052
rect 11054 20000 11060 20052
rect 11112 20000 11118 20052
rect 11330 20000 11336 20052
rect 11388 20040 11394 20052
rect 11517 20043 11575 20049
rect 11517 20040 11529 20043
rect 11388 20012 11529 20040
rect 11388 20000 11394 20012
rect 11517 20009 11529 20012
rect 11563 20009 11575 20043
rect 11974 20040 11980 20052
rect 11517 20003 11575 20009
rect 11624 20012 11980 20040
rect 4430 19972 4436 19984
rect 4172 19944 4436 19972
rect 2038 19864 2044 19916
rect 2096 19864 2102 19916
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 1765 19839 1823 19845
rect 1765 19805 1777 19839
rect 1811 19805 1823 19839
rect 1765 19799 1823 19805
rect 1780 19768 1808 19799
rect 3050 19796 3056 19848
rect 3108 19836 3114 19848
rect 4172 19845 4200 19944
rect 4430 19932 4436 19944
rect 4488 19972 4494 19984
rect 4724 19972 4752 20000
rect 4488 19944 4752 19972
rect 4488 19932 4494 19944
rect 4246 19864 4252 19916
rect 4304 19864 4310 19916
rect 4982 19864 4988 19916
rect 5040 19904 5046 19916
rect 5442 19904 5448 19916
rect 5040 19876 5448 19904
rect 5040 19864 5046 19876
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 8481 19907 8539 19913
rect 8481 19873 8493 19907
rect 8527 19904 8539 19907
rect 8938 19904 8944 19916
rect 8527 19876 8944 19904
rect 8527 19873 8539 19876
rect 8481 19867 8539 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 11333 19907 11391 19913
rect 11333 19873 11345 19907
rect 11379 19904 11391 19907
rect 11624 19904 11652 20012
rect 11974 20000 11980 20012
rect 12032 20000 12038 20052
rect 12710 20040 12716 20052
rect 12360 20012 12716 20040
rect 11379 19876 11652 19904
rect 11701 19907 11759 19913
rect 11379 19873 11391 19876
rect 11333 19867 11391 19873
rect 11701 19873 11713 19907
rect 11747 19904 11759 19907
rect 11974 19904 11980 19916
rect 11747 19876 11980 19904
rect 11747 19873 11759 19876
rect 11701 19867 11759 19873
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 12158 19864 12164 19916
rect 12216 19864 12222 19916
rect 12250 19864 12256 19916
rect 12308 19864 12314 19916
rect 4157 19839 4215 19845
rect 3108 19808 3174 19836
rect 3108 19796 3114 19808
rect 4157 19805 4169 19839
rect 4203 19805 4215 19839
rect 4157 19799 4215 19805
rect 5166 19796 5172 19848
rect 5224 19796 5230 19848
rect 5258 19796 5264 19848
rect 5316 19796 5322 19848
rect 7561 19839 7619 19845
rect 7561 19805 7573 19839
rect 7607 19836 7619 19839
rect 7650 19836 7656 19848
rect 7607 19808 7656 19836
rect 7607 19805 7619 19808
rect 7561 19799 7619 19805
rect 7650 19796 7656 19808
rect 7708 19836 7714 19848
rect 7708 19808 8064 19836
rect 7708 19796 7714 19808
rect 1412 19740 1808 19768
rect 1412 19712 1440 19740
rect 1394 19660 1400 19712
rect 1452 19660 1458 19712
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 1670 19700 1676 19712
rect 1627 19672 1676 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 1670 19660 1676 19672
rect 1728 19660 1734 19712
rect 3513 19703 3571 19709
rect 3513 19669 3525 19703
rect 3559 19700 3571 19703
rect 4154 19700 4160 19712
rect 3559 19672 4160 19700
rect 3559 19669 3571 19672
rect 3513 19663 3571 19669
rect 4154 19660 4160 19672
rect 4212 19660 4218 19712
rect 4525 19703 4583 19709
rect 4525 19669 4537 19703
rect 4571 19700 4583 19703
rect 4890 19700 4896 19712
rect 4571 19672 4896 19700
rect 4571 19669 4583 19672
rect 4525 19663 4583 19669
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 4982 19660 4988 19712
rect 5040 19660 5046 19712
rect 7558 19660 7564 19712
rect 7616 19700 7622 19712
rect 8036 19709 8064 19808
rect 8570 19796 8576 19848
rect 8628 19796 8634 19848
rect 9490 19836 9496 19848
rect 8680 19808 9496 19836
rect 8680 19768 8708 19808
rect 9490 19796 9496 19808
rect 9548 19836 9554 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 9548 19808 10241 19836
rect 9548 19796 9554 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 11238 19796 11244 19848
rect 11296 19796 11302 19848
rect 11425 19839 11483 19845
rect 11425 19805 11437 19839
rect 11471 19836 11483 19839
rect 11514 19836 11520 19848
rect 11471 19808 11520 19836
rect 11471 19805 11483 19808
rect 11425 19799 11483 19805
rect 11514 19796 11520 19808
rect 11572 19836 11578 19848
rect 11790 19836 11796 19848
rect 11572 19808 11796 19836
rect 11572 19796 11578 19808
rect 11790 19796 11796 19808
rect 11848 19836 11854 19848
rect 12268 19836 12296 19864
rect 12360 19845 12388 20012
rect 12710 20000 12716 20012
rect 12768 20000 12774 20052
rect 13170 20000 13176 20052
rect 13228 20000 13234 20052
rect 13354 20000 13360 20052
rect 13412 20000 13418 20052
rect 14182 20000 14188 20052
rect 14240 20000 14246 20052
rect 15289 20043 15347 20049
rect 15289 20009 15301 20043
rect 15335 20040 15347 20043
rect 15378 20040 15384 20052
rect 15335 20012 15384 20040
rect 15335 20009 15347 20012
rect 15289 20003 15347 20009
rect 15378 20000 15384 20012
rect 15436 20000 15442 20052
rect 15470 20000 15476 20052
rect 15528 20040 15534 20052
rect 15565 20043 15623 20049
rect 15565 20040 15577 20043
rect 15528 20012 15577 20040
rect 15528 20000 15534 20012
rect 15565 20009 15577 20012
rect 15611 20009 15623 20043
rect 15565 20003 15623 20009
rect 16669 20043 16727 20049
rect 16669 20009 16681 20043
rect 16715 20040 16727 20043
rect 16850 20040 16856 20052
rect 16715 20012 16856 20040
rect 16715 20009 16727 20012
rect 16669 20003 16727 20009
rect 16850 20000 16856 20012
rect 16908 20000 16914 20052
rect 16942 20000 16948 20052
rect 17000 20040 17006 20052
rect 17129 20043 17187 20049
rect 17129 20040 17141 20043
rect 17000 20012 17141 20040
rect 17000 20000 17006 20012
rect 17129 20009 17141 20012
rect 17175 20009 17187 20043
rect 17129 20003 17187 20009
rect 17589 20043 17647 20049
rect 17589 20009 17601 20043
rect 17635 20040 17647 20043
rect 17678 20040 17684 20052
rect 17635 20012 17684 20040
rect 17635 20009 17647 20012
rect 17589 20003 17647 20009
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 17862 20000 17868 20052
rect 17920 20000 17926 20052
rect 17954 20000 17960 20052
rect 18012 20040 18018 20052
rect 20990 20040 20996 20052
rect 18012 20012 20996 20040
rect 18012 20000 18018 20012
rect 20990 20000 20996 20012
rect 21048 20000 21054 20052
rect 22462 20000 22468 20052
rect 22520 20040 22526 20052
rect 22649 20043 22707 20049
rect 22649 20040 22661 20043
rect 22520 20012 22661 20040
rect 22520 20000 22526 20012
rect 22649 20009 22661 20012
rect 22695 20009 22707 20043
rect 22649 20003 22707 20009
rect 23845 20043 23903 20049
rect 23845 20009 23857 20043
rect 23891 20040 23903 20043
rect 24118 20040 24124 20052
rect 23891 20012 24124 20040
rect 23891 20009 23903 20012
rect 23845 20003 23903 20009
rect 12621 19975 12679 19981
rect 12621 19941 12633 19975
rect 12667 19941 12679 19975
rect 12621 19935 12679 19941
rect 11848 19808 12296 19836
rect 12345 19839 12403 19845
rect 11848 19796 11854 19808
rect 12345 19805 12357 19839
rect 12391 19805 12403 19839
rect 12345 19799 12403 19805
rect 12434 19796 12440 19848
rect 12492 19796 12498 19848
rect 12636 19836 12664 19935
rect 14090 19904 14096 19916
rect 13648 19876 14096 19904
rect 13648 19845 13676 19876
rect 14090 19864 14096 19876
rect 14148 19864 14154 19916
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 12636 19808 13553 19836
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19805 13691 19839
rect 13633 19799 13691 19805
rect 13814 19796 13820 19848
rect 13872 19796 13878 19848
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19836 13967 19839
rect 14200 19836 14228 20000
rect 14737 19975 14795 19981
rect 14737 19941 14749 19975
rect 14783 19972 14795 19975
rect 18601 19975 18659 19981
rect 18601 19972 18613 19975
rect 14783 19944 18613 19972
rect 14783 19941 14795 19944
rect 14737 19935 14795 19941
rect 15102 19864 15108 19916
rect 15160 19904 15166 19916
rect 15160 19876 15516 19904
rect 15160 19864 15166 19876
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 13955 19808 14228 19836
rect 14936 19808 15209 19836
rect 13955 19805 13967 19808
rect 13909 19799 13967 19805
rect 14936 19780 14964 19808
rect 15197 19805 15209 19808
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 15378 19796 15384 19848
rect 15436 19796 15442 19848
rect 15488 19845 15516 19876
rect 15672 19848 15700 19944
rect 16850 19904 16856 19916
rect 16224 19876 16856 19904
rect 15473 19839 15531 19845
rect 15473 19805 15485 19839
rect 15519 19805 15531 19839
rect 15473 19799 15531 19805
rect 15654 19796 15660 19848
rect 15712 19796 15718 19848
rect 16114 19796 16120 19848
rect 16172 19836 16178 19848
rect 16224 19845 16252 19876
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 16960 19845 16988 19944
rect 18601 19941 18613 19944
rect 18647 19972 18659 19975
rect 18782 19972 18788 19984
rect 18647 19944 18788 19972
rect 18647 19941 18659 19944
rect 18601 19935 18659 19941
rect 18782 19932 18788 19944
rect 18840 19932 18846 19984
rect 20441 19975 20499 19981
rect 20441 19972 20453 19975
rect 20088 19944 20453 19972
rect 17221 19907 17279 19913
rect 17221 19873 17233 19907
rect 17267 19904 17279 19907
rect 19058 19904 19064 19916
rect 17267 19876 19064 19904
rect 17267 19873 17279 19876
rect 17221 19867 17279 19873
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 16172 19808 16221 19836
rect 16172 19796 16178 19808
rect 16209 19805 16221 19808
rect 16255 19805 16267 19839
rect 16209 19799 16267 19805
rect 16485 19839 16543 19845
rect 16485 19805 16497 19839
rect 16531 19836 16543 19839
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16531 19808 16773 19836
rect 16531 19805 16543 19808
rect 16485 19799 16543 19805
rect 16761 19805 16773 19808
rect 16807 19805 16819 19839
rect 16761 19799 16819 19805
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 8496 19740 8708 19768
rect 8496 19712 8524 19740
rect 9030 19728 9036 19780
rect 9088 19728 9094 19780
rect 9861 19771 9919 19777
rect 9861 19737 9873 19771
rect 9907 19768 9919 19771
rect 12250 19768 12256 19780
rect 9907 19740 12256 19768
rect 9907 19737 9919 19740
rect 9861 19731 9919 19737
rect 12250 19728 12256 19740
rect 12308 19728 12314 19780
rect 12621 19771 12679 19777
rect 12621 19737 12633 19771
rect 12667 19768 12679 19771
rect 13446 19768 13452 19780
rect 12667 19740 13452 19768
rect 12667 19737 12679 19740
rect 12621 19731 12679 19737
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 14918 19728 14924 19780
rect 14976 19728 14982 19780
rect 7653 19703 7711 19709
rect 7653 19700 7665 19703
rect 7616 19672 7665 19700
rect 7616 19660 7622 19672
rect 7653 19669 7665 19672
rect 7699 19669 7711 19703
rect 7653 19663 7711 19669
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8478 19700 8484 19712
rect 8067 19672 8484 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8478 19660 8484 19672
rect 8536 19660 8542 19712
rect 8754 19660 8760 19712
rect 8812 19660 8818 19712
rect 10134 19660 10140 19712
rect 10192 19660 10198 19712
rect 12158 19660 12164 19712
rect 12216 19700 12222 19712
rect 14277 19703 14335 19709
rect 14277 19700 14289 19703
rect 12216 19672 14289 19700
rect 12216 19660 12222 19672
rect 14277 19669 14289 19672
rect 14323 19700 14335 19703
rect 14458 19700 14464 19712
rect 14323 19672 14464 19700
rect 14323 19669 14335 19672
rect 14277 19663 14335 19669
rect 14458 19660 14464 19672
rect 14516 19660 14522 19712
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 15436 19672 16129 19700
rect 15436 19660 15442 19672
rect 16117 19669 16129 19672
rect 16163 19700 16175 19703
rect 16206 19700 16212 19712
rect 16163 19672 16212 19700
rect 16163 19669 16175 19672
rect 16117 19663 16175 19669
rect 16206 19660 16212 19672
rect 16264 19700 16270 19712
rect 16301 19703 16359 19709
rect 16301 19700 16313 19703
rect 16264 19672 16313 19700
rect 16264 19660 16270 19672
rect 16301 19669 16313 19672
rect 16347 19700 16359 19703
rect 17236 19700 17264 19867
rect 19058 19864 19064 19876
rect 19116 19864 19122 19916
rect 17678 19796 17684 19848
rect 17736 19796 17742 19848
rect 17770 19796 17776 19848
rect 17828 19796 17834 19848
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 20088 19845 20116 19944
rect 20441 19941 20453 19944
rect 20487 19941 20499 19975
rect 20441 19935 20499 19941
rect 20254 19864 20260 19916
rect 20312 19864 20318 19916
rect 20349 19907 20407 19913
rect 20349 19873 20361 19907
rect 20395 19904 20407 19907
rect 20806 19904 20812 19916
rect 20395 19876 20812 19904
rect 20395 19873 20407 19876
rect 20349 19867 20407 19873
rect 20806 19864 20812 19876
rect 20864 19904 20870 19916
rect 22664 19904 22692 20003
rect 24118 20000 24124 20012
rect 24176 20000 24182 20052
rect 25777 20043 25835 20049
rect 25777 20009 25789 20043
rect 25823 20040 25835 20043
rect 25823 20012 26188 20040
rect 25823 20009 25835 20012
rect 25777 20003 25835 20009
rect 24029 19975 24087 19981
rect 24029 19972 24041 19975
rect 23584 19944 24041 19972
rect 22922 19904 22928 19916
rect 20864 19876 21956 19904
rect 22664 19876 22928 19904
rect 20864 19864 20870 19876
rect 21928 19848 21956 19876
rect 22922 19864 22928 19876
rect 22980 19904 22986 19916
rect 23584 19913 23612 19944
rect 24029 19941 24041 19944
rect 24075 19941 24087 19975
rect 26050 19972 26056 19984
rect 24029 19935 24087 19941
rect 25516 19944 26056 19972
rect 25516 19916 25544 19944
rect 23109 19907 23167 19913
rect 22980 19876 23060 19904
rect 22980 19864 22986 19876
rect 19521 19839 19579 19845
rect 19521 19836 19533 19839
rect 19392 19808 19533 19836
rect 19392 19796 19398 19808
rect 19521 19805 19533 19808
rect 19567 19805 19579 19839
rect 19521 19799 19579 19805
rect 19797 19839 19855 19845
rect 19797 19805 19809 19839
rect 19843 19805 19855 19839
rect 20073 19839 20131 19845
rect 20073 19836 20085 19839
rect 19797 19799 19855 19805
rect 19996 19808 20085 19836
rect 17954 19728 17960 19780
rect 18012 19728 18018 19780
rect 19812 19768 19840 19799
rect 19444 19740 19840 19768
rect 19444 19712 19472 19740
rect 19996 19712 20024 19808
rect 20073 19805 20085 19808
rect 20119 19805 20131 19839
rect 20073 19799 20131 19805
rect 20622 19796 20628 19848
rect 20680 19796 20686 19848
rect 20714 19796 20720 19848
rect 20772 19836 20778 19848
rect 20898 19836 20904 19848
rect 20772 19808 20904 19836
rect 20772 19796 20778 19808
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21910 19796 21916 19848
rect 21968 19796 21974 19848
rect 22738 19796 22744 19848
rect 22796 19796 22802 19848
rect 23032 19845 23060 19876
rect 23109 19873 23121 19907
rect 23155 19904 23167 19907
rect 23569 19907 23627 19913
rect 23155 19876 23520 19904
rect 23155 19873 23167 19876
rect 23109 19867 23167 19873
rect 23492 19845 23520 19876
rect 23569 19873 23581 19907
rect 23615 19873 23627 19907
rect 25498 19904 25504 19916
rect 23569 19867 23627 19873
rect 23676 19876 25504 19904
rect 23676 19848 23704 19876
rect 23017 19839 23075 19845
rect 23017 19805 23029 19839
rect 23063 19805 23075 19839
rect 23017 19799 23075 19805
rect 23201 19839 23259 19845
rect 23201 19805 23213 19839
rect 23247 19805 23259 19839
rect 23201 19799 23259 19805
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19805 23535 19839
rect 23477 19799 23535 19805
rect 20441 19771 20499 19777
rect 20441 19737 20453 19771
rect 20487 19768 20499 19771
rect 21082 19768 21088 19780
rect 20487 19740 21088 19768
rect 20487 19737 20499 19740
rect 20441 19731 20499 19737
rect 21082 19728 21088 19740
rect 21140 19728 21146 19780
rect 22756 19768 22784 19796
rect 23216 19768 23244 19799
rect 23658 19796 23664 19848
rect 23716 19796 23722 19848
rect 24136 19845 24164 19876
rect 25498 19864 25504 19876
rect 25556 19864 25562 19916
rect 23937 19839 23995 19845
rect 23937 19805 23949 19839
rect 23983 19805 23995 19839
rect 23937 19799 23995 19805
rect 24121 19839 24179 19845
rect 24121 19805 24133 19839
rect 24167 19805 24179 19839
rect 24121 19799 24179 19805
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25409 19839 25467 19845
rect 25409 19836 25421 19839
rect 25179 19808 25421 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 25409 19805 25421 19808
rect 25455 19805 25467 19839
rect 25409 19799 25467 19805
rect 22756 19740 23244 19768
rect 23290 19728 23296 19780
rect 23348 19768 23354 19780
rect 23952 19768 23980 19799
rect 24581 19771 24639 19777
rect 24581 19768 24593 19771
rect 23348 19740 24593 19768
rect 23348 19728 23354 19740
rect 24581 19737 24593 19740
rect 24627 19737 24639 19771
rect 24581 19731 24639 19737
rect 16347 19672 17264 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 19426 19660 19432 19712
rect 19484 19660 19490 19712
rect 19978 19660 19984 19712
rect 20036 19660 20042 19712
rect 22094 19660 22100 19712
rect 22152 19700 22158 19712
rect 22830 19700 22836 19712
rect 22152 19672 22836 19700
rect 22152 19660 22158 19672
rect 22830 19660 22836 19672
rect 22888 19700 22894 19712
rect 25424 19700 25452 19799
rect 25590 19796 25596 19848
rect 25648 19796 25654 19848
rect 25685 19839 25743 19845
rect 25685 19805 25697 19839
rect 25731 19836 25743 19839
rect 25774 19836 25780 19848
rect 25731 19808 25780 19836
rect 25731 19805 25743 19808
rect 25685 19799 25743 19805
rect 25774 19796 25780 19808
rect 25832 19796 25838 19848
rect 25869 19839 25927 19845
rect 25869 19805 25881 19839
rect 25915 19838 25927 19839
rect 25976 19838 26004 19944
rect 26050 19932 26056 19944
rect 26108 19932 26114 19984
rect 25915 19810 26004 19838
rect 26053 19839 26111 19845
rect 25915 19805 25927 19810
rect 25869 19799 25927 19805
rect 26053 19805 26065 19839
rect 26099 19805 26111 19839
rect 26160 19836 26188 20012
rect 28166 20000 28172 20052
rect 28224 20000 28230 20052
rect 34514 20000 34520 20052
rect 34572 20000 34578 20052
rect 27893 19975 27951 19981
rect 27893 19941 27905 19975
rect 27939 19941 27951 19975
rect 27893 19935 27951 19941
rect 27065 19907 27123 19913
rect 27065 19873 27077 19907
rect 27111 19904 27123 19907
rect 27522 19904 27528 19916
rect 27111 19876 27528 19904
rect 27111 19873 27123 19876
rect 27065 19867 27123 19873
rect 27522 19864 27528 19876
rect 27580 19864 27586 19916
rect 26237 19839 26295 19845
rect 26237 19836 26249 19839
rect 26160 19808 26249 19836
rect 26053 19799 26111 19805
rect 26237 19805 26249 19808
rect 26283 19805 26295 19839
rect 27798 19836 27804 19848
rect 27632 19823 27804 19836
rect 26237 19799 26295 19805
rect 27620 19817 27804 19823
rect 25501 19771 25559 19777
rect 25501 19737 25513 19771
rect 25547 19768 25559 19771
rect 26068 19768 26096 19799
rect 27620 19783 27632 19817
rect 27666 19808 27804 19817
rect 27666 19783 27678 19808
rect 27798 19796 27804 19808
rect 27856 19796 27862 19848
rect 27908 19836 27936 19935
rect 28184 19904 28212 20000
rect 32585 19975 32643 19981
rect 32585 19972 32597 19975
rect 31036 19944 32597 19972
rect 28721 19907 28779 19913
rect 28721 19904 28733 19907
rect 28184 19876 28733 19904
rect 28721 19873 28733 19876
rect 28767 19873 28779 19907
rect 28721 19867 28779 19873
rect 29638 19864 29644 19916
rect 29696 19904 29702 19916
rect 29733 19907 29791 19913
rect 29733 19904 29745 19907
rect 29696 19876 29745 19904
rect 29696 19864 29702 19876
rect 29733 19873 29745 19876
rect 29779 19904 29791 19907
rect 31036 19904 31064 19944
rect 32585 19941 32597 19944
rect 32631 19972 32643 19975
rect 32674 19972 32680 19984
rect 32631 19944 32680 19972
rect 32631 19941 32643 19944
rect 32585 19935 32643 19941
rect 32674 19932 32680 19944
rect 32732 19972 32738 19984
rect 32732 19944 32812 19972
rect 32732 19932 32738 19944
rect 29779 19876 31064 19904
rect 31481 19907 31539 19913
rect 29779 19873 29791 19876
rect 29733 19867 29791 19873
rect 31481 19873 31493 19907
rect 31527 19904 31539 19907
rect 31527 19876 31754 19904
rect 31527 19873 31539 19876
rect 31481 19867 31539 19873
rect 28442 19836 28448 19848
rect 27908 19808 28448 19836
rect 28442 19796 28448 19808
rect 28500 19836 28506 19848
rect 28813 19839 28871 19845
rect 28813 19836 28825 19839
rect 28500 19808 28825 19836
rect 28500 19796 28506 19808
rect 28813 19805 28825 19808
rect 28859 19805 28871 19839
rect 31726 19836 31754 19876
rect 31846 19864 31852 19916
rect 31904 19864 31910 19916
rect 32784 19913 32812 19944
rect 32769 19907 32827 19913
rect 32769 19873 32781 19907
rect 32815 19873 32827 19907
rect 32769 19867 32827 19873
rect 31941 19839 31999 19845
rect 31941 19836 31953 19839
rect 31726 19808 31953 19836
rect 28813 19799 28871 19805
rect 31941 19805 31953 19808
rect 31987 19836 31999 19839
rect 32122 19836 32128 19848
rect 31987 19808 32128 19836
rect 31987 19805 31999 19808
rect 31941 19799 31999 19805
rect 32122 19796 32128 19808
rect 32180 19796 32186 19848
rect 34514 19796 34520 19848
rect 34572 19836 34578 19848
rect 34701 19839 34759 19845
rect 34701 19836 34713 19839
rect 34572 19808 34713 19836
rect 34572 19796 34578 19808
rect 34701 19805 34713 19808
rect 34747 19805 34759 19839
rect 34701 19799 34759 19805
rect 27620 19780 27678 19783
rect 25547 19740 26096 19768
rect 25547 19737 25559 19740
rect 25501 19731 25559 19737
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 27614 19728 27620 19780
rect 27672 19728 27678 19780
rect 27890 19728 27896 19780
rect 27948 19728 27954 19780
rect 30009 19771 30067 19777
rect 30009 19768 30021 19771
rect 29196 19740 30021 19768
rect 26620 19700 26648 19728
rect 22888 19672 26648 19700
rect 27709 19703 27767 19709
rect 22888 19660 22894 19672
rect 27709 19669 27721 19703
rect 27755 19700 27767 19703
rect 27798 19700 27804 19712
rect 27755 19672 27804 19700
rect 27755 19669 27767 19672
rect 27709 19663 27767 19669
rect 27798 19660 27804 19672
rect 27856 19660 27862 19712
rect 29196 19709 29224 19740
rect 30009 19737 30021 19740
rect 30055 19737 30067 19771
rect 30009 19731 30067 19737
rect 30742 19728 30748 19780
rect 30800 19728 30806 19780
rect 33045 19771 33103 19777
rect 33045 19768 33057 19771
rect 32324 19740 33057 19768
rect 32324 19709 32352 19740
rect 33045 19737 33057 19740
rect 33091 19737 33103 19771
rect 34793 19771 34851 19777
rect 34793 19768 34805 19771
rect 34270 19740 34805 19768
rect 33045 19731 33103 19737
rect 34793 19737 34805 19740
rect 34839 19737 34851 19771
rect 34793 19731 34851 19737
rect 29181 19703 29239 19709
rect 29181 19669 29193 19703
rect 29227 19669 29239 19703
rect 29181 19663 29239 19669
rect 32309 19703 32367 19709
rect 32309 19669 32321 19703
rect 32355 19669 32367 19703
rect 32309 19663 32367 19669
rect 1104 19610 35236 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 35236 19610
rect 1104 19536 35236 19558
rect 4246 19456 4252 19508
rect 4304 19456 4310 19508
rect 4706 19456 4712 19508
rect 4764 19496 4770 19508
rect 5166 19496 5172 19508
rect 4764 19468 5172 19496
rect 4764 19456 4770 19468
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 5261 19499 5319 19505
rect 5261 19465 5273 19499
rect 5307 19496 5319 19499
rect 8570 19496 8576 19508
rect 5307 19468 8576 19496
rect 5307 19465 5319 19468
rect 5261 19459 5319 19465
rect 8570 19456 8576 19468
rect 8628 19456 8634 19508
rect 11790 19456 11796 19508
rect 11848 19456 11854 19508
rect 12066 19456 12072 19508
rect 12124 19496 12130 19508
rect 12802 19496 12808 19508
rect 12124 19468 12808 19496
rect 12124 19456 12130 19468
rect 12802 19456 12808 19468
rect 12860 19456 12866 19508
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19496 13323 19499
rect 13446 19496 13452 19508
rect 13311 19468 13452 19496
rect 13311 19465 13323 19468
rect 13265 19459 13323 19465
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 15654 19456 15660 19508
rect 15712 19456 15718 19508
rect 16117 19499 16175 19505
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 16206 19496 16212 19508
rect 16163 19468 16212 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 16206 19456 16212 19468
rect 16264 19456 16270 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 18012 19468 18245 19496
rect 18012 19456 18018 19468
rect 18233 19465 18245 19468
rect 18279 19465 18291 19499
rect 18233 19459 18291 19465
rect 18601 19499 18659 19505
rect 18601 19465 18613 19499
rect 18647 19465 18659 19499
rect 18601 19459 18659 19465
rect 2314 19388 2320 19440
rect 2372 19388 2378 19440
rect 4154 19428 4160 19440
rect 3988 19400 4160 19428
rect 1394 19320 1400 19372
rect 1452 19320 1458 19372
rect 3988 19369 4016 19400
rect 4154 19388 4160 19400
rect 4212 19428 4218 19440
rect 4212 19400 4476 19428
rect 4212 19388 4218 19400
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19329 4031 19363
rect 3973 19323 4031 19329
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19329 4399 19363
rect 4341 19323 4399 19329
rect 1673 19295 1731 19301
rect 1673 19261 1685 19295
rect 1719 19292 1731 19295
rect 1762 19292 1768 19304
rect 1719 19264 1768 19292
rect 1719 19261 1731 19264
rect 1673 19255 1731 19261
rect 1762 19252 1768 19264
rect 1820 19252 1826 19304
rect 4249 19295 4307 19301
rect 4249 19292 4261 19295
rect 3988 19264 4261 19292
rect 3605 19227 3663 19233
rect 3605 19224 3617 19227
rect 3068 19196 3617 19224
rect 3068 19168 3096 19196
rect 3605 19193 3617 19196
rect 3651 19193 3663 19227
rect 3605 19187 3663 19193
rect 3988 19168 4016 19264
rect 4249 19261 4261 19264
rect 4295 19261 4307 19295
rect 4249 19255 4307 19261
rect 4065 19227 4123 19233
rect 4065 19193 4077 19227
rect 4111 19224 4123 19227
rect 4356 19224 4384 19323
rect 4448 19301 4476 19400
rect 4982 19388 4988 19440
rect 5040 19388 5046 19440
rect 6730 19428 6736 19440
rect 6564 19400 6736 19428
rect 5000 19360 5028 19388
rect 6564 19372 6592 19400
rect 6730 19388 6736 19400
rect 6788 19388 6794 19440
rect 8481 19431 8539 19437
rect 8481 19428 8493 19431
rect 8050 19400 8493 19428
rect 8481 19397 8493 19400
rect 8527 19397 8539 19431
rect 8481 19391 8539 19397
rect 8754 19388 8760 19440
rect 8812 19428 8818 19440
rect 9125 19431 9183 19437
rect 9125 19428 9137 19431
rect 8812 19400 9137 19428
rect 8812 19388 8818 19400
rect 9125 19397 9137 19400
rect 9171 19397 9183 19431
rect 9125 19391 9183 19397
rect 10134 19388 10140 19440
rect 10192 19388 10198 19440
rect 11238 19388 11244 19440
rect 11296 19428 11302 19440
rect 11974 19428 11980 19440
rect 11296 19400 11980 19428
rect 11296 19388 11302 19400
rect 11974 19388 11980 19400
rect 12032 19428 12038 19440
rect 12437 19431 12495 19437
rect 12437 19428 12449 19431
rect 12032 19400 12449 19428
rect 12032 19388 12038 19400
rect 12437 19397 12449 19400
rect 12483 19428 12495 19431
rect 12526 19428 12532 19440
rect 12483 19400 12532 19428
rect 12483 19397 12495 19400
rect 12437 19391 12495 19397
rect 12526 19388 12532 19400
rect 12584 19388 12590 19440
rect 15672 19428 15700 19456
rect 16390 19428 16396 19440
rect 15672 19400 16396 19428
rect 16390 19388 16396 19400
rect 16448 19388 16454 19440
rect 17678 19388 17684 19440
rect 17736 19428 17742 19440
rect 18616 19428 18644 19459
rect 18782 19456 18788 19508
rect 18840 19496 18846 19508
rect 18840 19468 19196 19496
rect 18840 19456 18846 19468
rect 17736 19400 18644 19428
rect 17736 19388 17742 19400
rect 19058 19388 19064 19440
rect 19116 19388 19122 19440
rect 5077 19363 5135 19369
rect 5077 19360 5089 19363
rect 5000 19332 5089 19360
rect 5077 19329 5089 19332
rect 5123 19329 5135 19363
rect 5077 19323 5135 19329
rect 5258 19320 5264 19372
rect 5316 19360 5322 19372
rect 5537 19363 5595 19369
rect 5537 19360 5549 19363
rect 5316 19332 5549 19360
rect 5316 19320 5322 19332
rect 5537 19329 5549 19332
rect 5583 19329 5595 19363
rect 5537 19323 5595 19329
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 8573 19363 8631 19369
rect 8573 19360 8585 19363
rect 8496 19332 8585 19360
rect 8496 19304 8524 19332
rect 8573 19329 8585 19332
rect 8619 19329 8631 19363
rect 8573 19323 8631 19329
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 11514 19360 11520 19372
rect 10919 19332 11520 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19360 17463 19363
rect 17862 19360 17868 19372
rect 17451 19332 17868 19360
rect 17451 19329 17463 19332
rect 17405 19323 17463 19329
rect 17862 19320 17868 19332
rect 17920 19360 17926 19372
rect 18785 19363 18843 19369
rect 18785 19360 18797 19363
rect 17920 19332 18797 19360
rect 17920 19320 17926 19332
rect 18785 19329 18797 19332
rect 18831 19329 18843 19363
rect 18785 19323 18843 19329
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19360 19027 19363
rect 19076 19360 19104 19388
rect 19168 19369 19196 19468
rect 20162 19456 20168 19508
rect 20220 19456 20226 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 20901 19499 20959 19505
rect 20901 19496 20913 19499
rect 20680 19468 20913 19496
rect 20680 19456 20686 19468
rect 20901 19465 20913 19468
rect 20947 19496 20959 19499
rect 21542 19496 21548 19508
rect 20947 19468 21548 19496
rect 20947 19465 20959 19468
rect 20901 19459 20959 19465
rect 21542 19456 21548 19468
rect 21600 19456 21606 19508
rect 21637 19499 21695 19505
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 22021 19499 22079 19505
rect 22021 19496 22033 19499
rect 21683 19468 22033 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 22021 19465 22033 19468
rect 22067 19496 22079 19499
rect 22067 19468 22508 19496
rect 22067 19465 22079 19468
rect 22021 19459 22079 19465
rect 20714 19428 20720 19440
rect 19812 19400 20720 19428
rect 19015 19332 19104 19360
rect 19153 19363 19211 19369
rect 19015 19329 19027 19332
rect 18969 19323 19027 19329
rect 19153 19329 19165 19363
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4798 19292 4804 19304
rect 4479 19264 4804 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 4893 19295 4951 19301
rect 4893 19261 4905 19295
rect 4939 19292 4951 19295
rect 5166 19292 5172 19304
rect 4939 19264 5172 19292
rect 4939 19261 4951 19264
rect 4893 19255 4951 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5626 19252 5632 19304
rect 5684 19252 5690 19304
rect 6825 19295 6883 19301
rect 6825 19292 6837 19295
rect 6656 19264 6837 19292
rect 5905 19227 5963 19233
rect 4111 19196 5028 19224
rect 4111 19193 4123 19196
rect 4065 19187 4123 19193
rect 5000 19168 5028 19196
rect 5905 19193 5917 19227
rect 5951 19224 5963 19227
rect 6656 19224 6684 19264
rect 6825 19261 6837 19264
rect 6871 19261 6883 19295
rect 6825 19255 6883 19261
rect 8478 19252 8484 19304
rect 8536 19252 8542 19304
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19292 8907 19295
rect 8895 19264 8984 19292
rect 8895 19261 8907 19264
rect 8849 19255 8907 19261
rect 5951 19196 6684 19224
rect 5951 19193 5963 19196
rect 5905 19187 5963 19193
rect 8956 19168 8984 19264
rect 14642 19252 14648 19304
rect 14700 19292 14706 19304
rect 15105 19295 15163 19301
rect 15105 19292 15117 19295
rect 14700 19264 15117 19292
rect 14700 19252 14706 19264
rect 15105 19261 15117 19264
rect 15151 19292 15163 19295
rect 15378 19292 15384 19304
rect 15151 19264 15384 19292
rect 15151 19261 15163 19264
rect 15105 19255 15163 19261
rect 15378 19252 15384 19264
rect 15436 19252 15442 19304
rect 17037 19295 17095 19301
rect 17037 19261 17049 19295
rect 17083 19292 17095 19295
rect 18046 19292 18052 19304
rect 17083 19264 18052 19292
rect 17083 19261 17095 19264
rect 17037 19255 17095 19261
rect 18046 19252 18052 19264
rect 18104 19292 18110 19304
rect 18322 19292 18328 19304
rect 18104 19264 18328 19292
rect 18104 19252 18110 19264
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 18414 19252 18420 19304
rect 18472 19252 18478 19304
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 17678 19184 17684 19236
rect 17736 19184 17742 19236
rect 3050 19116 3056 19168
rect 3108 19116 3114 19168
rect 3145 19159 3203 19165
rect 3145 19125 3157 19159
rect 3191 19156 3203 19159
rect 3418 19156 3424 19168
rect 3191 19128 3424 19156
rect 3191 19125 3203 19128
rect 3145 19119 3203 19125
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 3970 19116 3976 19168
rect 4028 19116 4034 19168
rect 4430 19116 4436 19168
rect 4488 19116 4494 19168
rect 4982 19116 4988 19168
rect 5040 19116 5046 19168
rect 5258 19116 5264 19168
rect 5316 19156 5322 19168
rect 5442 19156 5448 19168
rect 5316 19128 5448 19156
rect 5316 19116 5322 19128
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 8294 19116 8300 19168
rect 8352 19116 8358 19168
rect 8938 19116 8944 19168
rect 8996 19116 9002 19168
rect 18141 19159 18199 19165
rect 18141 19125 18153 19159
rect 18187 19156 18199 19159
rect 18322 19156 18328 19168
rect 18187 19128 18328 19156
rect 18187 19125 18199 19128
rect 18141 19119 18199 19125
rect 18322 19116 18328 19128
rect 18380 19156 18386 19168
rect 18524 19156 18552 19255
rect 18690 19252 18696 19304
rect 18748 19292 18754 19304
rect 18892 19292 18920 19323
rect 19334 19320 19340 19372
rect 19392 19360 19398 19372
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19392 19332 19533 19360
rect 19392 19320 19398 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 19812 19369 19840 19400
rect 20714 19388 20720 19400
rect 20772 19388 20778 19440
rect 21269 19431 21327 19437
rect 21269 19397 21281 19431
rect 21315 19428 21327 19431
rect 21821 19431 21879 19437
rect 21821 19428 21833 19431
rect 21315 19400 21833 19428
rect 21315 19397 21327 19400
rect 21269 19391 21327 19397
rect 21821 19397 21833 19400
rect 21867 19428 21879 19431
rect 22373 19431 22431 19437
rect 22373 19428 22385 19431
rect 21867 19400 22385 19428
rect 21867 19397 21879 19400
rect 21821 19391 21879 19397
rect 22373 19397 22385 19400
rect 22419 19397 22431 19431
rect 22373 19391 22431 19397
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19668 19332 19717 19360
rect 19668 19320 19674 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 19978 19360 19984 19372
rect 19935 19332 19984 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 19978 19320 19984 19332
rect 20036 19320 20042 19372
rect 20809 19363 20867 19369
rect 20809 19329 20821 19363
rect 20855 19360 20867 19363
rect 20898 19360 20904 19372
rect 20855 19332 20904 19360
rect 20855 19329 20867 19332
rect 20809 19323 20867 19329
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 21082 19320 21088 19372
rect 21140 19360 21146 19372
rect 21361 19363 21419 19369
rect 21361 19360 21373 19363
rect 21140 19332 21373 19360
rect 21140 19320 21146 19332
rect 21361 19329 21373 19332
rect 21407 19329 21419 19363
rect 21361 19323 21419 19329
rect 21545 19363 21603 19369
rect 21545 19329 21557 19363
rect 21591 19329 21603 19363
rect 21545 19323 21603 19329
rect 18748 19264 18920 19292
rect 20916 19292 20944 19320
rect 21560 19292 21588 19323
rect 21634 19320 21640 19372
rect 21692 19320 21698 19372
rect 22281 19363 22339 19369
rect 22281 19329 22293 19363
rect 22327 19360 22339 19363
rect 22480 19360 22508 19468
rect 22738 19456 22744 19508
rect 22796 19496 22802 19508
rect 22833 19499 22891 19505
rect 22833 19496 22845 19499
rect 22796 19468 22845 19496
rect 22796 19456 22802 19468
rect 22833 19465 22845 19468
rect 22879 19465 22891 19499
rect 22833 19459 22891 19465
rect 23474 19456 23480 19508
rect 23532 19496 23538 19508
rect 23569 19499 23627 19505
rect 23569 19496 23581 19499
rect 23532 19468 23581 19496
rect 23532 19456 23538 19468
rect 23569 19465 23581 19468
rect 23615 19465 23627 19499
rect 23569 19459 23627 19465
rect 25958 19456 25964 19508
rect 26016 19496 26022 19508
rect 26145 19499 26203 19505
rect 26145 19496 26157 19499
rect 26016 19468 26157 19496
rect 26016 19456 26022 19468
rect 26145 19465 26157 19468
rect 26191 19465 26203 19499
rect 26145 19459 26203 19465
rect 29638 19456 29644 19508
rect 29696 19456 29702 19508
rect 30742 19456 30748 19508
rect 30800 19456 30806 19508
rect 31846 19456 31852 19508
rect 31904 19496 31910 19508
rect 31941 19499 31999 19505
rect 31941 19496 31953 19499
rect 31904 19468 31953 19496
rect 31904 19456 31910 19468
rect 31941 19465 31953 19468
rect 31987 19465 31999 19499
rect 31941 19459 31999 19465
rect 32490 19456 32496 19508
rect 32548 19456 32554 19508
rect 25593 19431 25651 19437
rect 25593 19397 25605 19431
rect 25639 19428 25651 19431
rect 26418 19428 26424 19440
rect 25639 19400 26424 19428
rect 25639 19397 25651 19400
rect 25593 19391 25651 19397
rect 26418 19388 26424 19400
rect 26476 19388 26482 19440
rect 22327 19332 22508 19360
rect 22557 19363 22615 19369
rect 22327 19329 22339 19332
rect 22281 19323 22339 19329
rect 22557 19329 22569 19363
rect 22603 19329 22615 19363
rect 22557 19323 22615 19329
rect 22094 19292 22100 19304
rect 20916 19264 21588 19292
rect 21652 19264 22100 19292
rect 18748 19252 18754 19264
rect 19058 19184 19064 19236
rect 19116 19184 19122 19236
rect 21652 19156 21680 19264
rect 22094 19252 22100 19264
rect 22152 19252 22158 19304
rect 22572 19292 22600 19323
rect 22922 19320 22928 19372
rect 22980 19360 22986 19372
rect 25225 19363 25283 19369
rect 25225 19360 25237 19363
rect 22980 19332 25237 19360
rect 22980 19320 22986 19332
rect 25225 19329 25237 19332
rect 25271 19329 25283 19363
rect 25225 19323 25283 19329
rect 25869 19363 25927 19369
rect 25869 19329 25881 19363
rect 25915 19360 25927 19363
rect 26694 19360 26700 19372
rect 25915 19332 26700 19360
rect 25915 19329 25927 19332
rect 25869 19323 25927 19329
rect 22480 19264 22600 19292
rect 25240 19292 25268 19323
rect 26694 19320 26700 19332
rect 26752 19320 26758 19372
rect 30650 19360 30656 19372
rect 30484 19332 30656 19360
rect 25590 19292 25596 19304
rect 25240 19264 25596 19292
rect 22480 19224 22508 19264
rect 25590 19252 25596 19264
rect 25648 19292 25654 19304
rect 26513 19295 26571 19301
rect 26513 19292 26525 19295
rect 25648 19264 26525 19292
rect 25648 19252 25654 19264
rect 26513 19261 26525 19264
rect 26559 19261 26571 19295
rect 26513 19255 26571 19261
rect 22020 19196 22508 19224
rect 18380 19128 21680 19156
rect 18380 19116 18386 19128
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 22020 19165 22048 19196
rect 24578 19184 24584 19236
rect 24636 19224 24642 19236
rect 24765 19227 24823 19233
rect 24765 19224 24777 19227
rect 24636 19196 24777 19224
rect 24636 19184 24642 19196
rect 24765 19193 24777 19196
rect 24811 19193 24823 19227
rect 24765 19187 24823 19193
rect 22005 19159 22063 19165
rect 22005 19156 22017 19159
rect 21784 19128 22017 19156
rect 21784 19116 21790 19128
rect 22005 19125 22017 19128
rect 22051 19125 22063 19159
rect 22005 19119 22063 19125
rect 22186 19116 22192 19168
rect 22244 19116 22250 19168
rect 22554 19116 22560 19168
rect 22612 19116 22618 19168
rect 24305 19159 24363 19165
rect 24305 19125 24317 19159
rect 24351 19156 24363 19159
rect 24670 19156 24676 19168
rect 24351 19128 24676 19156
rect 24351 19125 24363 19128
rect 24305 19119 24363 19125
rect 24670 19116 24676 19128
rect 24728 19116 24734 19168
rect 25774 19116 25780 19168
rect 25832 19116 25838 19168
rect 30190 19116 30196 19168
rect 30248 19156 30254 19168
rect 30484 19165 30512 19332
rect 30650 19320 30656 19332
rect 30708 19320 30714 19372
rect 31662 19360 31668 19372
rect 31623 19332 31668 19360
rect 31662 19320 31668 19332
rect 31720 19360 31726 19372
rect 32125 19363 32183 19369
rect 31720 19332 32076 19360
rect 31720 19320 31726 19332
rect 31938 19252 31944 19304
rect 31996 19252 32002 19304
rect 32048 19292 32076 19332
rect 32125 19329 32137 19363
rect 32171 19360 32183 19363
rect 32398 19360 32404 19372
rect 32171 19332 32404 19360
rect 32171 19329 32183 19332
rect 32125 19323 32183 19329
rect 32217 19295 32275 19301
rect 32217 19292 32229 19295
rect 32048 19264 32229 19292
rect 32217 19261 32229 19264
rect 32263 19261 32275 19295
rect 32217 19255 32275 19261
rect 31757 19227 31815 19233
rect 31757 19193 31769 19227
rect 31803 19224 31815 19227
rect 32324 19224 32352 19332
rect 32398 19320 32404 19332
rect 32456 19320 32462 19372
rect 31803 19196 32352 19224
rect 31803 19193 31815 19196
rect 31757 19187 31815 19193
rect 30469 19159 30527 19165
rect 30469 19156 30481 19159
rect 30248 19128 30481 19156
rect 30248 19116 30254 19128
rect 30469 19125 30481 19128
rect 30515 19125 30527 19159
rect 30469 19119 30527 19125
rect 32122 19116 32128 19168
rect 32180 19116 32186 19168
rect 34241 19159 34299 19165
rect 34241 19125 34253 19159
rect 34287 19156 34299 19159
rect 34330 19156 34336 19168
rect 34287 19128 34336 19156
rect 34287 19125 34299 19128
rect 34241 19119 34299 19125
rect 34330 19116 34336 19128
rect 34388 19156 34394 19168
rect 34514 19156 34520 19168
rect 34388 19128 34520 19156
rect 34388 19116 34394 19128
rect 34514 19116 34520 19128
rect 34572 19116 34578 19168
rect 1104 19066 35248 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 35248 19066
rect 1104 18992 35248 19014
rect 4706 18912 4712 18964
rect 4764 18912 4770 18964
rect 4890 18912 4896 18964
rect 4948 18912 4954 18964
rect 5537 18955 5595 18961
rect 5537 18921 5549 18955
rect 5583 18952 5595 18955
rect 5626 18952 5632 18964
rect 5583 18924 5632 18952
rect 5583 18921 5595 18924
rect 5537 18915 5595 18921
rect 5626 18912 5632 18924
rect 5684 18912 5690 18964
rect 8297 18955 8355 18961
rect 8297 18921 8309 18955
rect 8343 18952 8355 18955
rect 9030 18952 9036 18964
rect 8343 18924 9036 18952
rect 8343 18921 8355 18924
rect 8297 18915 8355 18921
rect 9030 18912 9036 18924
rect 9088 18912 9094 18964
rect 10226 18952 10232 18964
rect 9784 18924 10232 18952
rect 3970 18776 3976 18828
rect 4028 18816 4034 18828
rect 4724 18816 4752 18912
rect 4908 18884 4936 18912
rect 9784 18896 9812 18924
rect 10226 18912 10232 18924
rect 10284 18952 10290 18964
rect 10965 18955 11023 18961
rect 10965 18952 10977 18955
rect 10284 18924 10977 18952
rect 10284 18912 10290 18924
rect 10965 18921 10977 18924
rect 11011 18921 11023 18955
rect 10965 18915 11023 18921
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 14550 18952 14556 18964
rect 13504 18924 14556 18952
rect 13504 18912 13510 18924
rect 14550 18912 14556 18924
rect 14608 18912 14614 18964
rect 17589 18955 17647 18961
rect 17589 18921 17601 18955
rect 17635 18952 17647 18955
rect 19610 18952 19616 18964
rect 17635 18924 19616 18952
rect 17635 18921 17647 18924
rect 17589 18915 17647 18921
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 22186 18912 22192 18964
rect 22244 18952 22250 18964
rect 22465 18955 22523 18961
rect 22465 18952 22477 18955
rect 22244 18924 22477 18952
rect 22244 18912 22250 18924
rect 22465 18921 22477 18924
rect 22511 18952 22523 18955
rect 23385 18955 23443 18961
rect 23385 18952 23397 18955
rect 22511 18924 23397 18952
rect 22511 18921 22523 18924
rect 22465 18915 22523 18921
rect 23385 18921 23397 18924
rect 23431 18921 23443 18955
rect 23385 18915 23443 18921
rect 24857 18955 24915 18961
rect 24857 18921 24869 18955
rect 24903 18952 24915 18955
rect 25774 18952 25780 18964
rect 24903 18924 25780 18952
rect 24903 18921 24915 18924
rect 24857 18915 24915 18921
rect 25774 18912 25780 18924
rect 25832 18912 25838 18964
rect 26694 18912 26700 18964
rect 26752 18912 26758 18964
rect 27890 18912 27896 18964
rect 27948 18952 27954 18964
rect 27948 18924 28856 18952
rect 27948 18912 27954 18924
rect 4908 18856 5764 18884
rect 5736 18816 5764 18856
rect 9766 18844 9772 18896
rect 9824 18844 9830 18896
rect 12805 18887 12863 18893
rect 12805 18884 12817 18887
rect 10704 18856 12817 18884
rect 10704 18828 10732 18856
rect 12805 18853 12817 18856
rect 12851 18853 12863 18887
rect 12805 18847 12863 18853
rect 17144 18856 18276 18884
rect 6825 18819 6883 18825
rect 6825 18816 6837 18819
rect 4028 18788 4292 18816
rect 4724 18788 5396 18816
rect 5736 18788 6837 18816
rect 4028 18776 4034 18788
rect 3329 18751 3387 18757
rect 3329 18717 3341 18751
rect 3375 18717 3387 18751
rect 3329 18711 3387 18717
rect 3050 18572 3056 18624
rect 3108 18572 3114 18624
rect 3344 18612 3372 18711
rect 3418 18708 3424 18760
rect 3476 18748 3482 18760
rect 4264 18757 4292 18788
rect 5368 18757 5396 18788
rect 6825 18785 6837 18788
rect 6871 18785 6883 18819
rect 6825 18779 6883 18785
rect 10686 18776 10692 18828
rect 10744 18776 10750 18828
rect 11238 18776 11244 18828
rect 11296 18776 11302 18828
rect 12820 18816 12848 18847
rect 17144 18825 17172 18856
rect 17129 18819 17187 18825
rect 12820 18788 13676 18816
rect 4249 18751 4307 18757
rect 3476 18720 4200 18748
rect 3476 18708 3482 18720
rect 3605 18683 3663 18689
rect 3605 18649 3617 18683
rect 3651 18680 3663 18683
rect 4065 18683 4123 18689
rect 4065 18680 4077 18683
rect 3651 18652 4077 18680
rect 3651 18649 3663 18652
rect 3605 18643 3663 18649
rect 4065 18649 4077 18652
rect 4111 18649 4123 18683
rect 4172 18680 4200 18720
rect 4249 18717 4261 18751
rect 4295 18748 4307 18751
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 4295 18720 5273 18748
rect 4295 18717 4307 18720
rect 4249 18711 4307 18717
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 5353 18751 5411 18757
rect 5353 18717 5365 18751
rect 5399 18717 5411 18751
rect 5353 18711 5411 18717
rect 5276 18680 5304 18711
rect 6546 18708 6552 18760
rect 6604 18708 6610 18760
rect 8294 18708 8300 18760
rect 8352 18748 8358 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 8352 18720 9321 18748
rect 8352 18708 8358 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 10410 18708 10416 18760
rect 10468 18748 10474 18760
rect 10597 18751 10655 18757
rect 10597 18748 10609 18751
rect 10468 18720 10609 18748
rect 10468 18708 10474 18720
rect 10597 18717 10609 18720
rect 10643 18748 10655 18751
rect 11256 18748 11284 18776
rect 10643 18720 11284 18748
rect 11425 18751 11483 18757
rect 10643 18717 10655 18720
rect 10597 18711 10655 18717
rect 11425 18717 11437 18751
rect 11471 18748 11483 18751
rect 11471 18720 11560 18748
rect 11471 18717 11483 18720
rect 11425 18711 11483 18717
rect 4172 18652 5212 18680
rect 5276 18652 5488 18680
rect 4065 18643 4123 18649
rect 5184 18624 5212 18652
rect 5460 18624 5488 18652
rect 7558 18640 7564 18692
rect 7616 18640 7622 18692
rect 9861 18683 9919 18689
rect 9861 18649 9873 18683
rect 9907 18680 9919 18683
rect 10870 18680 10876 18692
rect 9907 18652 10876 18680
rect 9907 18649 9919 18652
rect 9861 18643 9919 18649
rect 10870 18640 10876 18652
rect 10928 18640 10934 18692
rect 4890 18612 4896 18624
rect 3344 18584 4896 18612
rect 4890 18572 4896 18584
rect 4948 18572 4954 18624
rect 5166 18572 5172 18624
rect 5224 18572 5230 18624
rect 5442 18572 5448 18624
rect 5500 18572 5506 18624
rect 8478 18572 8484 18624
rect 8536 18612 8542 18624
rect 8665 18615 8723 18621
rect 8665 18612 8677 18615
rect 8536 18584 8677 18612
rect 8536 18572 8542 18584
rect 8665 18581 8677 18584
rect 8711 18581 8723 18615
rect 8665 18575 8723 18581
rect 9582 18572 9588 18624
rect 9640 18612 9646 18624
rect 10229 18615 10287 18621
rect 10229 18612 10241 18615
rect 9640 18584 10241 18612
rect 9640 18572 9646 18584
rect 10229 18581 10241 18584
rect 10275 18581 10287 18615
rect 10229 18575 10287 18581
rect 11054 18572 11060 18624
rect 11112 18612 11118 18624
rect 11532 18612 11560 18720
rect 11606 18708 11612 18760
rect 11664 18748 11670 18760
rect 13648 18757 13676 18788
rect 17129 18785 17141 18819
rect 17175 18785 17187 18819
rect 17129 18779 17187 18785
rect 17328 18788 17908 18816
rect 17328 18760 17356 18788
rect 12069 18751 12127 18757
rect 12069 18748 12081 18751
rect 11664 18720 12081 18748
rect 11664 18708 11670 18720
rect 12069 18717 12081 18720
rect 12115 18748 12127 18751
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 12115 18720 13277 18748
rect 12115 18717 12127 18720
rect 12069 18711 12127 18717
rect 13265 18717 13277 18720
rect 13311 18748 13323 18751
rect 13541 18751 13599 18757
rect 13541 18748 13553 18751
rect 13311 18720 13553 18748
rect 13311 18717 13323 18720
rect 13265 18711 13323 18717
rect 13541 18717 13553 18720
rect 13587 18717 13599 18751
rect 13541 18711 13599 18717
rect 13633 18751 13691 18757
rect 13633 18717 13645 18751
rect 13679 18717 13691 18751
rect 15102 18748 15108 18760
rect 13633 18711 13691 18717
rect 13740 18720 15108 18748
rect 11701 18683 11759 18689
rect 11701 18649 11713 18683
rect 11747 18680 11759 18683
rect 11790 18680 11796 18692
rect 11747 18652 11796 18680
rect 11747 18649 11759 18652
rect 11701 18643 11759 18649
rect 11790 18640 11796 18652
rect 11848 18640 11854 18692
rect 13357 18683 13415 18689
rect 13357 18680 13369 18683
rect 13280 18652 13369 18680
rect 13280 18624 13308 18652
rect 13357 18649 13369 18652
rect 13403 18649 13415 18683
rect 13556 18680 13584 18711
rect 13740 18680 13768 18720
rect 15102 18708 15108 18720
rect 15160 18708 15166 18760
rect 17218 18708 17224 18760
rect 17276 18708 17282 18760
rect 17310 18708 17316 18760
rect 17368 18708 17374 18760
rect 17880 18757 17908 18788
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17451 18720 17693 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 17865 18751 17923 18757
rect 17865 18717 17877 18751
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18717 18199 18751
rect 18248 18748 18276 18856
rect 18598 18844 18604 18896
rect 18656 18884 18662 18896
rect 18877 18887 18935 18893
rect 18877 18884 18889 18887
rect 18656 18856 18889 18884
rect 18656 18844 18662 18856
rect 18877 18853 18889 18856
rect 18923 18884 18935 18887
rect 18966 18884 18972 18896
rect 18923 18856 18972 18884
rect 18923 18853 18935 18856
rect 18877 18847 18935 18853
rect 18966 18844 18972 18856
rect 19024 18844 19030 18896
rect 21910 18844 21916 18896
rect 21968 18844 21974 18896
rect 22925 18887 22983 18893
rect 22925 18853 22937 18887
rect 22971 18884 22983 18887
rect 23753 18887 23811 18893
rect 22971 18856 23704 18884
rect 22971 18853 22983 18856
rect 22925 18847 22983 18853
rect 18325 18819 18383 18825
rect 18325 18785 18337 18819
rect 18371 18816 18383 18819
rect 19334 18816 19340 18828
rect 18371 18788 19340 18816
rect 18371 18785 18383 18788
rect 18325 18779 18383 18785
rect 19334 18776 19340 18788
rect 19392 18776 19398 18828
rect 22373 18819 22431 18825
rect 22373 18785 22385 18819
rect 22419 18816 22431 18819
rect 22554 18816 22560 18828
rect 22419 18788 22560 18816
rect 22419 18785 22431 18788
rect 22373 18779 22431 18785
rect 22554 18776 22560 18788
rect 22612 18816 22618 18828
rect 23477 18819 23535 18825
rect 23477 18816 23489 18819
rect 22612 18788 23489 18816
rect 22612 18776 22618 18788
rect 23477 18785 23489 18788
rect 23523 18785 23535 18819
rect 23676 18816 23704 18856
rect 23753 18853 23765 18887
rect 23799 18884 23811 18887
rect 27614 18884 27620 18896
rect 23799 18856 27620 18884
rect 23799 18853 23811 18856
rect 23753 18847 23811 18853
rect 27614 18844 27620 18856
rect 27672 18884 27678 18896
rect 28445 18887 28503 18893
rect 28445 18884 28457 18887
rect 27672 18856 28457 18884
rect 27672 18844 27678 18856
rect 28445 18853 28457 18856
rect 28491 18853 28503 18887
rect 28445 18847 28503 18853
rect 25682 18816 25688 18828
rect 23676 18788 25688 18816
rect 23477 18779 23535 18785
rect 25682 18776 25688 18788
rect 25740 18776 25746 18828
rect 25802 18819 25860 18825
rect 25802 18816 25814 18819
rect 25792 18785 25814 18816
rect 25848 18785 25860 18819
rect 25792 18779 25860 18785
rect 18506 18748 18512 18760
rect 18248 18720 18512 18748
rect 18141 18711 18199 18717
rect 13556 18652 13768 18680
rect 13357 18643 13415 18649
rect 13998 18640 14004 18692
rect 14056 18680 14062 18692
rect 16114 18680 16120 18692
rect 14056 18652 16120 18680
rect 14056 18640 14062 18652
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 17420 18680 17448 18711
rect 18156 18680 18184 18711
rect 18506 18708 18512 18720
rect 18564 18748 18570 18760
rect 19058 18748 19064 18760
rect 18564 18720 19064 18748
rect 18564 18708 18570 18720
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18748 20683 18751
rect 20671 18720 20760 18748
rect 20671 18717 20683 18720
rect 20625 18711 20683 18717
rect 20732 18692 20760 18720
rect 20898 18708 20904 18760
rect 20956 18708 20962 18760
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 16224 18652 17448 18680
rect 17512 18652 18184 18680
rect 16224 18624 16252 18652
rect 12437 18615 12495 18621
rect 12437 18612 12449 18615
rect 11112 18584 12449 18612
rect 11112 18572 11118 18584
rect 12437 18581 12449 18584
rect 12483 18612 12495 18615
rect 13170 18612 13176 18624
rect 12483 18584 13176 18612
rect 12483 18581 12495 18584
rect 12437 18575 12495 18581
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 13262 18572 13268 18624
rect 13320 18572 13326 18624
rect 16206 18572 16212 18624
rect 16264 18572 16270 18624
rect 17218 18572 17224 18624
rect 17276 18612 17282 18624
rect 17512 18612 17540 18652
rect 20714 18640 20720 18692
rect 20772 18680 20778 18692
rect 21082 18680 21088 18692
rect 20772 18652 21088 18680
rect 20772 18640 20778 18652
rect 21082 18640 21088 18652
rect 21140 18640 21146 18692
rect 21284 18680 21312 18711
rect 21358 18708 21364 18760
rect 21416 18748 21422 18760
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 21416 18720 21649 18748
rect 21416 18708 21422 18720
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 21818 18708 21824 18760
rect 21876 18748 21882 18760
rect 22005 18751 22063 18757
rect 22005 18748 22017 18751
rect 21876 18720 22017 18748
rect 21876 18708 21882 18720
rect 22005 18717 22017 18720
rect 22051 18717 22063 18751
rect 22005 18711 22063 18717
rect 22462 18708 22468 18760
rect 22520 18748 22526 18760
rect 22649 18751 22707 18757
rect 22649 18748 22661 18751
rect 22520 18720 22661 18748
rect 22520 18708 22526 18720
rect 22649 18717 22661 18720
rect 22695 18717 22707 18751
rect 22649 18711 22707 18717
rect 22741 18751 22799 18757
rect 22741 18717 22753 18751
rect 22787 18748 22799 18751
rect 23198 18748 23204 18760
rect 22787 18720 23204 18748
rect 22787 18717 22799 18720
rect 22741 18711 22799 18717
rect 21542 18680 21548 18692
rect 21284 18652 21548 18680
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 22664 18680 22692 18711
rect 23198 18708 23204 18720
rect 23256 18757 23262 18760
rect 23256 18751 23314 18757
rect 23256 18717 23268 18751
rect 23302 18748 23314 18751
rect 24397 18751 24455 18757
rect 24397 18748 24409 18751
rect 23302 18720 23349 18748
rect 24136 18720 24409 18748
rect 23302 18717 23314 18720
rect 23256 18711 23314 18717
rect 23256 18708 23262 18711
rect 23109 18683 23167 18689
rect 23109 18680 23121 18683
rect 22664 18652 23121 18680
rect 23109 18649 23121 18652
rect 23155 18649 23167 18683
rect 23109 18643 23167 18649
rect 17276 18584 17540 18612
rect 17276 18572 17282 18584
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24136 18621 24164 18720
rect 24397 18717 24409 18720
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 24486 18708 24492 18760
rect 24544 18708 24550 18760
rect 24670 18708 24676 18760
rect 24728 18748 24734 18760
rect 25317 18751 25375 18757
rect 25317 18748 25329 18751
rect 24728 18720 25329 18748
rect 24728 18708 24734 18720
rect 25240 18621 25268 18720
rect 25317 18717 25329 18720
rect 25363 18717 25375 18751
rect 25792 18748 25820 18779
rect 26142 18776 26148 18828
rect 26200 18816 26206 18828
rect 28828 18825 28856 18924
rect 31938 18844 31944 18896
rect 31996 18884 32002 18896
rect 31996 18856 32628 18884
rect 31996 18844 32002 18856
rect 26973 18819 27031 18825
rect 26973 18816 26985 18819
rect 26200 18788 26985 18816
rect 26200 18776 26206 18788
rect 26053 18751 26111 18757
rect 26053 18748 26065 18751
rect 25792 18720 25912 18748
rect 25317 18711 25375 18717
rect 25884 18692 25912 18720
rect 25976 18720 26065 18748
rect 25866 18640 25872 18692
rect 25924 18640 25930 18692
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 23900 18584 24133 18612
rect 23900 18572 23906 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 24121 18575 24179 18581
rect 25225 18615 25283 18621
rect 25225 18581 25237 18615
rect 25271 18612 25283 18615
rect 25406 18612 25412 18624
rect 25271 18584 25412 18612
rect 25271 18581 25283 18584
rect 25225 18575 25283 18581
rect 25406 18572 25412 18584
rect 25464 18572 25470 18624
rect 25590 18572 25596 18624
rect 25648 18572 25654 18624
rect 25682 18572 25688 18624
rect 25740 18572 25746 18624
rect 25976 18621 26004 18720
rect 26053 18717 26065 18720
rect 26099 18717 26111 18751
rect 26053 18711 26111 18717
rect 26234 18708 26240 18760
rect 26292 18708 26298 18760
rect 26528 18757 26556 18788
rect 26973 18785 26985 18788
rect 27019 18785 27031 18819
rect 26973 18779 27031 18785
rect 27985 18819 28043 18825
rect 27985 18785 27997 18819
rect 28031 18816 28043 18819
rect 28353 18819 28411 18825
rect 28353 18816 28365 18819
rect 28031 18788 28365 18816
rect 28031 18785 28043 18788
rect 27985 18779 28043 18785
rect 28353 18785 28365 18788
rect 28399 18785 28411 18819
rect 28353 18779 28411 18785
rect 28813 18819 28871 18825
rect 28813 18785 28825 18819
rect 28859 18785 28871 18819
rect 28813 18779 28871 18785
rect 31297 18819 31355 18825
rect 31297 18785 31309 18819
rect 31343 18816 31355 18819
rect 31662 18816 31668 18828
rect 31343 18788 31668 18816
rect 31343 18785 31355 18788
rect 31297 18779 31355 18785
rect 31662 18776 31668 18788
rect 31720 18816 31726 18828
rect 32033 18819 32091 18825
rect 31720 18776 31754 18816
rect 32033 18785 32045 18819
rect 32079 18816 32091 18819
rect 32493 18819 32551 18825
rect 32493 18816 32505 18819
rect 32079 18788 32505 18816
rect 32079 18785 32091 18788
rect 32033 18779 32091 18785
rect 32493 18785 32505 18788
rect 32539 18785 32551 18819
rect 32493 18779 32551 18785
rect 26513 18751 26571 18757
rect 26513 18717 26525 18751
rect 26559 18717 26571 18751
rect 26513 18711 26571 18717
rect 26786 18708 26792 18760
rect 26844 18748 26850 18760
rect 27798 18748 27804 18760
rect 26844 18720 27804 18748
rect 26844 18708 26850 18720
rect 27798 18708 27804 18720
rect 27856 18748 27862 18760
rect 27893 18751 27951 18757
rect 27893 18748 27905 18751
rect 27856 18720 27905 18748
rect 27856 18708 27862 18720
rect 27893 18717 27905 18720
rect 27939 18717 27951 18751
rect 27893 18711 27951 18717
rect 29365 18751 29423 18757
rect 29365 18717 29377 18751
rect 29411 18748 29423 18751
rect 29546 18748 29552 18760
rect 29411 18720 29552 18748
rect 29411 18717 29423 18720
rect 29365 18711 29423 18717
rect 29546 18708 29552 18720
rect 29604 18708 29610 18760
rect 31726 18748 31754 18776
rect 32600 18760 32628 18856
rect 32674 18776 32680 18828
rect 32732 18816 32738 18828
rect 32769 18819 32827 18825
rect 32769 18816 32781 18819
rect 32732 18788 32781 18816
rect 32732 18776 32738 18788
rect 32769 18785 32781 18788
rect 32815 18816 32827 18819
rect 33042 18816 33048 18828
rect 32815 18788 33048 18816
rect 32815 18785 32827 18788
rect 32769 18779 32827 18785
rect 33042 18776 33048 18788
rect 33100 18776 33106 18828
rect 31941 18751 31999 18757
rect 31941 18748 31953 18751
rect 31726 18720 31953 18748
rect 31941 18717 31953 18720
rect 31987 18717 31999 18751
rect 31941 18711 31999 18717
rect 32398 18708 32404 18760
rect 32456 18708 32462 18760
rect 32582 18708 32588 18760
rect 32640 18708 32646 18760
rect 34330 18708 34336 18760
rect 34388 18748 34394 18760
rect 34701 18751 34759 18757
rect 34701 18748 34713 18751
rect 34388 18720 34713 18748
rect 34388 18708 34394 18720
rect 34701 18717 34713 18720
rect 34747 18717 34759 18751
rect 34701 18711 34759 18717
rect 29825 18683 29883 18689
rect 29825 18680 29837 18683
rect 29104 18652 29837 18680
rect 25961 18615 26019 18621
rect 25961 18581 25973 18615
rect 26007 18581 26019 18615
rect 25961 18575 26019 18581
rect 28261 18615 28319 18621
rect 28261 18581 28273 18615
rect 28307 18612 28319 18615
rect 29104 18612 29132 18652
rect 29825 18649 29837 18652
rect 29871 18649 29883 18683
rect 29825 18643 29883 18649
rect 30282 18640 30288 18692
rect 30340 18640 30346 18692
rect 33045 18683 33103 18689
rect 33045 18680 33057 18683
rect 32324 18652 33057 18680
rect 32324 18621 32352 18652
rect 33045 18649 33057 18652
rect 33091 18649 33103 18683
rect 34793 18683 34851 18689
rect 34793 18680 34805 18683
rect 34270 18652 34805 18680
rect 33045 18643 33103 18649
rect 34793 18649 34805 18652
rect 34839 18649 34851 18683
rect 34793 18643 34851 18649
rect 28307 18584 29132 18612
rect 32309 18615 32367 18621
rect 28307 18581 28319 18584
rect 28261 18575 28319 18581
rect 32309 18581 32321 18615
rect 32355 18581 32367 18615
rect 32309 18575 32367 18581
rect 34514 18572 34520 18624
rect 34572 18572 34578 18624
rect 1104 18522 35236 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 35236 18522
rect 1104 18448 35236 18470
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 13740 18380 14105 18408
rect 12526 18300 12532 18352
rect 12584 18340 12590 18352
rect 13740 18349 13768 18380
rect 14093 18377 14105 18380
rect 14139 18377 14151 18411
rect 14093 18371 14151 18377
rect 14200 18380 17448 18408
rect 13173 18343 13231 18349
rect 12584 18312 13032 18340
rect 12584 18300 12590 18312
rect 13004 18284 13032 18312
rect 13173 18309 13185 18343
rect 13219 18340 13231 18343
rect 13633 18343 13691 18349
rect 13633 18340 13645 18343
rect 13219 18312 13645 18340
rect 13219 18309 13231 18312
rect 13173 18303 13231 18309
rect 13633 18309 13645 18312
rect 13679 18309 13691 18343
rect 13633 18303 13691 18309
rect 13725 18343 13783 18349
rect 13725 18309 13737 18343
rect 13771 18309 13783 18343
rect 13725 18303 13783 18309
rect 13998 18300 14004 18352
rect 14056 18300 14062 18352
rect 4798 18232 4804 18284
rect 4856 18232 4862 18284
rect 4982 18232 4988 18284
rect 5040 18272 5046 18284
rect 5261 18275 5319 18281
rect 5261 18272 5273 18275
rect 5040 18244 5273 18272
rect 5040 18232 5046 18244
rect 5261 18241 5273 18244
rect 5307 18241 5319 18275
rect 5261 18235 5319 18241
rect 5442 18232 5448 18284
rect 5500 18232 5506 18284
rect 10505 18275 10563 18281
rect 10505 18241 10517 18275
rect 10551 18272 10563 18275
rect 10686 18272 10692 18284
rect 10551 18244 10692 18272
rect 10551 18241 10563 18244
rect 10505 18235 10563 18241
rect 10686 18232 10692 18244
rect 10744 18272 10750 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10744 18244 10977 18272
rect 10744 18232 10750 18244
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 10965 18235 11023 18241
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18241 11299 18275
rect 11241 18235 11299 18241
rect 4893 18207 4951 18213
rect 4893 18173 4905 18207
rect 4939 18204 4951 18207
rect 5353 18207 5411 18213
rect 5353 18204 5365 18207
rect 4939 18176 5365 18204
rect 4939 18173 4951 18176
rect 4893 18167 4951 18173
rect 5353 18173 5365 18176
rect 5399 18173 5411 18207
rect 5353 18167 5411 18173
rect 5169 18139 5227 18145
rect 5169 18105 5181 18139
rect 5215 18136 5227 18139
rect 8294 18136 8300 18148
rect 5215 18108 8300 18136
rect 5215 18105 5227 18108
rect 5169 18099 5227 18105
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18136 8447 18139
rect 8435 18108 8984 18136
rect 8435 18105 8447 18108
rect 8389 18099 8447 18105
rect 8956 18080 8984 18108
rect 10870 18096 10876 18148
rect 10928 18136 10934 18148
rect 11256 18136 11284 18235
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11388 18244 11730 18272
rect 11388 18232 11394 18244
rect 12802 18232 12808 18284
rect 12860 18232 12866 18284
rect 12986 18232 12992 18284
rect 13044 18232 13050 18284
rect 13078 18232 13084 18284
rect 13136 18232 13142 18284
rect 13262 18232 13268 18284
rect 13320 18232 13326 18284
rect 13446 18232 13452 18284
rect 13504 18281 13510 18284
rect 13504 18275 13553 18281
rect 13504 18241 13507 18275
rect 13541 18241 13553 18275
rect 13504 18235 13553 18241
rect 13504 18232 13510 18235
rect 13814 18232 13820 18284
rect 13872 18232 13878 18284
rect 11790 18164 11796 18216
rect 11848 18164 11854 18216
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 12667 18176 13369 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 13357 18173 13369 18176
rect 13403 18204 13415 18207
rect 14200 18204 14228 18380
rect 15657 18343 15715 18349
rect 14292 18312 14688 18340
rect 14292 18284 14320 18312
rect 14274 18232 14280 18284
rect 14332 18232 14338 18284
rect 14660 18281 14688 18312
rect 15657 18309 15669 18343
rect 15703 18340 15715 18343
rect 17310 18340 17316 18352
rect 15703 18312 17316 18340
rect 15703 18309 15715 18312
rect 15657 18303 15715 18309
rect 17310 18300 17316 18312
rect 17368 18300 17374 18352
rect 17420 18284 17448 18380
rect 17586 18368 17592 18420
rect 17644 18408 17650 18420
rect 17865 18411 17923 18417
rect 17865 18408 17877 18411
rect 17644 18380 17877 18408
rect 17644 18368 17650 18380
rect 17865 18377 17877 18380
rect 17911 18377 17923 18411
rect 17865 18371 17923 18377
rect 21637 18411 21695 18417
rect 21637 18377 21649 18411
rect 21683 18408 21695 18411
rect 21726 18408 21732 18420
rect 21683 18380 21732 18408
rect 21683 18377 21695 18380
rect 21637 18371 21695 18377
rect 21726 18368 21732 18380
rect 21784 18368 21790 18420
rect 23382 18368 23388 18420
rect 23440 18408 23446 18420
rect 24213 18411 24271 18417
rect 23440 18380 24072 18408
rect 23440 18368 23446 18380
rect 17681 18343 17739 18349
rect 17681 18309 17693 18343
rect 17727 18340 17739 18343
rect 18233 18343 18291 18349
rect 18233 18340 18245 18343
rect 17727 18312 18245 18340
rect 17727 18309 17739 18312
rect 17681 18303 17739 18309
rect 18233 18309 18245 18312
rect 18279 18309 18291 18343
rect 18233 18303 18291 18309
rect 23474 18300 23480 18352
rect 23532 18340 23538 18352
rect 24044 18349 24072 18380
rect 24213 18377 24225 18411
rect 24259 18408 24271 18411
rect 24486 18408 24492 18420
rect 24259 18380 24492 18408
rect 24259 18377 24271 18380
rect 24213 18371 24271 18377
rect 24486 18368 24492 18380
rect 24544 18368 24550 18420
rect 24578 18368 24584 18420
rect 24636 18408 24642 18420
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 24636 18380 24869 18408
rect 24636 18368 24642 18380
rect 24857 18377 24869 18380
rect 24903 18408 24915 18411
rect 25685 18411 25743 18417
rect 24903 18380 25636 18408
rect 24903 18377 24915 18380
rect 24857 18371 24915 18377
rect 25608 18352 25636 18380
rect 25685 18377 25697 18411
rect 25731 18408 25743 18411
rect 26234 18408 26240 18420
rect 25731 18380 26240 18408
rect 25731 18377 25743 18380
rect 25685 18371 25743 18377
rect 26234 18368 26240 18380
rect 26292 18368 26298 18420
rect 30282 18368 30288 18420
rect 30340 18368 30346 18420
rect 34514 18368 34520 18420
rect 34572 18368 34578 18420
rect 23845 18343 23903 18349
rect 23845 18340 23857 18343
rect 23532 18312 23857 18340
rect 23532 18300 23538 18312
rect 23845 18309 23857 18312
rect 23891 18309 23903 18343
rect 24044 18343 24119 18349
rect 24044 18312 24073 18343
rect 23845 18303 23903 18309
rect 24061 18309 24073 18312
rect 24107 18340 24119 18343
rect 24107 18312 25268 18340
rect 24107 18309 24119 18312
rect 24061 18303 24119 18309
rect 14553 18275 14611 18281
rect 14553 18241 14565 18275
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14645 18275 14703 18281
rect 14645 18241 14657 18275
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 14829 18275 14887 18281
rect 14829 18241 14841 18275
rect 14875 18241 14887 18275
rect 14829 18235 14887 18241
rect 13403 18176 14228 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 14366 18164 14372 18216
rect 14424 18164 14430 18216
rect 12897 18139 12955 18145
rect 10928 18108 12480 18136
rect 10928 18096 10934 18108
rect 12452 18080 12480 18108
rect 12897 18105 12909 18139
rect 12943 18136 12955 18139
rect 13722 18136 13728 18148
rect 12943 18108 13728 18136
rect 12943 18105 12955 18108
rect 12897 18099 12955 18105
rect 13722 18096 13728 18108
rect 13780 18136 13786 18148
rect 14568 18136 14596 18235
rect 13780 18108 14596 18136
rect 13780 18096 13786 18108
rect 8478 18028 8484 18080
rect 8536 18068 8542 18080
rect 8757 18071 8815 18077
rect 8757 18068 8769 18071
rect 8536 18040 8769 18068
rect 8536 18028 8542 18040
rect 8757 18037 8769 18040
rect 8803 18037 8815 18071
rect 8757 18031 8815 18037
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 9125 18071 9183 18077
rect 9125 18068 9137 18071
rect 8996 18040 9137 18068
rect 8996 18028 9002 18040
rect 9125 18037 9137 18040
rect 9171 18037 9183 18071
rect 9125 18031 9183 18037
rect 12434 18028 12440 18080
rect 12492 18028 12498 18080
rect 13078 18028 13084 18080
rect 13136 18068 13142 18080
rect 14277 18071 14335 18077
rect 14277 18068 14289 18071
rect 13136 18040 14289 18068
rect 13136 18028 13142 18040
rect 14277 18037 14289 18040
rect 14323 18068 14335 18071
rect 14844 18068 14872 18235
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 15286 18232 15292 18284
rect 15344 18232 15350 18284
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 15013 18207 15071 18213
rect 15013 18173 15025 18207
rect 15059 18204 15071 18207
rect 15488 18204 15516 18235
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15838 18232 15844 18284
rect 15896 18232 15902 18284
rect 15930 18232 15936 18284
rect 15988 18272 15994 18284
rect 16025 18275 16083 18281
rect 16025 18272 16037 18275
rect 15988 18244 16037 18272
rect 15988 18232 15994 18244
rect 16025 18241 16037 18244
rect 16071 18241 16083 18275
rect 16025 18235 16083 18241
rect 16206 18232 16212 18284
rect 16264 18232 16270 18284
rect 17034 18232 17040 18284
rect 17092 18232 17098 18284
rect 17221 18275 17279 18281
rect 17221 18241 17233 18275
rect 17267 18272 17279 18275
rect 17402 18272 17408 18284
rect 17267 18244 17408 18272
rect 17267 18241 17279 18244
rect 17221 18235 17279 18241
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 17494 18232 17500 18284
rect 17552 18232 17558 18284
rect 17586 18232 17592 18284
rect 17644 18232 17650 18284
rect 17957 18275 18015 18281
rect 17957 18241 17969 18275
rect 18003 18272 18015 18275
rect 18003 18244 18184 18272
rect 18003 18241 18015 18244
rect 17957 18235 18015 18241
rect 16666 18204 16672 18216
rect 15059 18176 16672 18204
rect 15059 18173 15071 18176
rect 15013 18167 15071 18173
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 17129 18207 17187 18213
rect 17129 18173 17141 18207
rect 17175 18204 17187 18207
rect 18049 18207 18107 18213
rect 18049 18204 18061 18207
rect 17175 18176 18061 18204
rect 17175 18173 17187 18176
rect 17129 18167 17187 18173
rect 18049 18173 18061 18176
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 17218 18096 17224 18148
rect 17276 18136 17282 18148
rect 17313 18139 17371 18145
rect 17313 18136 17325 18139
rect 17276 18108 17325 18136
rect 17276 18096 17282 18108
rect 17313 18105 17325 18108
rect 17359 18136 17371 18139
rect 17402 18136 17408 18148
rect 17359 18108 17408 18136
rect 17359 18105 17371 18108
rect 17313 18099 17371 18105
rect 17402 18096 17408 18108
rect 17460 18096 17466 18148
rect 14323 18040 14872 18068
rect 14323 18037 14335 18040
rect 14277 18031 14335 18037
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15930 18068 15936 18080
rect 15436 18040 15936 18068
rect 15436 18028 15442 18040
rect 15930 18028 15936 18040
rect 15988 18028 15994 18080
rect 16482 18028 16488 18080
rect 16540 18068 16546 18080
rect 18156 18068 18184 18244
rect 19702 18232 19708 18284
rect 19760 18232 19766 18284
rect 20346 18232 20352 18284
rect 20404 18232 20410 18284
rect 21358 18232 21364 18284
rect 21416 18232 21422 18284
rect 21453 18275 21511 18281
rect 21453 18241 21465 18275
rect 21499 18272 21511 18275
rect 21818 18272 21824 18284
rect 21499 18244 21824 18272
rect 21499 18241 21511 18244
rect 21453 18235 21511 18241
rect 21818 18232 21824 18244
rect 21876 18232 21882 18284
rect 18233 18207 18291 18213
rect 18233 18173 18245 18207
rect 18279 18204 18291 18207
rect 18506 18204 18512 18216
rect 18279 18176 18512 18204
rect 18279 18173 18291 18176
rect 18233 18167 18291 18173
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 23860 18204 23888 18303
rect 24302 18232 24308 18284
rect 24360 18232 24366 18284
rect 24489 18276 24547 18281
rect 24412 18275 24547 18276
rect 24412 18248 24501 18275
rect 24412 18204 24440 18248
rect 24489 18241 24501 18248
rect 24535 18241 24547 18275
rect 24489 18235 24547 18241
rect 25240 18216 25268 18312
rect 25590 18300 25596 18352
rect 25648 18300 25654 18352
rect 25777 18343 25835 18349
rect 25777 18309 25789 18343
rect 25823 18340 25835 18343
rect 25958 18340 25964 18352
rect 25823 18312 25964 18340
rect 25823 18309 25835 18312
rect 25777 18303 25835 18309
rect 25682 18232 25688 18284
rect 25740 18272 25746 18284
rect 25792 18272 25820 18303
rect 25958 18300 25964 18312
rect 26016 18300 26022 18352
rect 25740 18244 25820 18272
rect 25740 18232 25746 18244
rect 23860 18176 24440 18204
rect 25222 18164 25228 18216
rect 25280 18164 25286 18216
rect 25406 18164 25412 18216
rect 25464 18164 25470 18216
rect 20714 18096 20720 18148
rect 20772 18096 20778 18148
rect 23750 18096 23756 18148
rect 23808 18136 23814 18148
rect 25130 18136 25136 18148
rect 23808 18108 25136 18136
rect 23808 18096 23814 18108
rect 24044 18077 24072 18108
rect 25130 18096 25136 18108
rect 25188 18136 25194 18148
rect 25792 18136 25820 18244
rect 25866 18232 25872 18284
rect 25924 18232 25930 18284
rect 30190 18272 30196 18284
rect 30024 18244 30196 18272
rect 25188 18108 25820 18136
rect 25188 18096 25194 18108
rect 16540 18040 18184 18068
rect 24029 18071 24087 18077
rect 16540 18028 16546 18040
rect 24029 18037 24041 18071
rect 24075 18068 24087 18071
rect 24075 18040 24109 18068
rect 24075 18037 24087 18040
rect 24029 18031 24087 18037
rect 24394 18028 24400 18080
rect 24452 18028 24458 18080
rect 25222 18028 25228 18080
rect 25280 18068 25286 18080
rect 25884 18068 25912 18232
rect 30024 18080 30052 18244
rect 30190 18232 30196 18244
rect 30248 18232 30254 18284
rect 34532 18272 34560 18368
rect 34701 18275 34759 18281
rect 34701 18272 34713 18275
rect 34532 18244 34713 18272
rect 34701 18241 34713 18244
rect 34747 18241 34759 18275
rect 34701 18235 34759 18241
rect 34790 18232 34796 18284
rect 34848 18232 34854 18284
rect 34425 18207 34483 18213
rect 34425 18173 34437 18207
rect 34471 18204 34483 18207
rect 34808 18204 34836 18232
rect 34471 18176 34836 18204
rect 34471 18173 34483 18176
rect 34425 18167 34483 18173
rect 26050 18068 26056 18080
rect 25280 18040 26056 18068
rect 25280 18028 25286 18040
rect 26050 18028 26056 18040
rect 26108 18068 26114 18080
rect 26145 18071 26203 18077
rect 26145 18068 26157 18071
rect 26108 18040 26157 18068
rect 26108 18028 26114 18040
rect 26145 18037 26157 18040
rect 26191 18037 26203 18071
rect 26145 18031 26203 18037
rect 30006 18028 30012 18080
rect 30064 18028 30070 18080
rect 32677 18071 32735 18077
rect 32677 18037 32689 18071
rect 32723 18068 32735 18071
rect 33042 18068 33048 18080
rect 32723 18040 33048 18068
rect 32723 18037 32735 18040
rect 32677 18031 32735 18037
rect 33042 18028 33048 18040
rect 33100 18028 33106 18080
rect 1104 17978 35248 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 35248 17978
rect 1104 17904 35248 17926
rect 5166 17824 5172 17876
rect 5224 17824 5230 17876
rect 6546 17824 6552 17876
rect 6604 17824 6610 17876
rect 8294 17824 8300 17876
rect 8352 17824 8358 17876
rect 13633 17867 13691 17873
rect 13633 17833 13645 17867
rect 13679 17864 13691 17867
rect 13814 17864 13820 17876
rect 13679 17836 13820 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 14185 17867 14243 17873
rect 14185 17833 14197 17867
rect 14231 17864 14243 17867
rect 14274 17864 14280 17876
rect 14231 17836 14280 17864
rect 14231 17833 14243 17836
rect 14185 17827 14243 17833
rect 1670 17688 1676 17740
rect 1728 17688 1734 17740
rect 5258 17728 5264 17740
rect 5000 17700 5264 17728
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 1412 17592 1440 17623
rect 1412 17564 1532 17592
rect 1504 17524 1532 17564
rect 2314 17552 2320 17604
rect 2372 17552 2378 17604
rect 3050 17592 3056 17604
rect 2976 17564 3056 17592
rect 2976 17524 3004 17564
rect 3050 17552 3056 17564
rect 3108 17592 3114 17604
rect 3108 17564 3464 17592
rect 3108 17552 3114 17564
rect 3436 17536 3464 17564
rect 4890 17552 4896 17604
rect 4948 17592 4954 17604
rect 5000 17601 5028 17700
rect 5258 17688 5264 17700
rect 5316 17688 5322 17740
rect 6362 17688 6368 17740
rect 6420 17728 6426 17740
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 6420 17700 6469 17728
rect 6420 17688 6426 17700
rect 6457 17697 6469 17700
rect 6503 17728 6515 17731
rect 6564 17728 6592 17824
rect 6503 17700 6592 17728
rect 8312 17728 8340 17824
rect 13722 17756 13728 17808
rect 13780 17756 13786 17808
rect 9217 17731 9275 17737
rect 9217 17728 9229 17731
rect 8312 17700 9229 17728
rect 6503 17697 6515 17700
rect 6457 17691 6515 17697
rect 9217 17697 9229 17700
rect 9263 17697 9275 17731
rect 9217 17691 9275 17697
rect 11330 17688 11336 17740
rect 11388 17728 11394 17740
rect 11425 17731 11483 17737
rect 11425 17728 11437 17731
rect 11388 17700 11437 17728
rect 11388 17688 11394 17700
rect 11425 17697 11437 17700
rect 11471 17697 11483 17731
rect 11425 17691 11483 17697
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 13740 17728 13768 17756
rect 14200 17728 14228 17827
rect 14274 17824 14280 17836
rect 14332 17824 14338 17876
rect 14642 17824 14648 17876
rect 14700 17824 14706 17876
rect 15194 17824 15200 17876
rect 15252 17824 15258 17876
rect 15286 17824 15292 17876
rect 15344 17864 15350 17876
rect 15381 17867 15439 17873
rect 15381 17864 15393 17867
rect 15344 17836 15393 17864
rect 15344 17824 15350 17836
rect 15381 17833 15393 17836
rect 15427 17833 15439 17867
rect 15381 17827 15439 17833
rect 15838 17824 15844 17876
rect 15896 17864 15902 17876
rect 16482 17864 16488 17876
rect 15896 17836 16488 17864
rect 15896 17824 15902 17836
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 16761 17867 16819 17873
rect 16761 17833 16773 17867
rect 16807 17833 16819 17867
rect 16761 17827 16819 17833
rect 17129 17867 17187 17873
rect 17129 17833 17141 17867
rect 17175 17864 17187 17867
rect 17494 17864 17500 17876
rect 17175 17836 17500 17864
rect 17175 17833 17187 17836
rect 17129 17827 17187 17833
rect 13587 17700 13768 17728
rect 13832 17700 14228 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 8481 17663 8539 17669
rect 8481 17629 8493 17663
rect 8527 17629 8539 17663
rect 8481 17623 8539 17629
rect 4985 17595 5043 17601
rect 4985 17592 4997 17595
rect 4948 17564 4997 17592
rect 4948 17552 4954 17564
rect 4985 17561 4997 17564
rect 5031 17561 5043 17595
rect 4985 17555 5043 17561
rect 6730 17552 6736 17604
rect 6788 17552 6794 17604
rect 8389 17595 8447 17601
rect 8389 17592 8401 17595
rect 7958 17564 8401 17592
rect 8389 17561 8401 17564
rect 8435 17561 8447 17595
rect 8389 17555 8447 17561
rect 8496 17536 8524 17623
rect 8938 17620 8944 17672
rect 8996 17620 9002 17672
rect 11701 17663 11759 17669
rect 11701 17629 11713 17663
rect 11747 17660 11759 17663
rect 11790 17660 11796 17672
rect 11747 17632 11796 17660
rect 11747 17629 11759 17632
rect 11701 17623 11759 17629
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 13832 17669 13860 17700
rect 13725 17663 13783 17669
rect 13725 17660 13737 17663
rect 13320 17632 13737 17660
rect 13320 17620 13326 17632
rect 13725 17629 13737 17632
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 13817 17663 13875 17669
rect 13817 17629 13829 17663
rect 13863 17629 13875 17663
rect 13817 17623 13875 17629
rect 8956 17592 8984 17620
rect 8956 17564 9628 17592
rect 9600 17536 9628 17564
rect 9950 17552 9956 17604
rect 10008 17552 10014 17604
rect 10965 17595 11023 17601
rect 10965 17592 10977 17595
rect 10520 17564 10977 17592
rect 1504 17496 3004 17524
rect 3142 17484 3148 17536
rect 3200 17484 3206 17536
rect 3418 17484 3424 17536
rect 3476 17484 3482 17536
rect 4154 17484 4160 17536
rect 4212 17524 4218 17536
rect 5185 17527 5243 17533
rect 5185 17524 5197 17527
rect 4212 17496 5197 17524
rect 4212 17484 4218 17496
rect 5185 17493 5197 17496
rect 5231 17493 5243 17527
rect 5185 17487 5243 17493
rect 5350 17484 5356 17536
rect 5408 17484 5414 17536
rect 8202 17484 8208 17536
rect 8260 17484 8266 17536
rect 8478 17484 8484 17536
rect 8536 17484 8542 17536
rect 9582 17484 9588 17536
rect 9640 17524 9646 17536
rect 10520 17524 10548 17564
rect 10965 17561 10977 17564
rect 11011 17561 11023 17595
rect 13740 17592 13768 17623
rect 13998 17620 14004 17672
rect 14056 17620 14062 17672
rect 14090 17620 14096 17672
rect 14148 17620 14154 17672
rect 14274 17620 14280 17672
rect 14332 17660 14338 17672
rect 14660 17660 14688 17824
rect 15930 17756 15936 17808
rect 15988 17796 15994 17808
rect 16776 17796 16804 17827
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 20625 17867 20683 17873
rect 20625 17833 20637 17867
rect 20671 17864 20683 17867
rect 21358 17864 21364 17876
rect 20671 17836 21364 17864
rect 20671 17833 20683 17836
rect 20625 17827 20683 17833
rect 21358 17824 21364 17836
rect 21416 17824 21422 17876
rect 22922 17824 22928 17876
rect 22980 17864 22986 17876
rect 23201 17867 23259 17873
rect 23201 17864 23213 17867
rect 22980 17836 23213 17864
rect 22980 17824 22986 17836
rect 23201 17833 23213 17836
rect 23247 17864 23259 17867
rect 23290 17864 23296 17876
rect 23247 17836 23296 17864
rect 23247 17833 23259 17836
rect 23201 17827 23259 17833
rect 23290 17824 23296 17836
rect 23348 17824 23354 17876
rect 23474 17824 23480 17876
rect 23532 17864 23538 17876
rect 23753 17867 23811 17873
rect 23753 17864 23765 17867
rect 23532 17836 23765 17864
rect 23532 17824 23538 17836
rect 23753 17833 23765 17836
rect 23799 17864 23811 17867
rect 24213 17867 24271 17873
rect 24213 17864 24225 17867
rect 23799 17836 24225 17864
rect 23799 17833 23811 17836
rect 23753 17827 23811 17833
rect 24213 17833 24225 17836
rect 24259 17833 24271 17867
rect 24213 17827 24271 17833
rect 25130 17824 25136 17876
rect 25188 17864 25194 17876
rect 25869 17867 25927 17873
rect 25869 17864 25881 17867
rect 25188 17836 25881 17864
rect 25188 17824 25194 17836
rect 25869 17833 25881 17836
rect 25915 17864 25927 17867
rect 25958 17864 25964 17876
rect 25915 17836 25964 17864
rect 25915 17833 25927 17836
rect 25869 17827 25927 17833
rect 25958 17824 25964 17836
rect 26016 17824 26022 17876
rect 26326 17824 26332 17876
rect 26384 17864 26390 17876
rect 26602 17864 26608 17876
rect 26384 17836 26608 17864
rect 26384 17824 26390 17836
rect 26602 17824 26608 17836
rect 26660 17824 26666 17876
rect 15988 17768 16804 17796
rect 15988 17756 15994 17768
rect 20990 17756 20996 17808
rect 21048 17756 21054 17808
rect 14936 17700 16068 17728
rect 14936 17669 14964 17700
rect 14921 17663 14979 17669
rect 14921 17660 14933 17663
rect 14332 17632 14688 17660
rect 14752 17632 14933 17660
rect 14332 17620 14338 17632
rect 14016 17592 14044 17620
rect 14366 17592 14372 17604
rect 13740 17564 14372 17592
rect 10965 17555 11023 17561
rect 14366 17552 14372 17564
rect 14424 17552 14430 17604
rect 14752 17536 14780 17632
rect 14921 17629 14933 17632
rect 14967 17629 14979 17663
rect 14921 17623 14979 17629
rect 15289 17663 15347 17669
rect 15289 17629 15301 17663
rect 15335 17660 15347 17663
rect 15470 17660 15476 17672
rect 15335 17632 15476 17660
rect 15335 17629 15347 17632
rect 15289 17623 15347 17629
rect 15470 17620 15476 17632
rect 15528 17620 15534 17672
rect 15580 17669 15608 17700
rect 15565 17663 15623 17669
rect 15565 17629 15577 17663
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 15657 17663 15715 17669
rect 15657 17629 15669 17663
rect 15703 17629 15715 17663
rect 15841 17663 15899 17669
rect 15841 17660 15853 17663
rect 15657 17623 15715 17629
rect 15764 17632 15853 17660
rect 15672 17592 15700 17623
rect 15028 17564 15700 17592
rect 15028 17536 15056 17564
rect 9640 17496 10548 17524
rect 10689 17527 10747 17533
rect 9640 17484 9646 17496
rect 10689 17493 10701 17527
rect 10735 17524 10747 17527
rect 11238 17524 11244 17536
rect 10735 17496 11244 17524
rect 10735 17493 10747 17496
rect 10689 17487 10747 17493
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 12342 17484 12348 17536
rect 12400 17484 12406 17536
rect 12713 17527 12771 17533
rect 12713 17493 12725 17527
rect 12759 17524 12771 17527
rect 12986 17524 12992 17536
rect 12759 17496 12992 17524
rect 12759 17493 12771 17496
rect 12713 17487 12771 17493
rect 12986 17484 12992 17496
rect 13044 17484 13050 17536
rect 13170 17484 13176 17536
rect 13228 17524 13234 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 13228 17496 13461 17524
rect 13228 17484 13234 17496
rect 13449 17493 13461 17496
rect 13495 17524 13507 17527
rect 14090 17524 14096 17536
rect 13495 17496 14096 17524
rect 13495 17493 13507 17496
rect 13449 17487 13507 17493
rect 14090 17484 14096 17496
rect 14148 17484 14154 17536
rect 14734 17484 14740 17536
rect 14792 17484 14798 17536
rect 15010 17484 15016 17536
rect 15068 17484 15074 17536
rect 15105 17527 15163 17533
rect 15105 17493 15117 17527
rect 15151 17524 15163 17527
rect 15378 17524 15384 17536
rect 15151 17496 15384 17524
rect 15151 17493 15163 17496
rect 15105 17487 15163 17493
rect 15378 17484 15384 17496
rect 15436 17484 15442 17536
rect 15470 17484 15476 17536
rect 15528 17524 15534 17536
rect 15764 17524 15792 17632
rect 15841 17629 15853 17632
rect 15887 17629 15899 17663
rect 15841 17623 15899 17629
rect 15930 17620 15936 17672
rect 15988 17620 15994 17672
rect 16040 17669 16068 17700
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17678 17728 17684 17740
rect 16724 17700 17684 17728
rect 16724 17688 16730 17700
rect 17678 17688 17684 17700
rect 17736 17728 17742 17740
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 17736 17700 18153 17728
rect 17736 17688 17742 17700
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 18141 17691 18199 17697
rect 19061 17731 19119 17737
rect 19061 17697 19073 17731
rect 19107 17728 19119 17731
rect 19702 17728 19708 17740
rect 19107 17700 19708 17728
rect 19107 17697 19119 17700
rect 19061 17691 19119 17697
rect 19702 17688 19708 17700
rect 19760 17688 19766 17740
rect 20346 17688 20352 17740
rect 20404 17688 20410 17740
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 16301 17663 16359 17669
rect 16301 17629 16313 17663
rect 16347 17660 16359 17663
rect 16574 17660 16580 17672
rect 16347 17632 16580 17660
rect 16347 17629 16359 17632
rect 16301 17623 16359 17629
rect 16114 17552 16120 17604
rect 16172 17552 16178 17604
rect 16316 17524 16344 17623
rect 16574 17620 16580 17632
rect 16632 17620 16638 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17660 16819 17663
rect 16807 17632 16896 17660
rect 16807 17629 16819 17632
rect 16761 17623 16819 17629
rect 16868 17536 16896 17632
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 18325 17663 18383 17669
rect 18325 17629 18337 17663
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 15528 17496 16344 17524
rect 15528 17484 15534 17496
rect 16850 17484 16856 17536
rect 16908 17484 16914 17536
rect 17034 17484 17040 17536
rect 17092 17524 17098 17536
rect 17770 17524 17776 17536
rect 17092 17496 17776 17524
rect 17092 17484 17098 17496
rect 17770 17484 17776 17496
rect 17828 17524 17834 17536
rect 18340 17524 18368 17623
rect 19334 17620 19340 17672
rect 19392 17620 19398 17672
rect 19426 17620 19432 17672
rect 19484 17660 19490 17672
rect 19521 17663 19579 17669
rect 19521 17660 19533 17663
rect 19484 17632 19533 17660
rect 19484 17620 19490 17632
rect 19521 17629 19533 17632
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 20533 17663 20591 17669
rect 20533 17629 20545 17663
rect 20579 17660 20591 17663
rect 20717 17663 20775 17669
rect 20579 17632 20668 17660
rect 20579 17629 20591 17632
rect 20533 17623 20591 17629
rect 20640 17536 20668 17632
rect 20717 17629 20729 17663
rect 20763 17660 20775 17663
rect 21008 17660 21036 17756
rect 25590 17688 25596 17740
rect 25648 17728 25654 17740
rect 26510 17728 26516 17740
rect 25648 17700 26516 17728
rect 25648 17688 25654 17700
rect 26510 17688 26516 17700
rect 26568 17688 26574 17740
rect 20763 17632 21036 17660
rect 20763 17629 20775 17632
rect 20717 17623 20775 17629
rect 24762 17620 24768 17672
rect 24820 17660 24826 17672
rect 26786 17660 26792 17672
rect 24820 17632 26792 17660
rect 24820 17620 24826 17632
rect 26786 17620 26792 17632
rect 26844 17620 26850 17672
rect 17828 17496 18368 17524
rect 17828 17484 17834 17496
rect 20622 17484 20628 17536
rect 20680 17484 20686 17536
rect 22922 17484 22928 17536
rect 22980 17484 22986 17536
rect 25130 17484 25136 17536
rect 25188 17524 25194 17536
rect 25406 17524 25412 17536
rect 25188 17496 25412 17524
rect 25188 17484 25194 17496
rect 25406 17484 25412 17496
rect 25464 17524 25470 17536
rect 25501 17527 25559 17533
rect 25501 17524 25513 17527
rect 25464 17496 25513 17524
rect 25464 17484 25470 17496
rect 25501 17493 25513 17496
rect 25547 17493 25559 17527
rect 25501 17487 25559 17493
rect 26050 17484 26056 17536
rect 26108 17524 26114 17536
rect 26237 17527 26295 17533
rect 26237 17524 26249 17527
rect 26108 17496 26249 17524
rect 26108 17484 26114 17496
rect 26237 17493 26249 17496
rect 26283 17493 26295 17527
rect 26237 17487 26295 17493
rect 1104 17434 35236 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 35236 17434
rect 1104 17360 35236 17382
rect 2314 17280 2320 17332
rect 2372 17280 2378 17332
rect 3142 17280 3148 17332
rect 3200 17280 3206 17332
rect 4341 17323 4399 17329
rect 4341 17289 4353 17323
rect 4387 17320 4399 17323
rect 4982 17320 4988 17332
rect 4387 17292 4988 17320
rect 4387 17289 4399 17292
rect 4341 17283 4399 17289
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 5350 17280 5356 17332
rect 5408 17280 5414 17332
rect 6730 17280 6736 17332
rect 6788 17280 6794 17332
rect 8202 17280 8208 17332
rect 8260 17320 8266 17332
rect 8260 17292 8800 17320
rect 8260 17280 8266 17292
rect 934 17144 940 17196
rect 992 17184 998 17196
rect 1397 17187 1455 17193
rect 1397 17184 1409 17187
rect 992 17156 1409 17184
rect 992 17144 998 17156
rect 1397 17153 1409 17156
rect 1443 17153 1455 17187
rect 1397 17147 1455 17153
rect 2225 17187 2283 17193
rect 2225 17153 2237 17187
rect 2271 17184 2283 17187
rect 2866 17184 2872 17196
rect 2271 17156 2872 17184
rect 2271 17153 2283 17156
rect 2225 17147 2283 17153
rect 2866 17144 2872 17156
rect 2924 17184 2930 17196
rect 3160 17184 3188 17280
rect 3421 17187 3479 17193
rect 3421 17184 3433 17187
rect 2924 17156 3004 17184
rect 3160 17156 3433 17184
rect 2924 17144 2930 17156
rect 2866 17048 2872 17060
rect 1596 17020 2872 17048
rect 1596 16989 1624 17020
rect 2866 17008 2872 17020
rect 2924 17008 2930 17060
rect 1581 16983 1639 16989
rect 1581 16949 1593 16983
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 2976 16980 3004 17156
rect 3421 17153 3433 17156
rect 3467 17184 3479 17187
rect 3881 17187 3939 17193
rect 3881 17184 3893 17187
rect 3467 17156 3893 17184
rect 3467 17153 3479 17156
rect 3421 17147 3479 17153
rect 3881 17153 3893 17156
rect 3927 17153 3939 17187
rect 4154 17184 4160 17196
rect 3881 17147 3939 17153
rect 3988 17156 4160 17184
rect 3988 17128 4016 17156
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 5261 17187 5319 17193
rect 5261 17184 5273 17187
rect 4672 17156 5273 17184
rect 4672 17144 4678 17156
rect 5261 17153 5273 17156
rect 5307 17153 5319 17187
rect 5261 17147 5319 17153
rect 3510 17076 3516 17128
rect 3568 17076 3574 17128
rect 3970 17076 3976 17128
rect 4028 17076 4034 17128
rect 4062 17076 4068 17128
rect 4120 17076 4126 17128
rect 5368 17125 5396 17280
rect 6748 17252 6776 17280
rect 5644 17224 6776 17252
rect 5644 17125 5672 17224
rect 7374 17212 7380 17264
rect 7432 17212 7438 17264
rect 8772 17261 8800 17292
rect 9950 17280 9956 17332
rect 10008 17280 10014 17332
rect 12342 17280 12348 17332
rect 12400 17320 12406 17332
rect 12400 17280 12434 17320
rect 15746 17280 15752 17332
rect 15804 17320 15810 17332
rect 15933 17323 15991 17329
rect 15933 17320 15945 17323
rect 15804 17292 15945 17320
rect 15804 17280 15810 17292
rect 15933 17289 15945 17292
rect 15979 17289 15991 17323
rect 15933 17283 15991 17289
rect 16022 17280 16028 17332
rect 16080 17320 16086 17332
rect 16666 17320 16672 17332
rect 16080 17292 16672 17320
rect 16080 17280 16086 17292
rect 16666 17280 16672 17292
rect 16724 17320 16730 17332
rect 16942 17320 16948 17332
rect 16724 17292 16948 17320
rect 16724 17280 16730 17292
rect 16942 17280 16948 17292
rect 17000 17280 17006 17332
rect 17586 17280 17592 17332
rect 17644 17280 17650 17332
rect 20990 17280 20996 17332
rect 21048 17280 21054 17332
rect 21818 17280 21824 17332
rect 21876 17280 21882 17332
rect 22922 17280 22928 17332
rect 22980 17320 22986 17332
rect 24026 17320 24032 17332
rect 22980 17292 24032 17320
rect 22980 17280 22986 17292
rect 8757 17255 8815 17261
rect 8757 17221 8769 17255
rect 8803 17221 8815 17255
rect 8757 17215 8815 17221
rect 9398 17212 9404 17264
rect 9456 17252 9462 17264
rect 10962 17252 10968 17264
rect 9456 17224 10968 17252
rect 9456 17212 9462 17224
rect 10962 17212 10968 17224
rect 11020 17212 11026 17264
rect 11238 17212 11244 17264
rect 11296 17212 11302 17264
rect 11333 17255 11391 17261
rect 11333 17221 11345 17255
rect 11379 17252 11391 17255
rect 12406 17252 12434 17280
rect 15838 17252 15844 17264
rect 11379 17224 12296 17252
rect 12406 17224 15844 17252
rect 11379 17221 11391 17224
rect 11333 17215 11391 17221
rect 6362 17144 6368 17196
rect 6420 17144 6426 17196
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 8128 17156 8217 17184
rect 8128 17125 8156 17156
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17184 8539 17187
rect 9416 17184 9444 17212
rect 8527 17156 9444 17184
rect 9861 17187 9919 17193
rect 8527 17153 8539 17156
rect 8481 17147 8539 17153
rect 9861 17153 9873 17187
rect 9907 17184 9919 17187
rect 10321 17187 10379 17193
rect 10321 17184 10333 17187
rect 9907 17156 10333 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 10321 17153 10333 17156
rect 10367 17153 10379 17187
rect 10321 17147 10379 17153
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 11057 17187 11115 17193
rect 11057 17184 11069 17187
rect 10827 17156 11069 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 11057 17153 11069 17156
rect 11103 17153 11115 17187
rect 11057 17147 11115 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11256 17184 11284 17212
rect 11609 17187 11667 17193
rect 11609 17184 11621 17187
rect 11195 17156 11621 17184
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 11609 17153 11621 17156
rect 11655 17153 11667 17187
rect 12268 17184 12296 17224
rect 13078 17184 13084 17196
rect 12268 17156 13084 17184
rect 11609 17147 11667 17153
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17085 5411 17119
rect 5353 17079 5411 17085
rect 5629 17119 5687 17125
rect 5629 17085 5641 17119
rect 5675 17085 5687 17119
rect 6641 17119 6699 17125
rect 6641 17116 6653 17119
rect 5629 17079 5687 17085
rect 6472 17088 6653 17116
rect 3789 17051 3847 17057
rect 3789 17017 3801 17051
rect 3835 17048 3847 17051
rect 6472 17048 6500 17088
rect 6641 17085 6653 17088
rect 6687 17085 6699 17119
rect 6641 17079 6699 17085
rect 8113 17119 8171 17125
rect 8113 17085 8125 17119
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17116 9551 17119
rect 9766 17116 9772 17128
rect 9539 17088 9772 17116
rect 9539 17085 9551 17088
rect 9493 17079 9551 17085
rect 9766 17076 9772 17088
rect 9824 17076 9830 17128
rect 3835 17020 6500 17048
rect 3835 17017 3847 17020
rect 3789 17011 3847 17017
rect 8018 17008 8024 17060
rect 8076 17048 8082 17060
rect 8478 17048 8484 17060
rect 8076 17020 8484 17048
rect 8076 17008 8082 17020
rect 8478 17008 8484 17020
rect 8536 17048 8542 17060
rect 9876 17048 9904 17147
rect 11072 17116 11100 17147
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 13630 17144 13636 17196
rect 13688 17144 13694 17196
rect 13998 17144 14004 17196
rect 14056 17144 14062 17196
rect 14277 17190 14335 17193
rect 14108 17187 14335 17190
rect 14108 17162 14289 17187
rect 11974 17116 11980 17128
rect 11072 17088 11980 17116
rect 11974 17076 11980 17088
rect 12032 17076 12038 17128
rect 12161 17119 12219 17125
rect 12161 17085 12173 17119
rect 12207 17116 12219 17119
rect 12618 17116 12624 17128
rect 12207 17088 12624 17116
rect 12207 17085 12219 17088
rect 12161 17079 12219 17085
rect 12618 17076 12624 17088
rect 12676 17076 12682 17128
rect 13096 17116 13124 17144
rect 14108 17116 14136 17162
rect 14277 17153 14289 17162
rect 14323 17184 14335 17187
rect 14458 17184 14464 17196
rect 14323 17156 14464 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14458 17144 14464 17156
rect 14516 17144 14522 17196
rect 14645 17187 14703 17193
rect 14645 17153 14657 17187
rect 14691 17153 14703 17187
rect 14645 17147 14703 17153
rect 13096 17088 14136 17116
rect 8536 17020 9904 17048
rect 8536 17008 8542 17020
rect 12986 17008 12992 17060
rect 13044 17048 13050 17060
rect 13044 17020 13308 17048
rect 13044 17008 13050 17020
rect 3602 16980 3608 16992
rect 2823 16952 3608 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4614 16980 4620 16992
rect 4203 16952 4620 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4614 16940 4620 16952
rect 4672 16940 4678 16992
rect 13280 16989 13308 17020
rect 13265 16983 13323 16989
rect 13265 16949 13277 16983
rect 13311 16980 13323 16983
rect 14366 16980 14372 16992
rect 13311 16952 14372 16980
rect 13311 16949 13323 16952
rect 13265 16943 13323 16949
rect 14366 16940 14372 16952
rect 14424 16980 14430 16992
rect 14660 16980 14688 17147
rect 14844 17116 14872 17224
rect 15838 17212 15844 17224
rect 15896 17252 15902 17264
rect 15896 17224 17264 17252
rect 15896 17212 15902 17224
rect 14918 17144 14924 17196
rect 14976 17144 14982 17196
rect 15010 17144 15016 17196
rect 15068 17184 15074 17196
rect 15197 17187 15255 17193
rect 15197 17184 15209 17187
rect 15068 17156 15209 17184
rect 15068 17144 15074 17156
rect 15197 17153 15209 17156
rect 15243 17184 15255 17187
rect 15565 17187 15623 17193
rect 15565 17184 15577 17187
rect 15243 17156 15577 17184
rect 15243 17153 15255 17156
rect 15197 17147 15255 17153
rect 15565 17153 15577 17156
rect 15611 17184 15623 17187
rect 16025 17187 16083 17193
rect 16025 17184 16037 17187
rect 15611 17156 16037 17184
rect 15611 17153 15623 17156
rect 15565 17147 15623 17153
rect 16025 17153 16037 17156
rect 16071 17184 16083 17187
rect 16114 17184 16120 17196
rect 16071 17156 16120 17184
rect 16071 17153 16083 17156
rect 16025 17147 16083 17153
rect 16114 17144 16120 17156
rect 16172 17144 16178 17196
rect 16209 17187 16267 17193
rect 16209 17153 16221 17187
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 15473 17119 15531 17125
rect 15473 17116 15485 17119
rect 14844 17088 15485 17116
rect 15473 17085 15485 17088
rect 15519 17085 15531 17119
rect 15473 17079 15531 17085
rect 15657 17119 15715 17125
rect 15657 17085 15669 17119
rect 15703 17085 15715 17119
rect 15657 17079 15715 17085
rect 14734 17008 14740 17060
rect 14792 17048 14798 17060
rect 15672 17048 15700 17079
rect 15746 17076 15752 17128
rect 15804 17076 15810 17128
rect 16224 17048 16252 17147
rect 16758 17144 16764 17196
rect 16816 17144 16822 17196
rect 16942 17144 16948 17196
rect 17000 17144 17006 17196
rect 17236 17193 17264 17224
rect 17402 17212 17408 17264
rect 17460 17212 17466 17264
rect 21008 17252 21036 17280
rect 20824 17224 21036 17252
rect 22373 17255 22431 17261
rect 17221 17187 17279 17193
rect 17221 17153 17233 17187
rect 17267 17153 17279 17187
rect 17221 17147 17279 17153
rect 17310 17144 17316 17196
rect 17368 17184 17374 17196
rect 17770 17184 17776 17196
rect 17368 17156 17776 17184
rect 17368 17144 17374 17156
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 18138 17144 18144 17196
rect 18196 17184 18202 17196
rect 19426 17184 19432 17196
rect 18196 17156 19432 17184
rect 18196 17144 18202 17156
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 20824 17193 20852 17224
rect 22373 17221 22385 17255
rect 22419 17252 22431 17255
rect 22419 17224 22968 17252
rect 22419 17221 22431 17224
rect 22373 17215 22431 17221
rect 22940 17196 22968 17224
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 22097 17187 22155 17193
rect 22097 17184 22109 17187
rect 20809 17147 20867 17153
rect 20916 17156 22109 17184
rect 16393 17119 16451 17125
rect 16393 17085 16405 17119
rect 16439 17116 16451 17119
rect 16850 17116 16856 17128
rect 16439 17088 16856 17116
rect 16439 17085 16451 17088
rect 16393 17079 16451 17085
rect 16850 17076 16856 17088
rect 16908 17116 16914 17128
rect 17497 17119 17555 17125
rect 17497 17116 17509 17119
rect 16908 17088 17509 17116
rect 16908 17076 16914 17088
rect 17497 17085 17509 17088
rect 17543 17116 17555 17119
rect 18233 17119 18291 17125
rect 18233 17116 18245 17119
rect 17543 17088 18245 17116
rect 17543 17085 17555 17088
rect 17497 17079 17555 17085
rect 18233 17085 18245 17088
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 20622 17076 20628 17128
rect 20680 17116 20686 17128
rect 20717 17119 20775 17125
rect 20717 17116 20729 17119
rect 20680 17088 20729 17116
rect 20680 17076 20686 17088
rect 20717 17085 20729 17088
rect 20763 17116 20775 17119
rect 20916 17116 20944 17156
rect 22097 17153 22109 17156
rect 22143 17153 22155 17187
rect 22097 17147 22155 17153
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 22741 17187 22799 17193
rect 22741 17153 22753 17187
rect 22787 17153 22799 17187
rect 22741 17147 22799 17153
rect 20763 17088 20944 17116
rect 20763 17085 20775 17088
rect 20717 17079 20775 17085
rect 20990 17076 20996 17128
rect 21048 17076 21054 17128
rect 21634 17076 21640 17128
rect 21692 17076 21698 17128
rect 22005 17119 22063 17125
rect 22005 17085 22017 17119
rect 22051 17085 22063 17119
rect 22005 17079 22063 17085
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17116 22523 17119
rect 22756 17116 22784 17147
rect 22922 17144 22928 17196
rect 22980 17144 22986 17196
rect 23216 17193 23244 17292
rect 24026 17280 24032 17292
rect 24084 17280 24090 17332
rect 24394 17280 24400 17332
rect 24452 17320 24458 17332
rect 24452 17292 24624 17320
rect 24452 17280 24458 17292
rect 23293 17255 23351 17261
rect 23293 17221 23305 17255
rect 23339 17252 23351 17255
rect 23339 17224 24532 17252
rect 23339 17221 23351 17224
rect 23293 17215 23351 17221
rect 23201 17187 23259 17193
rect 23201 17153 23213 17187
rect 23247 17153 23259 17187
rect 23201 17147 23259 17153
rect 23385 17187 23443 17193
rect 23385 17153 23397 17187
rect 23431 17184 23443 17187
rect 23431 17156 23612 17184
rect 23431 17153 23443 17156
rect 23385 17147 23443 17153
rect 23477 17119 23535 17125
rect 23477 17116 23489 17119
rect 22511 17088 23489 17116
rect 22511 17085 22523 17088
rect 22465 17079 22523 17085
rect 23477 17085 23489 17088
rect 23523 17085 23535 17119
rect 23477 17079 23535 17085
rect 14792 17020 16252 17048
rect 21008 17048 21036 17076
rect 22020 17048 22048 17079
rect 21008 17020 22048 17048
rect 14792 17008 14798 17020
rect 23290 17008 23296 17060
rect 23348 17048 23354 17060
rect 23584 17048 23612 17156
rect 23658 17144 23664 17196
rect 23716 17144 23722 17196
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 23845 17187 23903 17193
rect 23845 17153 23857 17187
rect 23891 17153 23903 17187
rect 23845 17147 23903 17153
rect 23860 17048 23888 17147
rect 23934 17144 23940 17196
rect 23992 17193 23998 17196
rect 23992 17187 24041 17193
rect 23992 17153 23995 17187
rect 24029 17184 24041 17187
rect 24029 17156 24440 17184
rect 24029 17153 24041 17156
rect 23992 17147 24041 17153
rect 23992 17144 23998 17147
rect 24121 17119 24179 17125
rect 24121 17085 24133 17119
rect 24167 17085 24179 17119
rect 24121 17079 24179 17085
rect 23348 17020 23888 17048
rect 23348 17008 23354 17020
rect 24136 16992 24164 17079
rect 24412 17048 24440 17156
rect 24504 17125 24532 17224
rect 24596 17193 24624 17292
rect 25240 17292 26924 17320
rect 25240 17261 25268 17292
rect 25225 17255 25283 17261
rect 25225 17221 25237 17255
rect 25271 17221 25283 17255
rect 26237 17255 26295 17261
rect 26237 17252 26249 17255
rect 25225 17215 25283 17221
rect 25976 17224 26249 17252
rect 24581 17187 24639 17193
rect 24581 17153 24593 17187
rect 24627 17153 24639 17187
rect 24581 17147 24639 17153
rect 24489 17119 24547 17125
rect 24489 17085 24501 17119
rect 24535 17085 24547 17119
rect 25240 17116 25268 17215
rect 25872 17196 25924 17202
rect 25976 17193 26004 17224
rect 26237 17221 26249 17224
rect 26283 17221 26295 17255
rect 26237 17215 26295 17221
rect 26418 17212 26424 17264
rect 26476 17252 26482 17264
rect 26694 17252 26700 17264
rect 26476 17224 26700 17252
rect 26476 17212 26482 17224
rect 26694 17212 26700 17224
rect 26752 17212 26758 17264
rect 26896 17252 26924 17292
rect 26896 17224 27292 17252
rect 25961 17187 26019 17193
rect 25961 17153 25973 17187
rect 26007 17153 26019 17187
rect 25961 17147 26019 17153
rect 26145 17187 26203 17193
rect 26145 17153 26157 17187
rect 26191 17153 26203 17187
rect 26145 17147 26203 17153
rect 25872 17138 25924 17144
rect 24489 17079 24547 17085
rect 24596 17088 25268 17116
rect 24596 17048 24624 17088
rect 26050 17076 26056 17128
rect 26108 17116 26114 17128
rect 26160 17116 26188 17147
rect 26326 17144 26332 17196
rect 26384 17144 26390 17196
rect 26513 17187 26571 17193
rect 26513 17153 26525 17187
rect 26559 17153 26571 17187
rect 26513 17147 26571 17153
rect 26789 17187 26847 17193
rect 26789 17153 26801 17187
rect 26835 17185 26847 17187
rect 26896 17185 26924 17224
rect 27264 17193 27292 17224
rect 26835 17157 26924 17185
rect 26973 17187 27031 17193
rect 26835 17153 26847 17157
rect 26789 17147 26847 17153
rect 26973 17153 26985 17187
rect 27019 17153 27031 17187
rect 26973 17147 27031 17153
rect 27065 17187 27123 17193
rect 27065 17153 27077 17187
rect 27111 17153 27123 17187
rect 27065 17147 27123 17153
rect 27249 17187 27307 17193
rect 27249 17153 27261 17187
rect 27295 17153 27307 17187
rect 27249 17147 27307 17153
rect 26108 17088 26188 17116
rect 26528 17116 26556 17147
rect 26988 17116 27016 17147
rect 26528 17088 27016 17116
rect 26108 17076 26114 17088
rect 26528 17048 26556 17088
rect 24412 17020 24624 17048
rect 24872 17020 26556 17048
rect 24872 16992 24900 17020
rect 26694 17008 26700 17060
rect 26752 17048 26758 17060
rect 27080 17048 27108 17147
rect 26752 17020 27108 17048
rect 26752 17008 26758 17020
rect 15102 16980 15108 16992
rect 14424 16952 15108 16980
rect 14424 16940 14430 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 17402 16940 17408 16992
rect 17460 16980 17466 16992
rect 17678 16980 17684 16992
rect 17460 16952 17684 16980
rect 17460 16940 17466 16952
rect 17678 16940 17684 16952
rect 17736 16980 17742 16992
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17736 16952 17785 16980
rect 17736 16940 17742 16952
rect 17773 16949 17785 16952
rect 17819 16949 17831 16983
rect 17773 16943 17831 16949
rect 24118 16940 24124 16992
rect 24176 16980 24182 16992
rect 24213 16983 24271 16989
rect 24213 16980 24225 16983
rect 24176 16952 24225 16980
rect 24176 16940 24182 16952
rect 24213 16949 24225 16952
rect 24259 16949 24271 16983
rect 24213 16943 24271 16949
rect 24854 16940 24860 16992
rect 24912 16940 24918 16992
rect 26786 16940 26792 16992
rect 26844 16940 26850 16992
rect 27246 16940 27252 16992
rect 27304 16980 27310 16992
rect 27433 16983 27491 16989
rect 27433 16980 27445 16983
rect 27304 16952 27445 16980
rect 27304 16940 27310 16952
rect 27433 16949 27445 16952
rect 27479 16949 27491 16983
rect 27433 16943 27491 16949
rect 1104 16890 35248 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 35248 16890
rect 1104 16816 35248 16838
rect 3510 16736 3516 16788
rect 3568 16776 3574 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3568 16748 3801 16776
rect 3568 16736 3574 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 7374 16736 7380 16788
rect 7432 16776 7438 16788
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 7432 16748 7481 16776
rect 7432 16736 7438 16748
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7469 16739 7527 16745
rect 11238 16736 11244 16788
rect 11296 16736 11302 16788
rect 11517 16779 11575 16785
rect 11517 16745 11529 16779
rect 11563 16745 11575 16779
rect 11517 16739 11575 16745
rect 4062 16668 4068 16720
rect 4120 16708 4126 16720
rect 4157 16711 4215 16717
rect 4157 16708 4169 16711
rect 4120 16680 4169 16708
rect 4120 16668 4126 16680
rect 4157 16677 4169 16680
rect 4203 16677 4215 16711
rect 4157 16671 4215 16677
rect 10686 16668 10692 16720
rect 10744 16668 10750 16720
rect 11149 16711 11207 16717
rect 11149 16677 11161 16711
rect 11195 16708 11207 16711
rect 11256 16708 11284 16736
rect 11195 16680 11284 16708
rect 11195 16677 11207 16680
rect 11149 16671 11207 16677
rect 4080 16612 4660 16640
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4080 16581 4108 16612
rect 4632 16584 4660 16612
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 10704 16640 10732 16668
rect 11532 16652 11560 16739
rect 11974 16736 11980 16788
rect 12032 16736 12038 16788
rect 14458 16736 14464 16788
rect 14516 16736 14522 16788
rect 14734 16736 14740 16788
rect 14792 16736 14798 16788
rect 16758 16736 16764 16788
rect 16816 16736 16822 16788
rect 16942 16736 16948 16788
rect 17000 16736 17006 16788
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 18414 16776 18420 16788
rect 18104 16748 18420 16776
rect 18104 16736 18110 16748
rect 18414 16736 18420 16748
rect 18472 16736 18478 16788
rect 19426 16736 19432 16788
rect 19484 16736 19490 16788
rect 22922 16736 22928 16788
rect 22980 16776 22986 16788
rect 23753 16779 23811 16785
rect 23753 16776 23765 16779
rect 22980 16748 23765 16776
rect 22980 16736 22986 16748
rect 23753 16745 23765 16748
rect 23799 16745 23811 16779
rect 23753 16739 23811 16745
rect 24854 16736 24860 16788
rect 24912 16736 24918 16788
rect 25866 16736 25872 16788
rect 25924 16776 25930 16788
rect 26053 16779 26111 16785
rect 26053 16776 26065 16779
rect 25924 16748 26065 16776
rect 25924 16736 25930 16748
rect 26053 16745 26065 16748
rect 26099 16745 26111 16779
rect 26053 16739 26111 16745
rect 26234 16736 26240 16788
rect 26292 16776 26298 16788
rect 27801 16779 27859 16785
rect 27801 16776 27813 16779
rect 26292 16748 27813 16776
rect 26292 16736 26298 16748
rect 27801 16745 27813 16748
rect 27847 16745 27859 16779
rect 27801 16739 27859 16745
rect 11514 16640 11520 16652
rect 9640 16612 9720 16640
rect 10704 16612 11520 16640
rect 9640 16600 9646 16612
rect 4065 16575 4123 16581
rect 4065 16541 4077 16575
rect 4111 16541 4123 16575
rect 4065 16535 4123 16541
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4264 16504 4292 16535
rect 4614 16532 4620 16584
rect 4672 16532 4678 16584
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 7377 16575 7435 16581
rect 7377 16541 7389 16575
rect 7423 16572 7435 16575
rect 7423 16544 7972 16572
rect 7423 16541 7435 16544
rect 7377 16535 7435 16541
rect 5000 16504 5028 16532
rect 4264 16476 5028 16504
rect 7944 16445 7972 16544
rect 7929 16439 7987 16445
rect 7929 16405 7941 16439
rect 7975 16436 7987 16439
rect 8018 16436 8024 16448
rect 7975 16408 8024 16436
rect 7975 16405 7987 16408
rect 7929 16399 7987 16405
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 8478 16436 8484 16448
rect 8343 16408 8484 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 8478 16396 8484 16408
rect 8536 16436 8542 16448
rect 9692 16436 9720 16612
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 13538 16600 13544 16652
rect 13596 16640 13602 16652
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 13596 16612 13921 16640
rect 13596 16600 13602 16612
rect 13909 16609 13921 16612
rect 13955 16640 13967 16643
rect 13955 16612 14412 16640
rect 13955 16609 13967 16612
rect 13909 16603 13967 16609
rect 14384 16584 14412 16612
rect 13630 16532 13636 16584
rect 13688 16572 13694 16584
rect 14093 16575 14151 16581
rect 14093 16572 14105 16575
rect 13688 16544 14105 16572
rect 13688 16532 13694 16544
rect 14093 16541 14105 16544
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 14185 16575 14243 16581
rect 14185 16541 14197 16575
rect 14231 16541 14243 16575
rect 14185 16535 14243 16541
rect 11057 16507 11115 16513
rect 11057 16473 11069 16507
rect 11103 16504 11115 16507
rect 11517 16507 11575 16513
rect 11517 16504 11529 16507
rect 11103 16476 11529 16504
rect 11103 16473 11115 16476
rect 11057 16467 11115 16473
rect 11517 16473 11529 16476
rect 11563 16504 11575 16507
rect 12986 16504 12992 16516
rect 11563 16476 12992 16504
rect 11563 16473 11575 16476
rect 11517 16467 11575 16473
rect 12986 16464 12992 16476
rect 13044 16464 13050 16516
rect 13998 16464 14004 16516
rect 14056 16504 14062 16516
rect 14200 16504 14228 16535
rect 14366 16532 14372 16584
rect 14424 16532 14430 16584
rect 14476 16572 14504 16736
rect 16776 16708 16804 16736
rect 17037 16711 17095 16717
rect 17037 16708 17049 16711
rect 16776 16680 17049 16708
rect 17037 16677 17049 16680
rect 17083 16677 17095 16711
rect 17037 16671 17095 16677
rect 23290 16668 23296 16720
rect 23348 16708 23354 16720
rect 24673 16711 24731 16717
rect 24673 16708 24685 16711
rect 23348 16680 24685 16708
rect 23348 16668 23354 16680
rect 24673 16677 24685 16680
rect 24719 16677 24731 16711
rect 24673 16671 24731 16677
rect 16574 16600 16580 16652
rect 16632 16640 16638 16652
rect 16632 16612 17724 16640
rect 16632 16600 16638 16612
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14476 16544 14565 16572
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16761 16575 16819 16581
rect 16761 16572 16773 16575
rect 16724 16544 16773 16572
rect 16724 16532 16730 16544
rect 16761 16541 16773 16544
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16572 17279 16575
rect 17402 16572 17408 16584
rect 17267 16544 17408 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 14056 16476 14228 16504
rect 14056 16464 14062 16476
rect 9861 16439 9919 16445
rect 9861 16436 9873 16439
rect 8536 16408 9873 16436
rect 8536 16396 8542 16408
rect 9861 16405 9873 16408
rect 9907 16405 9919 16439
rect 9861 16399 9919 16405
rect 10321 16439 10379 16445
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10502 16436 10508 16448
rect 10367 16408 10508 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 10502 16396 10508 16408
rect 10560 16396 10566 16448
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11790 16436 11796 16448
rect 11747 16408 11796 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11790 16396 11796 16408
rect 11848 16396 11854 16448
rect 12434 16396 12440 16448
rect 12492 16436 12498 16448
rect 13170 16436 13176 16448
rect 12492 16408 13176 16436
rect 12492 16396 12498 16408
rect 13170 16396 13176 16408
rect 13228 16396 13234 16448
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 14090 16436 14096 16448
rect 13403 16408 14096 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 14200 16436 14228 16476
rect 14461 16507 14519 16513
rect 14461 16473 14473 16507
rect 14507 16504 14519 16507
rect 14734 16504 14740 16516
rect 14507 16476 14740 16504
rect 14507 16473 14519 16476
rect 14461 16467 14519 16473
rect 14734 16464 14740 16476
rect 14792 16504 14798 16516
rect 14918 16504 14924 16516
rect 14792 16476 14924 16504
rect 14792 16464 14798 16476
rect 14918 16464 14924 16476
rect 14976 16464 14982 16516
rect 16776 16504 16804 16535
rect 17402 16532 17408 16544
rect 17460 16532 17466 16584
rect 17696 16581 17724 16612
rect 21634 16600 21640 16652
rect 21692 16640 21698 16652
rect 22097 16643 22155 16649
rect 22097 16640 22109 16643
rect 21692 16612 22109 16640
rect 21692 16600 21698 16612
rect 22097 16609 22109 16612
rect 22143 16609 22155 16643
rect 22097 16603 22155 16609
rect 23385 16643 23443 16649
rect 23385 16609 23397 16643
rect 23431 16640 23443 16643
rect 23750 16640 23756 16652
rect 23431 16612 23756 16640
rect 23431 16609 23443 16612
rect 23385 16603 23443 16609
rect 17497 16575 17555 16581
rect 17497 16541 17509 16575
rect 17543 16541 17555 16575
rect 17497 16535 17555 16541
rect 17681 16575 17739 16581
rect 17681 16541 17693 16575
rect 17727 16572 17739 16575
rect 18138 16572 18144 16584
rect 17727 16544 18144 16572
rect 17727 16541 17739 16544
rect 17681 16535 17739 16541
rect 17512 16504 17540 16535
rect 18138 16532 18144 16544
rect 18196 16532 18202 16584
rect 19242 16532 19248 16584
rect 19300 16532 19306 16584
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16572 22431 16575
rect 22554 16572 22560 16584
rect 22419 16544 22560 16572
rect 22419 16541 22431 16544
rect 22373 16535 22431 16541
rect 22554 16532 22560 16544
rect 22612 16532 22618 16584
rect 16776 16476 17540 16504
rect 17788 16476 18644 16504
rect 17788 16448 17816 16476
rect 14366 16436 14372 16448
rect 14200 16408 14372 16436
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 17770 16396 17776 16448
rect 17828 16396 17834 16448
rect 18616 16436 18644 16476
rect 18690 16464 18696 16516
rect 18748 16504 18754 16516
rect 23400 16504 23428 16603
rect 23750 16600 23756 16612
rect 23808 16600 23814 16652
rect 24688 16640 24716 16671
rect 25958 16668 25964 16720
rect 26016 16708 26022 16720
rect 26697 16711 26755 16717
rect 26697 16708 26709 16711
rect 26016 16680 26709 16708
rect 26016 16668 26022 16680
rect 26697 16677 26709 16680
rect 26743 16708 26755 16711
rect 27433 16711 27491 16717
rect 27433 16708 27445 16711
rect 26743 16680 27445 16708
rect 26743 16677 26755 16680
rect 26697 16671 26755 16677
rect 27433 16677 27445 16680
rect 27479 16677 27491 16711
rect 27433 16671 27491 16677
rect 26050 16640 26056 16652
rect 24688 16612 25268 16640
rect 25240 16584 25268 16612
rect 25884 16612 26056 16640
rect 23934 16532 23940 16584
rect 23992 16532 23998 16584
rect 24118 16532 24124 16584
rect 24176 16532 24182 16584
rect 24394 16532 24400 16584
rect 24452 16572 24458 16584
rect 25041 16575 25099 16581
rect 25041 16572 25053 16575
rect 24452 16544 25053 16572
rect 24452 16532 24458 16544
rect 25041 16541 25053 16544
rect 25087 16541 25099 16575
rect 25041 16535 25099 16541
rect 25130 16532 25136 16584
rect 25188 16532 25194 16584
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 25884 16581 25912 16612
rect 26050 16600 26056 16612
rect 26108 16600 26114 16652
rect 27065 16643 27123 16649
rect 27065 16640 27077 16643
rect 26160 16612 27077 16640
rect 25317 16575 25375 16581
rect 25317 16541 25329 16575
rect 25363 16572 25375 16575
rect 25409 16575 25467 16581
rect 25409 16572 25421 16575
rect 25363 16544 25421 16572
rect 25363 16541 25375 16544
rect 25317 16535 25375 16541
rect 25409 16541 25421 16544
rect 25455 16541 25467 16575
rect 25409 16535 25467 16541
rect 25593 16575 25651 16581
rect 25593 16541 25605 16575
rect 25639 16541 25651 16575
rect 25869 16575 25927 16581
rect 25869 16572 25881 16575
rect 25593 16535 25651 16541
rect 25700 16544 25881 16572
rect 18748 16476 23428 16504
rect 18748 16464 18754 16476
rect 24026 16464 24032 16516
rect 24084 16504 24090 16516
rect 25148 16504 25176 16532
rect 25608 16504 25636 16535
rect 24084 16476 25636 16504
rect 24084 16464 24090 16476
rect 19426 16436 19432 16448
rect 18616 16408 19432 16436
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 23017 16439 23075 16445
rect 23017 16405 23029 16439
rect 23063 16436 23075 16439
rect 23566 16436 23572 16448
rect 23063 16408 23572 16436
rect 23063 16405 23075 16408
rect 23017 16399 23075 16405
rect 23566 16396 23572 16408
rect 23624 16396 23630 16448
rect 25406 16396 25412 16448
rect 25464 16436 25470 16448
rect 25700 16436 25728 16544
rect 25869 16541 25881 16544
rect 25915 16541 25927 16575
rect 25869 16535 25927 16541
rect 25958 16532 25964 16584
rect 26016 16532 26022 16584
rect 26160 16581 26188 16612
rect 27065 16609 27077 16612
rect 27111 16609 27123 16643
rect 30006 16640 30012 16652
rect 27065 16603 27123 16609
rect 29748 16612 30012 16640
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 26160 16504 26188 16535
rect 26234 16532 26240 16584
rect 26292 16532 26298 16584
rect 29748 16581 29776 16612
rect 30006 16600 30012 16612
rect 30064 16600 30070 16652
rect 26421 16575 26479 16581
rect 26421 16541 26433 16575
rect 26467 16572 26479 16575
rect 29733 16575 29791 16581
rect 26467 16544 26556 16572
rect 26467 16541 26479 16544
rect 26421 16535 26479 16541
rect 25976 16476 26188 16504
rect 25976 16448 26004 16476
rect 26528 16448 26556 16544
rect 29733 16541 29745 16575
rect 29779 16541 29791 16575
rect 29733 16535 29791 16541
rect 34517 16575 34575 16581
rect 34517 16541 34529 16575
rect 34563 16572 34575 16575
rect 34563 16544 35296 16572
rect 34563 16541 34575 16544
rect 34517 16535 34575 16541
rect 33597 16507 33655 16513
rect 33597 16473 33609 16507
rect 33643 16504 33655 16507
rect 34606 16504 34612 16516
rect 33643 16476 34612 16504
rect 33643 16473 33655 16476
rect 33597 16467 33655 16473
rect 34606 16464 34612 16476
rect 34664 16464 34670 16516
rect 25464 16408 25728 16436
rect 25777 16439 25835 16445
rect 25464 16396 25470 16408
rect 25777 16405 25789 16439
rect 25823 16436 25835 16439
rect 25866 16436 25872 16448
rect 25823 16408 25872 16436
rect 25823 16405 25835 16408
rect 25777 16399 25835 16405
rect 25866 16396 25872 16408
rect 25924 16396 25930 16448
rect 25958 16396 25964 16448
rect 26016 16396 26022 16448
rect 26234 16396 26240 16448
rect 26292 16396 26298 16448
rect 26510 16396 26516 16448
rect 26568 16396 26574 16448
rect 29638 16396 29644 16448
rect 29696 16396 29702 16448
rect 1104 16346 35236 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 35236 16346
rect 1104 16272 35236 16294
rect 10597 16235 10655 16241
rect 10597 16201 10609 16235
rect 10643 16232 10655 16235
rect 11054 16232 11060 16244
rect 10643 16204 11060 16232
rect 10643 16201 10655 16204
rect 10597 16195 10655 16201
rect 11054 16192 11060 16204
rect 11112 16192 11118 16244
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11379 16204 12664 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 3970 16124 3976 16176
rect 4028 16164 4034 16176
rect 4028 16136 5396 16164
rect 4028 16124 4034 16136
rect 3326 16056 3332 16108
rect 3384 16096 3390 16108
rect 4062 16096 4068 16108
rect 3384 16068 4068 16096
rect 3384 16056 3390 16068
rect 4062 16056 4068 16068
rect 4120 16096 4126 16108
rect 4433 16099 4491 16105
rect 4433 16096 4445 16099
rect 4120 16068 4445 16096
rect 4120 16056 4126 16068
rect 4433 16065 4445 16068
rect 4479 16065 4491 16099
rect 4433 16059 4491 16065
rect 4982 16056 4988 16108
rect 5040 16096 5046 16108
rect 5368 16105 5396 16136
rect 5442 16124 5448 16176
rect 5500 16164 5506 16176
rect 8481 16167 8539 16173
rect 8481 16164 8493 16167
rect 5500 16136 8493 16164
rect 5500 16124 5506 16136
rect 8481 16133 8493 16136
rect 8527 16133 8539 16167
rect 10137 16167 10195 16173
rect 10137 16164 10149 16167
rect 9706 16136 10149 16164
rect 8481 16127 8539 16133
rect 10137 16133 10149 16136
rect 10183 16133 10195 16167
rect 10137 16127 10195 16133
rect 5077 16099 5135 16105
rect 5077 16096 5089 16099
rect 5040 16068 5089 16096
rect 5040 16056 5046 16068
rect 5077 16065 5089 16068
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 5353 16099 5411 16105
rect 5353 16065 5365 16099
rect 5399 16065 5411 16099
rect 5353 16059 5411 16065
rect 4525 16031 4583 16037
rect 4525 15997 4537 16031
rect 4571 16028 4583 16031
rect 4893 16031 4951 16037
rect 4893 16028 4905 16031
rect 4571 16000 4905 16028
rect 4571 15997 4583 16000
rect 4525 15991 4583 15997
rect 4893 15997 4905 16000
rect 4939 15997 4951 16031
rect 5092 16028 5120 16059
rect 5460 16028 5488 16124
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16065 10287 16099
rect 11072 16096 11100 16192
rect 12529 16167 12587 16173
rect 12529 16164 12541 16167
rect 11900 16136 12541 16164
rect 11900 16105 11928 16136
rect 12529 16133 12541 16136
rect 12575 16133 12587 16167
rect 12529 16127 12587 16133
rect 12636 16108 12664 16204
rect 13630 16192 13636 16244
rect 13688 16232 13694 16244
rect 13725 16235 13783 16241
rect 13725 16232 13737 16235
rect 13688 16204 13737 16232
rect 13688 16192 13694 16204
rect 13725 16201 13737 16204
rect 13771 16232 13783 16235
rect 14642 16232 14648 16244
rect 13771 16204 14648 16232
rect 13771 16201 13783 16204
rect 13725 16195 13783 16201
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 15289 16235 15347 16241
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15746 16232 15752 16244
rect 15335 16204 15752 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 17313 16235 17371 16241
rect 17313 16201 17325 16235
rect 17359 16232 17371 16235
rect 18322 16232 18328 16244
rect 17359 16204 18328 16232
rect 17359 16201 17371 16204
rect 17313 16195 17371 16201
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18509 16235 18567 16241
rect 18509 16201 18521 16235
rect 18555 16232 18567 16235
rect 18598 16232 18604 16244
rect 18555 16204 18604 16232
rect 18555 16201 18567 16204
rect 18509 16195 18567 16201
rect 18598 16192 18604 16204
rect 18656 16192 18662 16244
rect 18966 16232 18972 16244
rect 18800 16204 18972 16232
rect 13541 16167 13599 16173
rect 13541 16133 13553 16167
rect 13587 16164 13599 16167
rect 14660 16164 14688 16192
rect 18800 16164 18828 16204
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 19153 16235 19211 16241
rect 19153 16201 19165 16235
rect 19199 16232 19211 16235
rect 19242 16232 19248 16244
rect 19199 16204 19248 16232
rect 19199 16201 19211 16204
rect 19153 16195 19211 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19334 16192 19340 16244
rect 19392 16192 19398 16244
rect 19426 16192 19432 16244
rect 19484 16192 19490 16244
rect 19889 16235 19947 16241
rect 19889 16201 19901 16235
rect 19935 16232 19947 16235
rect 20622 16232 20628 16244
rect 19935 16204 20628 16232
rect 19935 16201 19947 16204
rect 19889 16195 19947 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 23382 16232 23388 16244
rect 21008 16204 23388 16232
rect 19352 16164 19380 16192
rect 13587 16136 14136 16164
rect 14660 16136 15240 16164
rect 13587 16133 13599 16136
rect 13541 16127 13599 16133
rect 11701 16099 11759 16105
rect 11072 16094 11652 16096
rect 11701 16094 11713 16099
rect 11072 16068 11713 16094
rect 11624 16066 11713 16068
rect 10229 16059 10287 16065
rect 11701 16065 11713 16066
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16096 12311 16099
rect 12434 16096 12440 16108
rect 12299 16068 12440 16096
rect 12299 16065 12311 16068
rect 12253 16059 12311 16065
rect 5092 16000 5488 16028
rect 8205 16031 8263 16037
rect 4893 15991 4951 15997
rect 8205 15997 8217 16031
rect 8251 16028 8263 16031
rect 8478 16028 8484 16040
rect 8251 16000 8484 16028
rect 8251 15997 8263 16000
rect 8205 15991 8263 15997
rect 8478 15988 8484 16000
rect 8536 15988 8542 16040
rect 10244 16028 10272 16059
rect 10502 16028 10508 16040
rect 10244 16000 10508 16028
rect 10502 15988 10508 16000
rect 10560 15988 10566 16040
rect 11790 15988 11796 16040
rect 11848 16028 11854 16040
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 11848 16000 11989 16028
rect 11848 15988 11854 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 11977 15991 12035 15997
rect 12066 15988 12072 16040
rect 12124 15988 12130 16040
rect 4614 15920 4620 15972
rect 4672 15960 4678 15972
rect 5261 15963 5319 15969
rect 5261 15960 5273 15963
rect 4672 15932 5273 15960
rect 4672 15920 4678 15932
rect 5261 15929 5273 15932
rect 5307 15929 5319 15963
rect 5261 15923 5319 15929
rect 10965 15963 11023 15969
rect 10965 15929 10977 15963
rect 11011 15960 11023 15963
rect 12268 15960 12296 16059
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 12618 16056 12624 16108
rect 12676 16096 12682 16108
rect 12805 16099 12863 16105
rect 12805 16096 12817 16099
rect 12676 16068 12817 16096
rect 12676 16056 12682 16068
rect 12805 16065 12817 16068
rect 12851 16096 12863 16099
rect 13262 16096 13268 16108
rect 12851 16068 13268 16096
rect 12851 16065 12863 16068
rect 12805 16059 12863 16065
rect 13262 16056 13268 16068
rect 13320 16056 13326 16108
rect 12713 16031 12771 16037
rect 12713 16028 12725 16031
rect 11011 15932 12296 15960
rect 12360 16000 12725 16028
rect 11011 15929 11023 15932
rect 10965 15923 11023 15929
rect 4798 15852 4804 15904
rect 4856 15852 4862 15904
rect 9950 15852 9956 15904
rect 10008 15852 10014 15904
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12360 15892 12388 16000
rect 12713 15997 12725 16000
rect 12759 15997 12771 16031
rect 12713 15991 12771 15997
rect 13170 15988 13176 16040
rect 13228 16028 13234 16040
rect 13832 16028 13860 16136
rect 13909 16099 13967 16105
rect 13909 16065 13921 16099
rect 13955 16096 13967 16099
rect 13998 16096 14004 16108
rect 13955 16068 14004 16096
rect 13955 16065 13967 16068
rect 13909 16059 13967 16065
rect 13998 16056 14004 16068
rect 14056 16056 14062 16108
rect 14108 16105 14136 16136
rect 15212 16108 15240 16136
rect 15304 16136 18828 16164
rect 18892 16136 19380 16164
rect 19444 16164 19472 16192
rect 19521 16167 19579 16173
rect 19521 16164 19533 16167
rect 19444 16136 19533 16164
rect 14093 16099 14151 16105
rect 14093 16065 14105 16099
rect 14139 16096 14151 16099
rect 14274 16096 14280 16108
rect 14139 16068 14280 16096
rect 14139 16065 14151 16068
rect 14093 16059 14151 16065
rect 14274 16056 14280 16068
rect 14332 16056 14338 16108
rect 15194 16056 15200 16108
rect 15252 16056 15258 16108
rect 13228 16000 13860 16028
rect 13228 15988 13234 16000
rect 12437 15963 12495 15969
rect 12437 15929 12449 15963
rect 12483 15960 12495 15963
rect 15304 15960 15332 16136
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16096 15439 16099
rect 17770 16096 17776 16108
rect 15427 16068 17776 16096
rect 15427 16065 15439 16068
rect 15381 16059 15439 16065
rect 17770 16056 17776 16068
rect 17828 16056 17834 16108
rect 17954 16056 17960 16108
rect 18012 16056 18018 16108
rect 18049 16099 18107 16105
rect 18049 16065 18061 16099
rect 18095 16065 18107 16099
rect 18049 16059 18107 16065
rect 18141 16099 18199 16105
rect 18141 16065 18153 16099
rect 18187 16065 18199 16099
rect 18141 16059 18199 16065
rect 16390 15988 16396 16040
rect 16448 16028 16454 16040
rect 18064 16028 18092 16059
rect 16448 16000 18092 16028
rect 18156 16028 18184 16059
rect 18322 16056 18328 16108
rect 18380 16056 18386 16108
rect 18414 16056 18420 16108
rect 18472 16056 18478 16108
rect 18690 16056 18696 16108
rect 18748 16056 18754 16108
rect 18892 16105 18920 16136
rect 19521 16133 19533 16136
rect 19567 16133 19579 16167
rect 19521 16127 19579 16133
rect 19610 16124 19616 16176
rect 19668 16124 19674 16176
rect 21008 16173 21036 16204
rect 23382 16192 23388 16204
rect 23440 16192 23446 16244
rect 23658 16192 23664 16244
rect 23716 16232 23722 16244
rect 23716 16204 23980 16232
rect 23716 16192 23722 16204
rect 20073 16167 20131 16173
rect 20073 16164 20085 16167
rect 19904 16136 20085 16164
rect 19904 16108 19932 16136
rect 20073 16133 20085 16136
rect 20119 16133 20131 16167
rect 20993 16167 21051 16173
rect 20993 16164 21005 16167
rect 20073 16127 20131 16133
rect 20548 16136 21005 16164
rect 18785 16099 18843 16105
rect 18785 16065 18797 16099
rect 18831 16065 18843 16099
rect 18785 16059 18843 16065
rect 18877 16099 18935 16105
rect 18877 16065 18889 16099
rect 18923 16065 18935 16099
rect 18877 16059 18935 16065
rect 18708 16028 18736 16056
rect 18156 16000 18736 16028
rect 18800 16028 18828 16059
rect 18966 16056 18972 16108
rect 19024 16094 19030 16108
rect 19245 16099 19303 16105
rect 19245 16096 19257 16099
rect 19076 16094 19257 16096
rect 19024 16068 19257 16094
rect 19024 16066 19104 16068
rect 19024 16056 19030 16066
rect 19245 16065 19257 16068
rect 19291 16065 19303 16099
rect 19245 16059 19303 16065
rect 19393 16099 19451 16105
rect 19393 16065 19405 16099
rect 19439 16086 19451 16099
rect 19751 16099 19809 16105
rect 19439 16065 19564 16086
rect 19393 16059 19564 16065
rect 19751 16065 19763 16099
rect 19797 16065 19809 16099
rect 19751 16059 19809 16065
rect 19408 16058 19564 16059
rect 19536 16028 19564 16058
rect 19766 16028 19794 16059
rect 19886 16056 19892 16108
rect 19944 16056 19950 16108
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20548 16105 20576 16136
rect 20993 16133 21005 16136
rect 21039 16133 21051 16167
rect 23842 16164 23848 16176
rect 20993 16127 21051 16133
rect 21376 16136 23848 16164
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 20036 16068 20269 16096
rect 20036 16056 20042 16068
rect 20257 16065 20269 16068
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 20533 16099 20591 16105
rect 20533 16065 20545 16099
rect 20579 16065 20591 16099
rect 21174 16096 21180 16108
rect 20533 16059 20591 16065
rect 20640 16068 21180 16096
rect 20441 16031 20499 16037
rect 20441 16028 20453 16031
rect 18800 16000 19334 16028
rect 19536 16000 19656 16028
rect 19766 16000 20453 16028
rect 16448 15988 16454 16000
rect 12483 15932 15332 15960
rect 12483 15929 12495 15932
rect 12437 15923 12495 15929
rect 12032 15864 12388 15892
rect 12032 15852 12038 15864
rect 16758 15852 16764 15904
rect 16816 15892 16822 15904
rect 16868 15901 16896 16000
rect 17681 15963 17739 15969
rect 17681 15929 17693 15963
rect 17727 15960 17739 15963
rect 17862 15960 17868 15972
rect 17727 15932 17868 15960
rect 17727 15929 17739 15932
rect 17681 15923 17739 15929
rect 17862 15920 17868 15932
rect 17920 15960 17926 15972
rect 18156 15960 18184 16000
rect 17920 15932 18184 15960
rect 18693 15963 18751 15969
rect 17920 15920 17926 15932
rect 18693 15929 18705 15963
rect 18739 15960 18751 15963
rect 18800 15960 18828 16000
rect 18739 15932 18828 15960
rect 19306 15960 19334 16000
rect 19628 15960 19656 16000
rect 20441 15997 20453 16000
rect 20487 15997 20499 16031
rect 20441 15991 20499 15997
rect 19306 15932 19564 15960
rect 19628 15932 20024 15960
rect 18739 15929 18751 15932
rect 18693 15923 18751 15929
rect 16853 15895 16911 15901
rect 16853 15892 16865 15895
rect 16816 15864 16865 15892
rect 16816 15852 16822 15864
rect 16853 15861 16865 15864
rect 16899 15861 16911 15895
rect 16853 15855 16911 15861
rect 17034 15852 17040 15904
rect 17092 15892 17098 15904
rect 17954 15892 17960 15904
rect 17092 15864 17960 15892
rect 17092 15852 17098 15864
rect 17954 15852 17960 15864
rect 18012 15852 18018 15904
rect 18969 15895 19027 15901
rect 18969 15861 18981 15895
rect 19015 15892 19027 15895
rect 19334 15892 19340 15904
rect 19015 15864 19340 15892
rect 19015 15861 19027 15864
rect 18969 15855 19027 15861
rect 19334 15852 19340 15864
rect 19392 15852 19398 15904
rect 19536 15892 19564 15932
rect 19886 15892 19892 15904
rect 19536 15864 19892 15892
rect 19886 15852 19892 15864
rect 19944 15852 19950 15904
rect 19996 15892 20024 15932
rect 20070 15920 20076 15972
rect 20128 15960 20134 15972
rect 20548 15960 20576 16059
rect 20128 15932 20576 15960
rect 20128 15920 20134 15932
rect 20640 15901 20668 16068
rect 21174 16056 21180 16068
rect 21232 16056 21238 16108
rect 21376 16105 21404 16136
rect 23842 16124 23848 16136
rect 23900 16124 23906 16176
rect 23952 16164 23980 16204
rect 25222 16192 25228 16244
rect 25280 16232 25286 16244
rect 26142 16232 26148 16244
rect 25280 16204 26148 16232
rect 25280 16192 25286 16204
rect 26142 16192 26148 16204
rect 26200 16192 26206 16244
rect 32398 16192 32404 16244
rect 32456 16232 32462 16244
rect 32493 16235 32551 16241
rect 32493 16232 32505 16235
rect 32456 16204 32505 16232
rect 32456 16192 32462 16204
rect 32493 16201 32505 16204
rect 32539 16201 32551 16235
rect 32493 16195 32551 16201
rect 33042 16192 33048 16244
rect 33100 16192 33106 16244
rect 34885 16235 34943 16241
rect 34885 16201 34897 16235
rect 34931 16232 34943 16235
rect 35268 16232 35296 16544
rect 34931 16204 35296 16232
rect 34931 16201 34943 16204
rect 34885 16195 34943 16201
rect 28629 16167 28687 16173
rect 28629 16164 28641 16167
rect 23952 16136 28641 16164
rect 21361 16099 21419 16105
rect 21361 16065 21373 16099
rect 21407 16065 21419 16099
rect 21361 16059 21419 16065
rect 22005 16099 22063 16105
rect 22005 16065 22017 16099
rect 22051 16096 22063 16099
rect 22554 16096 22560 16108
rect 22051 16068 22560 16096
rect 22051 16065 22063 16068
rect 22005 16059 22063 16065
rect 21376 16028 21404 16059
rect 22554 16056 22560 16068
rect 22612 16056 22618 16108
rect 23290 16056 23296 16108
rect 23348 16056 23354 16108
rect 21008 16000 21404 16028
rect 21008 15904 21036 16000
rect 21634 15988 21640 16040
rect 21692 16028 21698 16040
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21692 16000 21925 16028
rect 21692 15988 21698 16000
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15960 21419 15963
rect 23952 15960 23980 16136
rect 28629 16133 28641 16136
rect 28675 16133 28687 16167
rect 28629 16127 28687 16133
rect 29638 16124 29644 16176
rect 29696 16124 29702 16176
rect 25406 16096 25412 16108
rect 21407 15932 23980 15960
rect 25240 16068 25412 16096
rect 21407 15929 21419 15932
rect 21361 15923 21419 15929
rect 25240 15904 25268 16068
rect 25406 16056 25412 16068
rect 25464 16056 25470 16108
rect 25593 16099 25651 16105
rect 25593 16065 25605 16099
rect 25639 16096 25651 16099
rect 25866 16096 25872 16108
rect 25639 16068 25872 16096
rect 25639 16065 25651 16068
rect 25593 16059 25651 16065
rect 25866 16056 25872 16068
rect 25924 16056 25930 16108
rect 25961 16099 26019 16105
rect 25961 16065 25973 16099
rect 26007 16065 26019 16099
rect 25961 16059 26019 16065
rect 25501 16031 25559 16037
rect 25501 15997 25513 16031
rect 25547 16028 25559 16031
rect 25976 16028 26004 16059
rect 26234 16056 26240 16108
rect 26292 16056 26298 16108
rect 31938 16056 31944 16108
rect 31996 16096 32002 16108
rect 32125 16099 32183 16105
rect 32125 16096 32137 16099
rect 31996 16068 32137 16096
rect 31996 16056 32002 16068
rect 32125 16065 32137 16068
rect 32171 16065 32183 16099
rect 32125 16059 32183 16065
rect 32306 16056 32312 16108
rect 32364 16056 32370 16108
rect 33060 16096 33088 16192
rect 34146 16124 34152 16176
rect 34204 16124 34210 16176
rect 33137 16099 33195 16105
rect 33137 16096 33149 16099
rect 33060 16068 33149 16096
rect 33137 16065 33149 16068
rect 33183 16065 33195 16099
rect 33137 16059 33195 16065
rect 25547 16000 26004 16028
rect 26789 16031 26847 16037
rect 25547 15997 25559 16000
rect 25501 15991 25559 15997
rect 26789 15997 26801 16031
rect 26835 16028 26847 16031
rect 26970 16028 26976 16040
rect 26835 16000 26976 16028
rect 26835 15997 26847 16000
rect 26789 15991 26847 15997
rect 26970 15988 26976 16000
rect 27028 15988 27034 16040
rect 28261 16031 28319 16037
rect 28261 15997 28273 16031
rect 28307 16028 28319 16031
rect 28353 16031 28411 16037
rect 28353 16028 28365 16031
rect 28307 16000 28365 16028
rect 28307 15997 28319 16000
rect 28261 15991 28319 15997
rect 28353 15997 28365 16000
rect 28399 15997 28411 16031
rect 28353 15991 28411 15997
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 19996 15864 20637 15892
rect 20625 15861 20637 15864
rect 20671 15861 20683 15895
rect 20625 15855 20683 15861
rect 20990 15852 20996 15904
rect 21048 15852 21054 15904
rect 22094 15852 22100 15904
rect 22152 15892 22158 15904
rect 22373 15895 22431 15901
rect 22373 15892 22385 15895
rect 22152 15864 22385 15892
rect 22152 15852 22158 15864
rect 22373 15861 22385 15864
rect 22419 15861 22431 15895
rect 22373 15855 22431 15861
rect 24949 15895 25007 15901
rect 24949 15861 24961 15895
rect 24995 15892 25007 15895
rect 25130 15892 25136 15904
rect 24995 15864 25136 15892
rect 24995 15861 25007 15864
rect 24949 15855 25007 15861
rect 25130 15852 25136 15864
rect 25188 15852 25194 15904
rect 25222 15852 25228 15904
rect 25280 15852 25286 15904
rect 28368 15892 28396 15991
rect 33410 15988 33416 16040
rect 33468 15988 33474 16040
rect 29270 15892 29276 15904
rect 28368 15864 29276 15892
rect 29270 15852 29276 15864
rect 29328 15852 29334 15904
rect 30101 15895 30159 15901
rect 30101 15861 30113 15895
rect 30147 15892 30159 15895
rect 31110 15892 31116 15904
rect 30147 15864 31116 15892
rect 30147 15861 30159 15864
rect 30101 15855 30159 15861
rect 31110 15852 31116 15864
rect 31168 15852 31174 15904
rect 1104 15802 35248 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 35248 15802
rect 1104 15728 35248 15750
rect 3326 15648 3332 15700
rect 3384 15648 3390 15700
rect 4798 15648 4804 15700
rect 4856 15648 4862 15700
rect 5074 15648 5080 15700
rect 5132 15688 5138 15700
rect 5261 15691 5319 15697
rect 5261 15688 5273 15691
rect 5132 15660 5273 15688
rect 5132 15648 5138 15660
rect 5261 15657 5273 15660
rect 5307 15657 5319 15691
rect 5261 15651 5319 15657
rect 12066 15648 12072 15700
rect 12124 15688 12130 15700
rect 12253 15691 12311 15697
rect 12253 15688 12265 15691
rect 12124 15660 12265 15688
rect 12124 15648 12130 15660
rect 12253 15657 12265 15660
rect 12299 15657 12311 15691
rect 12253 15651 12311 15657
rect 12621 15691 12679 15697
rect 12621 15657 12633 15691
rect 12667 15688 12679 15691
rect 12986 15688 12992 15700
rect 12667 15660 12992 15688
rect 12667 15657 12679 15660
rect 12621 15651 12679 15657
rect 12986 15648 12992 15660
rect 13044 15648 13050 15700
rect 13173 15691 13231 15697
rect 13173 15657 13185 15691
rect 13219 15688 13231 15691
rect 13354 15688 13360 15700
rect 13219 15660 13360 15688
rect 13219 15657 13231 15660
rect 13173 15651 13231 15657
rect 13354 15648 13360 15660
rect 13412 15648 13418 15700
rect 13538 15648 13544 15700
rect 13596 15648 13602 15700
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15657 14795 15691
rect 14737 15651 14795 15657
rect 4816 15552 4844 15648
rect 13081 15623 13139 15629
rect 13081 15589 13093 15623
rect 13127 15620 13139 15623
rect 14752 15620 14780 15651
rect 15194 15648 15200 15700
rect 15252 15648 15258 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 17862 15688 17868 15700
rect 17552 15660 17868 15688
rect 17552 15648 17558 15660
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18601 15691 18659 15697
rect 18601 15688 18613 15691
rect 18012 15660 18613 15688
rect 18012 15648 18018 15660
rect 18601 15657 18613 15660
rect 18647 15657 18659 15691
rect 18601 15651 18659 15657
rect 19429 15691 19487 15697
rect 19429 15657 19441 15691
rect 19475 15688 19487 15691
rect 19518 15688 19524 15700
rect 19475 15660 19524 15688
rect 19475 15657 19487 15660
rect 19429 15651 19487 15657
rect 13127 15592 14780 15620
rect 13127 15589 13139 15592
rect 13081 15583 13139 15589
rect 15102 15580 15108 15632
rect 15160 15620 15166 15632
rect 18322 15620 18328 15632
rect 15160 15592 18328 15620
rect 15160 15580 15166 15592
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 6273 15555 6331 15561
rect 6273 15552 6285 15555
rect 4816 15524 6285 15552
rect 6273 15521 6285 15524
rect 6319 15521 6331 15555
rect 6273 15515 6331 15521
rect 8478 15512 8484 15564
rect 8536 15552 8542 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 8536 15524 9597 15552
rect 8536 15512 8542 15524
rect 1581 15487 1639 15493
rect 1581 15453 1593 15487
rect 1627 15453 1639 15487
rect 1581 15447 1639 15453
rect 1596 15416 1624 15447
rect 3602 15444 3608 15496
rect 3660 15484 3666 15496
rect 4617 15487 4675 15493
rect 3660 15456 3832 15484
rect 3660 15444 3666 15456
rect 1596 15388 1716 15416
rect 1688 15360 1716 15388
rect 1854 15376 1860 15428
rect 1912 15376 1918 15428
rect 3513 15419 3571 15425
rect 3513 15416 3525 15419
rect 3082 15388 3525 15416
rect 3513 15385 3525 15388
rect 3559 15385 3571 15419
rect 3513 15379 3571 15385
rect 3804 15360 3832 15456
rect 4617 15453 4629 15487
rect 4663 15453 4675 15487
rect 4617 15447 4675 15453
rect 1670 15308 1676 15360
rect 1728 15308 1734 15360
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 3973 15351 4031 15357
rect 3973 15348 3985 15351
rect 3844 15320 3985 15348
rect 3844 15308 3850 15320
rect 3973 15317 3985 15320
rect 4019 15317 4031 15351
rect 4632 15348 4660 15447
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4764 15456 4813 15484
rect 4764 15444 4770 15456
rect 4801 15453 4813 15456
rect 4847 15484 4859 15487
rect 4847 15456 5672 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 5644 15428 5672 15456
rect 5902 15444 5908 15496
rect 5960 15484 5966 15496
rect 5997 15487 6055 15493
rect 5997 15484 6009 15487
rect 5960 15456 6009 15484
rect 5960 15444 5966 15456
rect 5997 15453 6009 15456
rect 6043 15453 6055 15487
rect 5997 15447 6055 15453
rect 8018 15444 8024 15496
rect 8076 15484 8082 15496
rect 8076 15456 8432 15484
rect 8076 15444 8082 15456
rect 4985 15419 5043 15425
rect 4985 15385 4997 15419
rect 5031 15416 5043 15419
rect 5169 15419 5227 15425
rect 5169 15416 5181 15419
rect 5031 15388 5181 15416
rect 5031 15385 5043 15388
rect 4985 15379 5043 15385
rect 5169 15385 5181 15388
rect 5215 15385 5227 15419
rect 5169 15379 5227 15385
rect 5442 15376 5448 15428
rect 5500 15376 5506 15428
rect 5626 15376 5632 15428
rect 5684 15376 5690 15428
rect 7929 15419 7987 15425
rect 7929 15416 7941 15419
rect 7498 15388 7941 15416
rect 7929 15385 7941 15388
rect 7975 15385 7987 15419
rect 7929 15379 7987 15385
rect 4890 15348 4896 15360
rect 4632 15320 4896 15348
rect 3973 15311 4031 15317
rect 4890 15308 4896 15320
rect 4948 15348 4954 15360
rect 5460 15348 5488 15376
rect 4948 15320 5488 15348
rect 4948 15308 4954 15320
rect 7742 15308 7748 15360
rect 7800 15308 7806 15360
rect 8404 15357 8432 15456
rect 8772 15360 8800 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15552 9919 15555
rect 9950 15552 9956 15564
rect 9907 15524 9956 15552
rect 9907 15521 9919 15524
rect 9861 15515 9919 15521
rect 9950 15512 9956 15524
rect 10008 15512 10014 15564
rect 12802 15512 12808 15564
rect 12860 15552 12866 15564
rect 13265 15555 13323 15561
rect 12860 15524 13216 15552
rect 12860 15512 12866 15524
rect 11974 15444 11980 15496
rect 12032 15484 12038 15496
rect 12069 15487 12127 15493
rect 12069 15484 12081 15487
rect 12032 15456 12081 15484
rect 12032 15444 12038 15456
rect 12069 15453 12081 15456
rect 12115 15453 12127 15487
rect 12069 15447 12127 15453
rect 12618 15444 12624 15496
rect 12676 15444 12682 15496
rect 12912 15493 12940 15524
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15453 12955 15487
rect 12897 15447 12955 15453
rect 12989 15487 13047 15493
rect 12989 15453 13001 15487
rect 13035 15453 13047 15487
rect 12989 15447 13047 15453
rect 10594 15376 10600 15428
rect 10652 15376 10658 15428
rect 11793 15419 11851 15425
rect 11793 15385 11805 15419
rect 11839 15416 11851 15419
rect 11885 15419 11943 15425
rect 11885 15416 11897 15419
rect 11839 15388 11897 15416
rect 11839 15385 11851 15388
rect 11793 15379 11851 15385
rect 11885 15385 11897 15388
rect 11931 15416 11943 15419
rect 12636 15416 12664 15444
rect 11931 15388 12664 15416
rect 12805 15419 12863 15425
rect 11931 15385 11943 15388
rect 11885 15379 11943 15385
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 13004 15416 13032 15447
rect 12851 15388 13032 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 8389 15351 8447 15357
rect 8389 15317 8401 15351
rect 8435 15348 8447 15351
rect 8570 15348 8576 15360
rect 8435 15320 8576 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 8754 15308 8760 15360
rect 8812 15308 8818 15360
rect 11330 15308 11336 15360
rect 11388 15308 11394 15360
rect 13188 15348 13216 15524
rect 13265 15521 13277 15555
rect 13311 15521 13323 15555
rect 13265 15515 13323 15521
rect 13817 15555 13875 15561
rect 13817 15521 13829 15555
rect 13863 15552 13875 15555
rect 14369 15555 14427 15561
rect 14369 15552 14381 15555
rect 13863 15524 14381 15552
rect 13863 15521 13875 15524
rect 13817 15515 13875 15521
rect 14369 15521 14381 15524
rect 14415 15521 14427 15555
rect 14369 15515 14427 15521
rect 13280 15416 13308 15515
rect 14458 15512 14464 15564
rect 14516 15552 14522 15564
rect 15197 15555 15255 15561
rect 14516 15524 14964 15552
rect 14516 15512 14522 15524
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15484 13415 15487
rect 13446 15484 13452 15496
rect 13403 15456 13452 15484
rect 13403 15453 13415 15456
rect 13357 15447 13415 15453
rect 13446 15444 13452 15456
rect 13504 15444 13510 15496
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 14274 15444 14280 15496
rect 14332 15444 14338 15496
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 14642 15484 14648 15496
rect 14599 15456 14648 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 14936 15416 14964 15524
rect 15197 15521 15209 15555
rect 15243 15552 15255 15555
rect 15286 15552 15292 15564
rect 15243 15524 15292 15552
rect 15243 15521 15255 15524
rect 15197 15515 15255 15521
rect 15286 15512 15292 15524
rect 15344 15552 15350 15564
rect 16485 15555 16543 15561
rect 15344 15524 15700 15552
rect 15344 15512 15350 15524
rect 15010 15444 15016 15496
rect 15068 15484 15074 15496
rect 15672 15493 15700 15524
rect 16485 15521 16497 15555
rect 16531 15552 16543 15555
rect 16666 15552 16672 15564
rect 16531 15524 16672 15552
rect 16531 15521 16543 15524
rect 16485 15515 16543 15521
rect 16666 15512 16672 15524
rect 16724 15512 16730 15564
rect 16868 15524 17908 15552
rect 15657 15487 15715 15493
rect 15068 15456 15608 15484
rect 15068 15444 15074 15456
rect 15289 15419 15347 15425
rect 15289 15416 15301 15419
rect 13280 15388 14872 15416
rect 14936 15388 15301 15416
rect 14734 15348 14740 15360
rect 13188 15320 14740 15348
rect 14734 15308 14740 15320
rect 14792 15308 14798 15360
rect 14844 15357 14872 15388
rect 15289 15385 15301 15388
rect 15335 15385 15347 15419
rect 15580 15416 15608 15456
rect 15657 15453 15669 15487
rect 15703 15453 15715 15487
rect 15657 15447 15715 15453
rect 16114 15444 16120 15496
rect 16172 15444 16178 15496
rect 16868 15428 16896 15524
rect 17880 15493 17908 15524
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 17236 15456 17693 15484
rect 16850 15416 16856 15428
rect 15580 15388 16856 15416
rect 15289 15379 15347 15385
rect 16850 15376 16856 15388
rect 16908 15376 16914 15428
rect 17236 15360 17264 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 17865 15487 17923 15493
rect 17865 15453 17877 15487
rect 17911 15453 17923 15487
rect 18340 15484 18368 15580
rect 18616 15552 18644 15651
rect 19518 15648 19524 15660
rect 19576 15648 19582 15700
rect 25501 15691 25559 15697
rect 25501 15657 25513 15691
rect 25547 15688 25559 15691
rect 25866 15688 25872 15700
rect 25547 15660 25872 15688
rect 25547 15657 25559 15660
rect 25501 15651 25559 15657
rect 25866 15648 25872 15660
rect 25924 15648 25930 15700
rect 29270 15648 29276 15700
rect 29328 15648 29334 15700
rect 32217 15691 32275 15697
rect 32217 15657 32229 15691
rect 32263 15688 32275 15691
rect 33410 15688 33416 15700
rect 32263 15660 33416 15688
rect 32263 15657 32275 15660
rect 32217 15651 32275 15657
rect 33410 15648 33416 15660
rect 33468 15648 33474 15700
rect 34146 15648 34152 15700
rect 34204 15648 34210 15700
rect 18966 15580 18972 15632
rect 19024 15620 19030 15632
rect 19024 15592 19840 15620
rect 19024 15580 19030 15592
rect 18616 15524 19564 15552
rect 19150 15484 19156 15496
rect 18340 15456 19156 15484
rect 17865 15447 17923 15453
rect 19150 15444 19156 15456
rect 19208 15484 19214 15496
rect 19536 15493 19564 15524
rect 19812 15493 19840 15592
rect 26970 15512 26976 15564
rect 27028 15552 27034 15564
rect 29288 15552 29316 15648
rect 31297 15623 31355 15629
rect 31297 15589 31309 15623
rect 31343 15620 31355 15623
rect 32306 15620 32312 15632
rect 31343 15592 32312 15620
rect 31343 15589 31355 15592
rect 31297 15583 31355 15589
rect 29549 15555 29607 15561
rect 29549 15552 29561 15555
rect 27028 15524 27108 15552
rect 29288 15524 29561 15552
rect 27028 15512 27034 15524
rect 19337 15487 19395 15493
rect 19337 15484 19349 15487
rect 19208 15456 19349 15484
rect 19208 15444 19214 15456
rect 19337 15453 19349 15456
rect 19383 15453 19395 15487
rect 19337 15447 19395 15453
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19613 15487 19671 15493
rect 19613 15453 19625 15487
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15453 19855 15487
rect 19797 15447 19855 15453
rect 23293 15487 23351 15493
rect 23293 15453 23305 15487
rect 23339 15484 23351 15487
rect 23382 15484 23388 15496
rect 23339 15456 23388 15484
rect 23339 15453 23351 15456
rect 23293 15447 23351 15453
rect 18325 15419 18383 15425
rect 18325 15385 18337 15419
rect 18371 15416 18383 15419
rect 18598 15416 18604 15428
rect 18371 15388 18604 15416
rect 18371 15385 18383 15388
rect 18325 15379 18383 15385
rect 18598 15376 18604 15388
rect 18656 15376 18662 15428
rect 18966 15376 18972 15428
rect 19024 15376 19030 15428
rect 19628 15416 19656 15447
rect 23382 15444 23388 15456
rect 23440 15444 23446 15496
rect 27080 15493 27108 15524
rect 29549 15521 29561 15524
rect 29595 15521 29607 15555
rect 29549 15515 29607 15521
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15453 23627 15487
rect 23569 15447 23627 15453
rect 26887 15487 26945 15493
rect 26887 15453 26899 15487
rect 26933 15484 26945 15487
rect 27065 15487 27123 15493
rect 26933 15456 27016 15484
rect 26933 15453 26945 15456
rect 26887 15447 26945 15453
rect 20070 15416 20076 15428
rect 19076 15388 20076 15416
rect 14829 15351 14887 15357
rect 14829 15317 14841 15351
rect 14875 15317 14887 15351
rect 14829 15311 14887 15317
rect 16666 15308 16672 15360
rect 16724 15348 16730 15360
rect 17034 15348 17040 15360
rect 16724 15320 17040 15348
rect 16724 15308 16730 15320
rect 17034 15308 17040 15320
rect 17092 15308 17098 15360
rect 17218 15308 17224 15360
rect 17276 15308 17282 15360
rect 17862 15308 17868 15360
rect 17920 15308 17926 15360
rect 18414 15308 18420 15360
rect 18472 15348 18478 15360
rect 18874 15348 18880 15360
rect 18472 15320 18880 15348
rect 18472 15308 18478 15320
rect 18874 15308 18880 15320
rect 18932 15348 18938 15360
rect 19076 15348 19104 15388
rect 20070 15376 20076 15388
rect 20128 15376 20134 15428
rect 22738 15376 22744 15428
rect 22796 15416 22802 15428
rect 23474 15416 23480 15428
rect 22796 15388 23480 15416
rect 22796 15376 22802 15388
rect 23474 15376 23480 15388
rect 23532 15416 23538 15428
rect 23584 15416 23612 15447
rect 23532 15388 23612 15416
rect 26988 15416 27016 15456
rect 27065 15453 27077 15487
rect 27111 15484 27123 15487
rect 27522 15484 27528 15496
rect 27111 15456 27528 15484
rect 27111 15453 27123 15456
rect 27065 15447 27123 15453
rect 27522 15444 27528 15456
rect 27580 15444 27586 15496
rect 31202 15444 31208 15496
rect 31260 15484 31266 15496
rect 31956 15493 31984 15592
rect 32306 15580 32312 15592
rect 32364 15580 32370 15632
rect 32582 15580 32588 15632
rect 32640 15580 32646 15632
rect 32033 15555 32091 15561
rect 32033 15521 32045 15555
rect 32079 15552 32091 15555
rect 32493 15555 32551 15561
rect 32493 15552 32505 15555
rect 32079 15524 32505 15552
rect 32079 15521 32091 15524
rect 32033 15515 32091 15521
rect 32493 15521 32505 15524
rect 32539 15521 32551 15555
rect 32493 15515 32551 15521
rect 32600 15493 32628 15580
rect 31389 15487 31447 15493
rect 31389 15484 31401 15487
rect 31260 15456 31401 15484
rect 31260 15444 31266 15456
rect 31389 15453 31401 15456
rect 31435 15453 31447 15487
rect 31389 15447 31447 15453
rect 31941 15487 31999 15493
rect 31941 15453 31953 15487
rect 31987 15453 31999 15487
rect 31941 15447 31999 15453
rect 32401 15487 32459 15493
rect 32401 15453 32413 15487
rect 32447 15453 32459 15487
rect 32401 15447 32459 15453
rect 32585 15487 32643 15493
rect 32585 15453 32597 15487
rect 32631 15453 32643 15487
rect 34057 15487 34115 15493
rect 34057 15484 34069 15487
rect 32585 15447 32643 15453
rect 33888 15456 34069 15484
rect 27154 15416 27160 15428
rect 26988 15388 27160 15416
rect 23532 15376 23538 15388
rect 27154 15376 27160 15388
rect 27212 15376 27218 15428
rect 28994 15376 29000 15428
rect 29052 15416 29058 15428
rect 29825 15419 29883 15425
rect 29825 15416 29837 15419
rect 29052 15388 29837 15416
rect 29052 15376 29058 15388
rect 29825 15385 29837 15388
rect 29871 15385 29883 15419
rect 31481 15419 31539 15425
rect 31481 15416 31493 15419
rect 31050 15388 31493 15416
rect 29825 15379 29883 15385
rect 31481 15385 31493 15388
rect 31527 15385 31539 15419
rect 32416 15416 32444 15447
rect 31481 15379 31539 15385
rect 31956 15388 32444 15416
rect 31956 15360 31984 15388
rect 33888 15360 33916 15456
rect 34057 15453 34069 15456
rect 34103 15484 34115 15487
rect 34330 15484 34336 15496
rect 34103 15456 34336 15484
rect 34103 15453 34115 15456
rect 34057 15447 34115 15453
rect 34330 15444 34336 15456
rect 34388 15444 34394 15496
rect 18932 15320 19104 15348
rect 18932 15308 18938 15320
rect 19334 15308 19340 15360
rect 19392 15348 19398 15360
rect 19705 15351 19763 15357
rect 19705 15348 19717 15351
rect 19392 15320 19717 15348
rect 19392 15308 19398 15320
rect 19705 15317 19717 15320
rect 19751 15348 19763 15351
rect 19978 15348 19984 15360
rect 19751 15320 19984 15348
rect 19751 15317 19763 15320
rect 19705 15311 19763 15317
rect 19978 15308 19984 15320
rect 20036 15308 20042 15360
rect 20990 15308 20996 15360
rect 21048 15308 21054 15360
rect 21082 15308 21088 15360
rect 21140 15348 21146 15360
rect 21361 15351 21419 15357
rect 21361 15348 21373 15351
rect 21140 15320 21373 15348
rect 21140 15308 21146 15320
rect 21361 15317 21373 15320
rect 21407 15317 21419 15351
rect 21361 15311 21419 15317
rect 21910 15308 21916 15360
rect 21968 15348 21974 15360
rect 23198 15348 23204 15360
rect 21968 15320 23204 15348
rect 21968 15308 21974 15320
rect 23198 15308 23204 15320
rect 23256 15308 23262 15360
rect 23385 15351 23443 15357
rect 23385 15317 23397 15351
rect 23431 15348 23443 15351
rect 23658 15348 23664 15360
rect 23431 15320 23664 15348
rect 23431 15317 23443 15320
rect 23385 15311 23443 15317
rect 23658 15308 23664 15320
rect 23716 15308 23722 15360
rect 23750 15308 23756 15360
rect 23808 15308 23814 15360
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 25222 15348 25228 15360
rect 25087 15320 25228 15348
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 25222 15308 25228 15320
rect 25280 15348 25286 15360
rect 25682 15348 25688 15360
rect 25280 15320 25688 15348
rect 25280 15308 25286 15320
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 25961 15351 26019 15357
rect 25961 15317 25973 15351
rect 26007 15348 26019 15351
rect 26510 15348 26516 15360
rect 26007 15320 26516 15348
rect 26007 15317 26019 15320
rect 25961 15311 26019 15317
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 27065 15351 27123 15357
rect 27065 15317 27077 15351
rect 27111 15348 27123 15351
rect 27614 15348 27620 15360
rect 27111 15320 27620 15348
rect 27111 15317 27123 15320
rect 27065 15311 27123 15317
rect 27614 15308 27620 15320
rect 27672 15308 27678 15360
rect 31938 15308 31944 15360
rect 31996 15308 32002 15360
rect 33870 15308 33876 15360
rect 33928 15308 33934 15360
rect 1104 15258 35236 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 35236 15258
rect 1104 15184 35236 15206
rect 1581 15147 1639 15153
rect 1581 15113 1593 15147
rect 1627 15144 1639 15147
rect 1854 15144 1860 15156
rect 1627 15116 1860 15144
rect 1627 15113 1639 15116
rect 1581 15107 1639 15113
rect 1854 15104 1860 15116
rect 1912 15104 1918 15156
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 10689 15147 10747 15153
rect 10689 15144 10701 15147
rect 10652 15116 10701 15144
rect 10652 15104 10658 15116
rect 10689 15113 10701 15116
rect 10735 15113 10747 15147
rect 10689 15107 10747 15113
rect 11330 15104 11336 15156
rect 11388 15144 11394 15156
rect 11388 15116 12296 15144
rect 11388 15104 11394 15116
rect 11241 15079 11299 15085
rect 11241 15045 11253 15079
rect 11287 15076 11299 15079
rect 11974 15076 11980 15088
rect 11287 15048 11980 15076
rect 11287 15045 11299 15048
rect 11241 15039 11299 15045
rect 11974 15036 11980 15048
rect 12032 15036 12038 15088
rect 934 14968 940 15020
rect 992 15008 998 15020
rect 1397 15011 1455 15017
rect 1397 15008 1409 15011
rect 992 14980 1409 15008
rect 992 14968 998 14980
rect 1397 14977 1409 14980
rect 1443 14977 1455 15011
rect 1397 14971 1455 14977
rect 7742 14968 7748 15020
rect 7800 15008 7806 15020
rect 8113 15011 8171 15017
rect 8113 15008 8125 15011
rect 7800 14980 8125 15008
rect 7800 14968 7806 14980
rect 8113 14977 8125 14980
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 14977 10655 15011
rect 10597 14971 10655 14977
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 10410 14940 10416 14952
rect 8987 14912 10416 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 3510 14764 3516 14816
rect 3568 14804 3574 14816
rect 5902 14804 5908 14816
rect 3568 14776 5908 14804
rect 3568 14764 3574 14776
rect 5902 14764 5908 14776
rect 5960 14764 5966 14816
rect 10428 14804 10456 14900
rect 10502 14832 10508 14884
rect 10560 14872 10566 14884
rect 10612 14872 10640 14971
rect 11606 14968 11612 15020
rect 11664 14968 11670 15020
rect 12268 15017 12296 15116
rect 14090 15104 14096 15156
rect 14148 15104 14154 15156
rect 14274 15104 14280 15156
rect 14332 15104 14338 15156
rect 22123 15147 22181 15153
rect 15212 15116 22094 15144
rect 15212 15076 15240 15116
rect 13110 15048 15240 15076
rect 15286 15036 15292 15088
rect 15344 15036 15350 15088
rect 16485 15079 16543 15085
rect 16485 15045 16497 15079
rect 16531 15076 16543 15079
rect 17310 15076 17316 15088
rect 16531 15048 17316 15076
rect 16531 15045 16543 15048
rect 16485 15039 16543 15045
rect 17310 15036 17316 15048
rect 17368 15036 17374 15088
rect 19150 15036 19156 15088
rect 19208 15036 19214 15088
rect 21453 15079 21511 15085
rect 20732 15048 21312 15076
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13725 15014 13783 15017
rect 13725 15011 13860 15014
rect 13725 15008 13737 15011
rect 13504 14980 13737 15008
rect 13504 14968 13510 14980
rect 13725 14977 13737 14980
rect 13771 15008 13860 15011
rect 13771 14986 14320 15008
rect 13771 14977 13783 14986
rect 13832 14980 14320 14986
rect 13725 14971 13783 14977
rect 13630 14900 13636 14952
rect 13688 14900 13694 14952
rect 14292 14940 14320 14980
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14424 14980 14872 15008
rect 14424 14968 14430 14980
rect 14734 14940 14740 14952
rect 14292 14912 14740 14940
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 14844 14949 14872 14980
rect 14918 14968 14924 15020
rect 14976 14968 14982 15020
rect 15102 14968 15108 15020
rect 15160 14968 15166 15020
rect 15304 15008 15332 15036
rect 16120 15020 16172 15026
rect 15473 15011 15531 15017
rect 15473 15008 15485 15011
rect 15304 14980 15485 15008
rect 15473 14977 15485 14980
rect 15519 14977 15531 15011
rect 15473 14971 15531 14977
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16172 14980 16681 15008
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 15120 14940 15148 14968
rect 16120 14962 16172 14968
rect 14875 14912 15148 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 16574 14900 16580 14952
rect 16632 14940 16638 14952
rect 16776 14940 16804 14971
rect 16850 14968 16856 15020
rect 16908 15008 16914 15020
rect 16945 15011 17003 15017
rect 16945 15008 16957 15011
rect 16908 14980 16957 15008
rect 16908 14968 16914 14980
rect 16945 14977 16957 14980
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 17494 14968 17500 15020
rect 17552 14968 17558 15020
rect 18966 14968 18972 15020
rect 19024 15008 19030 15020
rect 20732 15017 20760 15048
rect 21284 15020 21312 15048
rect 21453 15045 21465 15079
rect 21499 15076 21511 15079
rect 21910 15076 21916 15088
rect 21499 15048 21916 15076
rect 21499 15045 21511 15048
rect 21453 15039 21511 15045
rect 21910 15036 21916 15048
rect 21968 15036 21974 15088
rect 22066 15076 22094 15116
rect 22123 15113 22135 15147
rect 22169 15144 22181 15147
rect 22278 15144 22284 15156
rect 22169 15116 22284 15144
rect 22169 15113 22181 15116
rect 22123 15107 22181 15113
rect 22278 15104 22284 15116
rect 22336 15104 22342 15156
rect 22480 15116 26464 15144
rect 22480 15076 22508 15116
rect 22066 15048 22508 15076
rect 23198 15036 23204 15088
rect 23256 15036 23262 15088
rect 24397 15079 24455 15085
rect 24397 15045 24409 15079
rect 24443 15076 24455 15079
rect 24443 15048 25176 15076
rect 24443 15045 24455 15048
rect 24397 15039 24455 15045
rect 20717 15011 20775 15017
rect 20717 15008 20729 15011
rect 19024 14980 20729 15008
rect 19024 14968 19030 14980
rect 20717 14977 20729 14980
rect 20763 14977 20775 15011
rect 21082 15008 21088 15020
rect 20717 14971 20775 14977
rect 20824 14980 21088 15008
rect 17512 14940 17540 14968
rect 20824 14952 20852 14980
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 21266 14968 21272 15020
rect 21324 14968 21330 15020
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22373 15011 22431 15017
rect 22373 15008 22385 15011
rect 22152 14980 22385 15008
rect 22152 14968 22158 14980
rect 22373 14977 22385 14980
rect 22419 14977 22431 15011
rect 22373 14971 22431 14977
rect 22465 15011 22523 15017
rect 22465 14977 22477 15011
rect 22511 14977 22523 15011
rect 22465 14971 22523 14977
rect 16632 14912 17540 14940
rect 16632 14900 16638 14912
rect 20806 14900 20812 14952
rect 20864 14900 20870 14952
rect 22186 14940 22192 14952
rect 22066 14912 22192 14940
rect 22066 14872 22094 14912
rect 22186 14900 22192 14912
rect 22244 14900 22250 14952
rect 22480 14940 22508 14971
rect 22554 14968 22560 15020
rect 22612 15008 22618 15020
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22612 14980 22661 15008
rect 22612 14968 22618 14980
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 22741 15011 22799 15017
rect 22741 14977 22753 15011
rect 22787 15008 22799 15011
rect 22830 15008 22836 15020
rect 22787 14980 22836 15008
rect 22787 14977 22799 14980
rect 22741 14971 22799 14977
rect 22830 14968 22836 14980
rect 22888 14968 22894 15020
rect 23216 15008 23244 15036
rect 23477 15011 23535 15017
rect 23477 15008 23489 15011
rect 23216 14980 23489 15008
rect 23477 14977 23489 14980
rect 23523 14977 23535 15011
rect 23477 14971 23535 14977
rect 22480 14912 23060 14940
rect 10560 14844 22094 14872
rect 22138 14844 22508 14872
rect 10560 14832 10566 14844
rect 13814 14804 13820 14816
rect 10428 14776 13820 14804
rect 13814 14764 13820 14776
rect 13872 14764 13878 14816
rect 17218 14764 17224 14816
rect 17276 14804 17282 14816
rect 17497 14807 17555 14813
rect 17497 14804 17509 14807
rect 17276 14776 17509 14804
rect 17276 14764 17282 14776
rect 17497 14773 17509 14776
rect 17543 14773 17555 14807
rect 17497 14767 17555 14773
rect 20441 14807 20499 14813
rect 20441 14773 20453 14807
rect 20487 14804 20499 14807
rect 20806 14804 20812 14816
rect 20487 14776 20812 14804
rect 20487 14773 20499 14776
rect 20441 14767 20499 14773
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 22138 14813 22166 14844
rect 22480 14816 22508 14844
rect 23032 14816 23060 14912
rect 23492 14872 23520 14971
rect 23566 14968 23572 15020
rect 23624 15008 23630 15020
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23624 14980 23857 15008
rect 23624 14968 23630 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 24302 14968 24308 15020
rect 24360 14968 24366 15020
rect 24578 14968 24584 15020
rect 24636 14968 24642 15020
rect 24762 14968 24768 15020
rect 24820 14968 24826 15020
rect 25148 15017 25176 15048
rect 25133 15011 25191 15017
rect 25133 14977 25145 15011
rect 25179 15008 25191 15011
rect 25222 15008 25228 15020
rect 25179 14980 25228 15008
rect 25179 14977 25191 14980
rect 25133 14971 25191 14977
rect 25222 14968 25228 14980
rect 25280 14968 25286 15020
rect 23750 14900 23756 14952
rect 23808 14900 23814 14952
rect 25041 14943 25099 14949
rect 25041 14909 25053 14943
rect 25087 14909 25099 14943
rect 25041 14903 25099 14909
rect 24118 14872 24124 14884
rect 23492 14844 24124 14872
rect 24118 14832 24124 14844
rect 24176 14832 24182 14884
rect 24213 14875 24271 14881
rect 24213 14841 24225 14875
rect 24259 14872 24271 14875
rect 25056 14872 25084 14903
rect 26326 14900 26332 14952
rect 26384 14900 26390 14952
rect 26436 14940 26464 15116
rect 27154 15104 27160 15156
rect 27212 15144 27218 15156
rect 27212 15116 27568 15144
rect 27212 15104 27218 15116
rect 26528 15048 27476 15076
rect 26528 15017 26556 15048
rect 26513 15011 26571 15017
rect 26513 14977 26525 15011
rect 26559 14977 26571 15011
rect 26513 14971 26571 14977
rect 26697 15011 26755 15017
rect 26697 14977 26709 15011
rect 26743 14977 26755 15011
rect 26697 14971 26755 14977
rect 26602 14940 26608 14952
rect 26436 14912 26608 14940
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 26712 14940 26740 14971
rect 26786 14968 26792 15020
rect 26844 15008 26850 15020
rect 27157 15011 27215 15017
rect 27157 15008 27169 15011
rect 26844 14980 27169 15008
rect 26844 14968 26850 14980
rect 27157 14977 27169 14980
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27246 14968 27252 15020
rect 27304 14968 27310 15020
rect 27062 14940 27068 14952
rect 26712 14912 27068 14940
rect 27062 14900 27068 14912
rect 27120 14940 27126 14952
rect 27264 14940 27292 14968
rect 27120 14912 27292 14940
rect 27448 14940 27476 15048
rect 27540 15008 27568 15116
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 32217 15147 32275 15153
rect 27672 15116 27752 15144
rect 27672 15104 27678 15116
rect 27724 15076 27752 15116
rect 32217 15113 32229 15147
rect 32263 15144 32275 15147
rect 32582 15144 32588 15156
rect 32263 15116 32588 15144
rect 32263 15113 32275 15116
rect 32217 15107 32275 15113
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 27724 15048 28212 15076
rect 27709 15011 27767 15017
rect 27709 15008 27721 15011
rect 27540 14980 27721 15008
rect 27709 14977 27721 14980
rect 27755 14977 27767 15011
rect 27709 14971 27767 14977
rect 27798 14968 27804 15020
rect 27856 15008 27862 15020
rect 28184 15017 28212 15048
rect 27893 15011 27951 15017
rect 27893 15008 27905 15011
rect 27856 14980 27905 15008
rect 27856 14968 27862 14980
rect 27893 14977 27905 14980
rect 27939 14977 27951 15011
rect 27893 14971 27951 14977
rect 28169 15011 28227 15017
rect 28169 14977 28181 15011
rect 28215 14977 28227 15011
rect 28169 14971 28227 14977
rect 28353 15011 28411 15017
rect 28353 14977 28365 15011
rect 28399 14977 28411 15011
rect 29825 15011 29883 15017
rect 29825 15008 29837 15011
rect 28353 14971 28411 14977
rect 29656 14980 29837 15008
rect 27522 14940 27528 14952
rect 27448 14912 27528 14940
rect 27120 14900 27126 14912
rect 27522 14900 27528 14912
rect 27580 14940 27586 14952
rect 28077 14943 28135 14949
rect 28077 14940 28089 14943
rect 27580 14912 28089 14940
rect 27580 14900 27586 14912
rect 28077 14909 28089 14912
rect 28123 14940 28135 14943
rect 28368 14940 28396 14971
rect 28123 14912 28396 14940
rect 28123 14909 28135 14912
rect 28077 14903 28135 14909
rect 28994 14900 29000 14952
rect 29052 14900 29058 14952
rect 24259 14844 25084 14872
rect 24259 14841 24271 14844
rect 24213 14835 24271 14841
rect 26234 14832 26240 14884
rect 26292 14872 26298 14884
rect 26973 14875 27031 14881
rect 26973 14872 26985 14875
rect 26292 14844 26985 14872
rect 26292 14832 26298 14844
rect 26973 14841 26985 14844
rect 27019 14841 27031 14875
rect 29012 14872 29040 14900
rect 26973 14835 27031 14841
rect 27632 14844 29040 14872
rect 22097 14807 22166 14813
rect 22097 14773 22109 14807
rect 22143 14776 22166 14807
rect 22281 14807 22339 14813
rect 22143 14773 22155 14776
rect 22097 14767 22155 14773
rect 22281 14773 22293 14807
rect 22327 14804 22339 14807
rect 22370 14804 22376 14816
rect 22327 14776 22376 14804
rect 22327 14773 22339 14776
rect 22281 14767 22339 14773
rect 22370 14764 22376 14776
rect 22428 14764 22434 14816
rect 22462 14764 22468 14816
rect 22520 14764 22526 14816
rect 22922 14764 22928 14816
rect 22980 14764 22986 14816
rect 23014 14764 23020 14816
rect 23072 14764 23078 14816
rect 23106 14764 23112 14816
rect 23164 14804 23170 14816
rect 23201 14807 23259 14813
rect 23201 14804 23213 14807
rect 23164 14776 23213 14804
rect 23164 14764 23170 14776
rect 23201 14773 23213 14776
rect 23247 14773 23259 14807
rect 23201 14767 23259 14773
rect 25501 14807 25559 14813
rect 25501 14773 25513 14807
rect 25547 14804 25559 14807
rect 27632 14804 27660 14844
rect 25547 14776 27660 14804
rect 25547 14773 25559 14776
rect 25501 14767 25559 14773
rect 28258 14764 28264 14816
rect 28316 14764 28322 14816
rect 29454 14764 29460 14816
rect 29512 14804 29518 14816
rect 29656 14813 29684 14980
rect 29825 14977 29837 14980
rect 29871 15008 29883 15011
rect 30006 15008 30012 15020
rect 29871 14980 30012 15008
rect 29871 14977 29883 14980
rect 29825 14971 29883 14977
rect 30006 14968 30012 14980
rect 30064 15008 30070 15020
rect 30374 15008 30380 15020
rect 30064 14980 30380 15008
rect 30064 14968 30070 14980
rect 30374 14968 30380 14980
rect 30432 15008 30438 15020
rect 31202 15008 31208 15020
rect 30432 14980 31208 15008
rect 30432 14968 30438 14980
rect 31202 14968 31208 14980
rect 31260 14968 31266 15020
rect 31846 14968 31852 15020
rect 31904 15008 31910 15020
rect 32401 15011 32459 15017
rect 32401 15008 32413 15011
rect 31904 14980 32413 15008
rect 31904 14968 31910 14980
rect 32401 14977 32413 14980
rect 32447 15008 32459 15011
rect 32674 15008 32680 15020
rect 32447 14980 32680 15008
rect 32447 14977 32459 14980
rect 32401 14971 32459 14977
rect 32674 14968 32680 14980
rect 32732 14968 32738 15020
rect 29641 14807 29699 14813
rect 29641 14804 29653 14807
rect 29512 14776 29653 14804
rect 29512 14764 29518 14776
rect 29641 14773 29653 14776
rect 29687 14773 29699 14807
rect 29641 14767 29699 14773
rect 29914 14764 29920 14816
rect 29972 14764 29978 14816
rect 1104 14714 35248 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 35248 14714
rect 1104 14640 35248 14662
rect 4982 14560 4988 14612
rect 5040 14560 5046 14612
rect 5077 14603 5135 14609
rect 5077 14569 5089 14603
rect 5123 14600 5135 14603
rect 5166 14600 5172 14612
rect 5123 14572 5172 14600
rect 5123 14569 5135 14572
rect 5077 14563 5135 14569
rect 5166 14560 5172 14572
rect 5224 14560 5230 14612
rect 5258 14560 5264 14612
rect 5316 14560 5322 14612
rect 5350 14560 5356 14612
rect 5408 14560 5414 14612
rect 10689 14603 10747 14609
rect 10689 14569 10701 14603
rect 10735 14600 10747 14603
rect 11606 14600 11612 14612
rect 10735 14572 11612 14600
rect 10735 14569 10747 14572
rect 10689 14563 10747 14569
rect 11606 14560 11612 14572
rect 11664 14560 11670 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12621 14603 12679 14609
rect 12621 14600 12633 14603
rect 12032 14572 12633 14600
rect 12032 14560 12038 14572
rect 12621 14569 12633 14572
rect 12667 14600 12679 14603
rect 13630 14600 13636 14612
rect 12667 14572 13636 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 13909 14603 13967 14609
rect 13909 14569 13921 14603
rect 13955 14600 13967 14603
rect 14366 14600 14372 14612
rect 13955 14572 14372 14600
rect 13955 14569 13967 14572
rect 13909 14563 13967 14569
rect 14366 14560 14372 14572
rect 14424 14560 14430 14612
rect 14734 14560 14740 14612
rect 14792 14600 14798 14612
rect 16574 14600 16580 14612
rect 14792 14572 16580 14600
rect 14792 14560 14798 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 18874 14560 18880 14612
rect 18932 14560 18938 14612
rect 21174 14600 21180 14612
rect 20732 14572 21180 14600
rect 4341 14535 4399 14541
rect 4341 14501 4353 14535
rect 4387 14532 4399 14535
rect 5000 14532 5028 14560
rect 5368 14532 5396 14560
rect 4387 14504 5396 14532
rect 12989 14535 13047 14541
rect 4387 14501 4399 14504
rect 4341 14495 4399 14501
rect 12989 14501 13001 14535
rect 13035 14532 13047 14535
rect 13357 14535 13415 14541
rect 13357 14532 13369 14535
rect 13035 14504 13369 14532
rect 13035 14501 13047 14504
rect 12989 14495 13047 14501
rect 13357 14501 13369 14504
rect 13403 14532 13415 14535
rect 13446 14532 13452 14544
rect 13403 14504 13452 14532
rect 13403 14501 13415 14504
rect 13357 14495 13415 14501
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4356 14396 4384 14495
rect 13446 14492 13452 14504
rect 13504 14492 13510 14544
rect 13648 14532 13676 14560
rect 14553 14535 14611 14541
rect 14553 14532 14565 14535
rect 13648 14504 14565 14532
rect 14553 14501 14565 14504
rect 14599 14532 14611 14535
rect 14918 14532 14924 14544
rect 14599 14504 14924 14532
rect 14599 14501 14611 14504
rect 14553 14495 14611 14501
rect 14918 14492 14924 14504
rect 14976 14532 14982 14544
rect 15749 14535 15807 14541
rect 15749 14532 15761 14535
rect 14976 14504 15761 14532
rect 14976 14492 14982 14504
rect 15749 14501 15761 14504
rect 15795 14501 15807 14535
rect 15749 14495 15807 14501
rect 4985 14467 5043 14473
rect 4985 14433 4997 14467
rect 5031 14464 5043 14467
rect 5031 14436 5304 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 5276 14408 5304 14436
rect 5902 14424 5908 14476
rect 5960 14464 5966 14476
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 5960 14436 6561 14464
rect 5960 14424 5966 14436
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 8297 14467 8355 14473
rect 8297 14433 8309 14467
rect 8343 14464 8355 14467
rect 9217 14467 9275 14473
rect 9217 14464 9229 14467
rect 8343 14436 9229 14464
rect 8343 14433 8355 14436
rect 8297 14427 8355 14433
rect 9217 14433 9229 14436
rect 9263 14433 9275 14467
rect 15764 14464 15792 14495
rect 16669 14467 16727 14473
rect 16669 14464 16681 14467
rect 15764 14436 16681 14464
rect 9217 14427 9275 14433
rect 16669 14433 16681 14436
rect 16715 14464 16727 14467
rect 16758 14464 16764 14476
rect 16715 14436 16764 14464
rect 16715 14433 16727 14436
rect 16669 14427 16727 14433
rect 16758 14424 16764 14436
rect 16816 14464 16822 14476
rect 17586 14464 17592 14476
rect 16816 14436 17592 14464
rect 16816 14424 16822 14436
rect 4019 14368 4384 14396
rect 5077 14399 5135 14405
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 5077 14365 5089 14399
rect 5123 14365 5135 14399
rect 5077 14359 5135 14365
rect 4798 14288 4804 14340
rect 4856 14288 4862 14340
rect 5092 14328 5120 14359
rect 5258 14356 5264 14408
rect 5316 14356 5322 14408
rect 5534 14356 5540 14408
rect 5592 14356 5598 14408
rect 8570 14356 8576 14408
rect 8628 14356 8634 14408
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8812 14368 8953 14396
rect 8812 14356 8818 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 16853 14399 16911 14405
rect 16853 14396 16865 14399
rect 8941 14359 8999 14365
rect 15396 14368 16865 14396
rect 5552 14328 5580 14356
rect 5092 14300 5580 14328
rect 6825 14331 6883 14337
rect 6825 14297 6837 14331
rect 6871 14297 6883 14331
rect 8481 14331 8539 14337
rect 8481 14328 8493 14331
rect 8050 14300 8493 14328
rect 6825 14291 6883 14297
rect 8481 14297 8493 14300
rect 8527 14297 8539 14331
rect 8588 14328 8616 14356
rect 9122 14328 9128 14340
rect 8588 14300 9128 14328
rect 8481 14291 8539 14297
rect 3878 14220 3884 14272
rect 3936 14220 3942 14272
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5350 14260 5356 14272
rect 5132 14232 5356 14260
rect 5132 14220 5138 14232
rect 5350 14220 5356 14232
rect 5408 14260 5414 14272
rect 6546 14260 6552 14272
rect 5408 14232 6552 14260
rect 5408 14220 5414 14232
rect 6546 14220 6552 14232
rect 6604 14260 6610 14272
rect 6840 14260 6868 14291
rect 9122 14288 9128 14300
rect 9180 14288 9186 14340
rect 9766 14288 9772 14340
rect 9824 14288 9830 14340
rect 15396 14272 15424 14368
rect 16853 14365 16865 14368
rect 16899 14365 16911 14399
rect 16853 14359 16911 14365
rect 17218 14356 17224 14408
rect 17276 14356 17282 14408
rect 17420 14405 17448 14436
rect 17586 14424 17592 14436
rect 17644 14464 17650 14476
rect 17865 14467 17923 14473
rect 17865 14464 17877 14467
rect 17644 14436 17877 14464
rect 17644 14424 17650 14436
rect 17865 14433 17877 14436
rect 17911 14464 17923 14467
rect 18966 14464 18972 14476
rect 17911 14436 18972 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 18966 14424 18972 14436
rect 19024 14424 19030 14476
rect 20732 14464 20760 14572
rect 21174 14560 21180 14572
rect 21232 14600 21238 14612
rect 21361 14603 21419 14609
rect 21361 14600 21373 14603
rect 21232 14572 21373 14600
rect 21232 14560 21238 14572
rect 21361 14569 21373 14572
rect 21407 14569 21419 14603
rect 23937 14603 23995 14609
rect 21361 14563 21419 14569
rect 22112 14572 23796 14600
rect 20898 14492 20904 14544
rect 20956 14532 20962 14544
rect 22112 14532 22140 14572
rect 20956 14504 22140 14532
rect 22557 14535 22615 14541
rect 20956 14492 20962 14504
rect 22557 14501 22569 14535
rect 22603 14532 22615 14535
rect 22738 14532 22744 14544
rect 22603 14504 22744 14532
rect 22603 14501 22615 14504
rect 22557 14495 22615 14501
rect 22738 14492 22744 14504
rect 22796 14492 22802 14544
rect 23566 14532 23572 14544
rect 23308 14504 23572 14532
rect 20088 14436 20760 14464
rect 17405 14399 17463 14405
rect 17405 14365 17417 14399
rect 17451 14365 17463 14399
rect 17405 14359 17463 14365
rect 17236 14328 17264 14356
rect 17589 14331 17647 14337
rect 17589 14328 17601 14331
rect 16132 14300 17264 14328
rect 17420 14300 17601 14328
rect 6604 14232 6868 14260
rect 6604 14220 6610 14232
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 11517 14263 11575 14269
rect 11517 14260 11529 14263
rect 11204 14232 11529 14260
rect 11204 14220 11210 14232
rect 11517 14229 11529 14232
rect 11563 14229 11575 14263
rect 11517 14223 11575 14229
rect 15378 14220 15384 14272
rect 15436 14220 15442 14272
rect 15930 14220 15936 14272
rect 15988 14260 15994 14272
rect 16132 14269 16160 14300
rect 17420 14272 17448 14300
rect 17589 14297 17601 14300
rect 17635 14297 17647 14331
rect 20088 14328 20116 14436
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20622 14398 20628 14408
rect 20456 14396 20628 14398
rect 20211 14370 20628 14396
rect 20211 14368 20484 14370
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 20622 14356 20628 14370
rect 20680 14356 20686 14408
rect 20732 14405 20760 14436
rect 20809 14467 20867 14473
rect 20809 14433 20821 14467
rect 20855 14464 20867 14467
rect 21729 14467 21787 14473
rect 21729 14464 21741 14467
rect 20855 14436 21741 14464
rect 20855 14433 20867 14436
rect 20809 14427 20867 14433
rect 21729 14433 21741 14436
rect 21775 14433 21787 14467
rect 21729 14427 21787 14433
rect 22649 14467 22707 14473
rect 22649 14433 22661 14467
rect 22695 14464 22707 14467
rect 22922 14464 22928 14476
rect 22695 14436 22928 14464
rect 22695 14433 22707 14436
rect 22649 14427 22707 14433
rect 22922 14424 22928 14436
rect 22980 14424 22986 14476
rect 23017 14467 23075 14473
rect 23017 14433 23029 14467
rect 23063 14433 23075 14467
rect 23017 14427 23075 14433
rect 20717 14399 20775 14405
rect 20717 14365 20729 14399
rect 20763 14365 20775 14399
rect 20717 14359 20775 14365
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 20257 14331 20315 14337
rect 20257 14328 20269 14331
rect 20088 14300 20269 14328
rect 17589 14291 17647 14297
rect 20257 14297 20269 14300
rect 20303 14297 20315 14331
rect 20257 14291 20315 14297
rect 20438 14288 20444 14340
rect 20496 14288 20502 14340
rect 20640 14328 20668 14356
rect 21008 14328 21036 14359
rect 21266 14356 21272 14408
rect 21324 14396 21330 14408
rect 21361 14399 21419 14405
rect 21361 14396 21373 14399
rect 21324 14368 21373 14396
rect 21324 14356 21330 14368
rect 21361 14365 21373 14368
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21545 14399 21603 14405
rect 21545 14365 21557 14399
rect 21591 14396 21603 14399
rect 21818 14396 21824 14408
rect 21591 14368 21824 14396
rect 21591 14365 21603 14368
rect 21545 14359 21603 14365
rect 21560 14328 21588 14359
rect 21818 14356 21824 14368
rect 21876 14356 21882 14408
rect 22278 14356 22284 14408
rect 22336 14396 22342 14408
rect 22336 14368 22508 14396
rect 22336 14356 22342 14368
rect 20640 14300 21036 14328
rect 21100 14300 21588 14328
rect 16117 14263 16175 14269
rect 16117 14260 16129 14263
rect 15988 14232 16129 14260
rect 15988 14220 15994 14232
rect 16117 14229 16129 14232
rect 16163 14229 16175 14263
rect 16117 14223 16175 14229
rect 17034 14220 17040 14272
rect 17092 14220 17098 14272
rect 17402 14220 17408 14272
rect 17460 14220 17466 14272
rect 18966 14220 18972 14272
rect 19024 14260 19030 14272
rect 19334 14260 19340 14272
rect 19024 14232 19340 14260
rect 19024 14220 19030 14232
rect 19334 14220 19340 14232
rect 19392 14260 19398 14272
rect 19429 14263 19487 14269
rect 19429 14260 19441 14263
rect 19392 14232 19441 14260
rect 19392 14220 19398 14232
rect 19429 14229 19441 14232
rect 19475 14229 19487 14263
rect 19429 14223 19487 14229
rect 20070 14220 20076 14272
rect 20128 14220 20134 14272
rect 20346 14269 20352 14272
rect 20342 14223 20352 14269
rect 20346 14220 20352 14223
rect 20404 14220 20410 14272
rect 20530 14220 20536 14272
rect 20588 14220 20594 14272
rect 20806 14220 20812 14272
rect 20864 14260 20870 14272
rect 21100 14260 21128 14300
rect 20864 14232 21128 14260
rect 20864 14220 20870 14232
rect 21174 14220 21180 14272
rect 21232 14220 21238 14272
rect 21266 14220 21272 14272
rect 21324 14260 21330 14272
rect 22097 14263 22155 14269
rect 22097 14260 22109 14263
rect 21324 14232 22109 14260
rect 21324 14220 21330 14232
rect 22097 14229 22109 14232
rect 22143 14229 22155 14263
rect 22097 14223 22155 14229
rect 22370 14220 22376 14272
rect 22428 14220 22434 14272
rect 22480 14260 22508 14368
rect 22557 14331 22615 14337
rect 22557 14297 22569 14331
rect 22603 14328 22615 14331
rect 22922 14328 22928 14340
rect 22603 14300 22928 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 22922 14288 22928 14300
rect 22980 14288 22986 14340
rect 23032 14328 23060 14427
rect 23106 14356 23112 14408
rect 23164 14356 23170 14408
rect 23198 14356 23204 14408
rect 23256 14396 23262 14408
rect 23308 14396 23336 14504
rect 23566 14492 23572 14504
rect 23624 14492 23630 14544
rect 23768 14532 23796 14572
rect 23937 14569 23949 14603
rect 23983 14600 23995 14603
rect 24302 14600 24308 14612
rect 23983 14572 24308 14600
rect 23983 14569 23995 14572
rect 23937 14563 23995 14569
rect 24302 14560 24308 14572
rect 24360 14560 24366 14612
rect 24412 14572 26556 14600
rect 24412 14532 24440 14572
rect 26528 14544 26556 14572
rect 26602 14560 26608 14612
rect 26660 14600 26666 14612
rect 31846 14600 31852 14612
rect 26660 14572 31852 14600
rect 26660 14560 26666 14572
rect 31846 14560 31852 14572
rect 31904 14600 31910 14612
rect 32125 14603 32183 14609
rect 32125 14600 32137 14603
rect 31904 14572 32137 14600
rect 31904 14560 31910 14572
rect 32125 14569 32137 14572
rect 32171 14569 32183 14603
rect 32125 14563 32183 14569
rect 32953 14603 33011 14609
rect 32953 14569 32965 14603
rect 32999 14600 33011 14603
rect 33042 14600 33048 14612
rect 32999 14572 33048 14600
rect 32999 14569 33011 14572
rect 32953 14563 33011 14569
rect 23768 14504 24440 14532
rect 26510 14492 26516 14544
rect 26568 14492 26574 14544
rect 26786 14492 26792 14544
rect 26844 14532 26850 14544
rect 26844 14504 27200 14532
rect 26844 14492 26850 14504
rect 26973 14467 27031 14473
rect 26973 14433 26985 14467
rect 27019 14464 27031 14467
rect 27062 14464 27068 14476
rect 27019 14436 27068 14464
rect 27019 14433 27031 14436
rect 26973 14427 27031 14433
rect 27062 14424 27068 14436
rect 27120 14424 27126 14476
rect 23385 14399 23443 14405
rect 23385 14396 23397 14399
rect 23256 14368 23397 14396
rect 23256 14356 23262 14368
rect 23385 14365 23397 14368
rect 23431 14365 23443 14399
rect 23385 14359 23443 14365
rect 23474 14356 23480 14408
rect 23532 14356 23538 14408
rect 23658 14356 23664 14408
rect 23716 14356 23722 14408
rect 23750 14356 23756 14408
rect 23808 14356 23814 14408
rect 25498 14356 25504 14408
rect 25556 14356 25562 14408
rect 27172 14405 27200 14504
rect 28258 14492 28264 14544
rect 28316 14492 28322 14544
rect 29270 14492 29276 14544
rect 29328 14532 29334 14544
rect 32968 14532 32996 14563
rect 33042 14560 33048 14572
rect 33100 14560 33106 14612
rect 29328 14504 29592 14532
rect 29328 14492 29334 14504
rect 28077 14467 28135 14473
rect 28077 14433 28089 14467
rect 28123 14464 28135 14467
rect 28276 14464 28304 14492
rect 29564 14473 29592 14504
rect 30852 14504 32996 14532
rect 28123 14436 28304 14464
rect 29549 14467 29607 14473
rect 28123 14433 28135 14436
rect 28077 14427 28135 14433
rect 29549 14433 29561 14467
rect 29595 14464 29607 14467
rect 30852 14464 30880 14504
rect 31665 14467 31723 14473
rect 31665 14464 31677 14467
rect 29595 14436 30880 14464
rect 31312 14436 31677 14464
rect 29595 14433 29607 14436
rect 29549 14427 29607 14433
rect 31312 14408 31340 14436
rect 31665 14433 31677 14436
rect 31711 14433 31723 14467
rect 31665 14427 31723 14433
rect 31846 14424 31852 14476
rect 31904 14424 31910 14476
rect 34057 14467 34115 14473
rect 34057 14433 34069 14467
rect 34103 14464 34115 14467
rect 34103 14436 34652 14464
rect 34103 14433 34115 14436
rect 34057 14427 34115 14433
rect 25777 14399 25835 14405
rect 25777 14396 25789 14399
rect 25700 14368 25789 14396
rect 23676 14328 23704 14356
rect 23032 14300 23704 14328
rect 24578 14288 24584 14340
rect 24636 14288 24642 14340
rect 22830 14260 22836 14272
rect 22480 14232 22836 14260
rect 22830 14220 22836 14232
rect 22888 14220 22894 14272
rect 23293 14263 23351 14269
rect 23293 14229 23305 14263
rect 23339 14260 23351 14263
rect 24596 14260 24624 14288
rect 25700 14269 25728 14368
rect 25777 14365 25789 14368
rect 25823 14365 25835 14399
rect 25777 14359 25835 14365
rect 27157 14399 27215 14405
rect 27157 14365 27169 14399
rect 27203 14365 27215 14399
rect 27157 14359 27215 14365
rect 27982 14356 27988 14408
rect 28040 14356 28046 14408
rect 28166 14356 28172 14408
rect 28224 14396 28230 14408
rect 29454 14396 29460 14408
rect 28224 14368 29460 14396
rect 28224 14356 28230 14368
rect 29454 14356 29460 14368
rect 29512 14356 29518 14408
rect 31294 14356 31300 14408
rect 31352 14356 31358 14408
rect 31573 14399 31631 14405
rect 31573 14365 31585 14399
rect 31619 14365 31631 14399
rect 31573 14359 31631 14365
rect 34517 14399 34575 14405
rect 34517 14365 34529 14399
rect 34563 14365 34575 14399
rect 34517 14359 34575 14365
rect 29825 14331 29883 14337
rect 29825 14328 29837 14331
rect 28368 14300 29837 14328
rect 23339 14232 24624 14260
rect 25685 14263 25743 14269
rect 23339 14229 23351 14232
rect 23293 14223 23351 14229
rect 25685 14229 25697 14263
rect 25731 14229 25743 14263
rect 25685 14223 25743 14229
rect 25961 14263 26019 14269
rect 25961 14229 25973 14263
rect 26007 14260 26019 14263
rect 26418 14260 26424 14272
rect 26007 14232 26424 14260
rect 26007 14229 26019 14232
rect 25961 14223 26019 14229
rect 26418 14220 26424 14232
rect 26476 14220 26482 14272
rect 27341 14263 27399 14269
rect 27341 14229 27353 14263
rect 27387 14260 27399 14263
rect 27430 14260 27436 14272
rect 27387 14232 27436 14260
rect 27387 14229 27399 14232
rect 27341 14223 27399 14229
rect 27430 14220 27436 14232
rect 27488 14220 27494 14272
rect 28368 14269 28396 14300
rect 29825 14297 29837 14300
rect 29871 14297 29883 14331
rect 29825 14291 29883 14297
rect 29914 14288 29920 14340
rect 29972 14328 29978 14340
rect 31588 14328 31616 14359
rect 29972 14300 30314 14328
rect 31588 14300 31800 14328
rect 29972 14288 29978 14300
rect 31772 14272 31800 14300
rect 28353 14263 28411 14269
rect 28353 14229 28365 14263
rect 28399 14229 28411 14263
rect 28353 14223 28411 14229
rect 31297 14263 31355 14269
rect 31297 14229 31309 14263
rect 31343 14260 31355 14263
rect 31754 14260 31760 14272
rect 31343 14232 31760 14260
rect 31343 14229 31355 14232
rect 31297 14223 31355 14229
rect 31754 14220 31760 14232
rect 31812 14220 31818 14272
rect 31849 14263 31907 14269
rect 31849 14229 31861 14263
rect 31895 14260 31907 14263
rect 32214 14260 32220 14272
rect 31895 14232 32220 14260
rect 31895 14229 31907 14232
rect 31849 14223 31907 14229
rect 32214 14220 32220 14232
rect 32272 14220 32278 14272
rect 34532 14260 34560 14359
rect 34624 14340 34652 14436
rect 34606 14288 34612 14340
rect 34664 14288 34670 14340
rect 34532 14232 35296 14260
rect 1104 14170 35236 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 35236 14170
rect 1104 14096 35236 14118
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 4798 14056 4804 14068
rect 4387 14028 4804 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 5166 14016 5172 14068
rect 5224 14056 5230 14068
rect 5224 14028 6776 14056
rect 5224 14016 5230 14028
rect 2866 13948 2872 14000
rect 2924 13948 2930 14000
rect 3878 13948 3884 14000
rect 3936 13948 3942 14000
rect 5534 13988 5540 14000
rect 5092 13960 5540 13988
rect 5092 13929 5120 13960
rect 5534 13948 5540 13960
rect 5592 13988 5598 14000
rect 5592 13960 6684 13988
rect 5592 13948 5598 13960
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13889 5135 13923
rect 5077 13883 5135 13889
rect 2608 13852 2636 13883
rect 5350 13880 5356 13932
rect 5408 13880 5414 13932
rect 5721 13923 5779 13929
rect 5721 13918 5733 13923
rect 5644 13890 5733 13918
rect 3510 13852 3516 13864
rect 2608 13824 3516 13852
rect 3510 13812 3516 13824
rect 3568 13852 3574 13864
rect 4617 13855 4675 13861
rect 4617 13852 4629 13855
rect 3568 13824 4629 13852
rect 3568 13812 3574 13824
rect 4617 13821 4629 13824
rect 4663 13821 4675 13855
rect 5644 13852 5672 13890
rect 5721 13889 5733 13890
rect 5767 13889 5779 13923
rect 5721 13883 5779 13889
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 4617 13815 4675 13821
rect 5276 13824 5672 13852
rect 5813 13855 5871 13861
rect 5276 13796 5304 13824
rect 5813 13821 5825 13855
rect 5859 13852 5871 13855
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 5859 13824 6377 13852
rect 5859 13821 5871 13824
rect 5813 13815 5871 13821
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 6656 13852 6684 13960
rect 6748 13929 6776 14028
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8812 14028 9045 14056
rect 8812 14016 8818 14028
rect 9033 14025 9045 14028
rect 9079 14056 9091 14059
rect 9079 14028 9674 14056
rect 9079 14025 9091 14028
rect 9033 14019 9091 14025
rect 6733 13923 6791 13929
rect 6733 13889 6745 13923
rect 6779 13889 6791 13923
rect 6733 13883 6791 13889
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 6840 13852 6868 13883
rect 6656 13824 6868 13852
rect 9646 13852 9674 14028
rect 9766 14016 9772 14068
rect 9824 14016 9830 14068
rect 10229 14059 10287 14065
rect 10229 14025 10241 14059
rect 10275 14056 10287 14059
rect 10502 14056 10508 14068
rect 10275 14028 10508 14056
rect 10275 14025 10287 14028
rect 10229 14019 10287 14025
rect 9861 13923 9919 13929
rect 9861 13889 9873 13923
rect 9907 13920 9919 13923
rect 10244 13920 10272 14019
rect 10502 14016 10508 14028
rect 10560 14016 10566 14068
rect 11514 14016 11520 14068
rect 11572 14056 11578 14068
rect 13538 14056 13544 14068
rect 11572 14028 13544 14056
rect 11572 14016 11578 14028
rect 13538 14016 13544 14028
rect 13596 14056 13602 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13596 14028 13645 14056
rect 13596 14016 13602 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 14550 14016 14556 14068
rect 14608 14056 14614 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14608 14028 14749 14056
rect 14608 14016 14614 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 14752 13988 14780 14019
rect 16114 14016 16120 14068
rect 16172 14056 16178 14068
rect 20438 14056 20444 14068
rect 16172 14028 20444 14056
rect 16172 14016 16178 14028
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 21174 14016 21180 14068
rect 21232 14016 21238 14068
rect 21266 14016 21272 14068
rect 21324 14016 21330 14068
rect 21818 14016 21824 14068
rect 21876 14016 21882 14068
rect 23109 14059 23167 14065
rect 23109 14025 23121 14059
rect 23155 14056 23167 14059
rect 23382 14056 23388 14068
rect 23155 14028 23388 14056
rect 23155 14025 23167 14028
rect 23109 14019 23167 14025
rect 23382 14016 23388 14028
rect 23440 14056 23446 14068
rect 23750 14056 23756 14068
rect 23440 14028 23756 14056
rect 23440 14016 23446 14028
rect 23750 14016 23756 14028
rect 23808 14016 23814 14068
rect 25133 14059 25191 14065
rect 25133 14025 25145 14059
rect 25179 14056 25191 14059
rect 25498 14056 25504 14068
rect 25179 14028 25504 14056
rect 25179 14025 25191 14028
rect 25133 14019 25191 14025
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 26142 14056 26148 14068
rect 25608 14028 26148 14056
rect 17037 13991 17095 13997
rect 14752 13960 16988 13988
rect 9907 13892 10272 13920
rect 9907 13889 9919 13892
rect 9861 13883 9919 13889
rect 11146 13880 11152 13932
rect 11204 13880 11210 13932
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 15378 13920 15384 13932
rect 14691 13892 15384 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 11164 13852 11192 13880
rect 9646 13824 11192 13852
rect 6365 13815 6423 13821
rect 12802 13812 12808 13864
rect 12860 13812 12866 13864
rect 14093 13855 14151 13861
rect 14093 13821 14105 13855
rect 14139 13852 14151 13855
rect 14660 13852 14688 13883
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 15933 13923 15991 13929
rect 15933 13920 15945 13923
rect 15580 13892 15945 13920
rect 14139 13824 14688 13852
rect 14139 13821 14151 13824
rect 14093 13815 14151 13821
rect 5166 13744 5172 13796
rect 5224 13744 5230 13796
rect 5258 13744 5264 13796
rect 5316 13744 5322 13796
rect 6089 13787 6147 13793
rect 6089 13753 6101 13787
rect 6135 13784 6147 13787
rect 6914 13784 6920 13796
rect 6135 13756 6920 13784
rect 6135 13753 6147 13756
rect 6089 13747 6147 13753
rect 6914 13744 6920 13756
rect 6972 13744 6978 13796
rect 12894 13744 12900 13796
rect 12952 13784 12958 13796
rect 14108 13784 14136 13815
rect 12952 13756 14136 13784
rect 12952 13744 12958 13756
rect 14918 13744 14924 13796
rect 14976 13784 14982 13796
rect 15580 13793 15608 13892
rect 15933 13889 15945 13892
rect 15979 13920 15991 13923
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 15979 13892 16681 13920
rect 15979 13889 15991 13892
rect 15933 13883 15991 13889
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16850 13880 16856 13932
rect 16908 13880 16914 13932
rect 15749 13855 15807 13861
rect 15749 13821 15761 13855
rect 15795 13852 15807 13855
rect 15838 13852 15844 13864
rect 15795 13824 15844 13852
rect 15795 13821 15807 13824
rect 15749 13815 15807 13821
rect 15197 13787 15255 13793
rect 15197 13784 15209 13787
rect 14976 13756 15209 13784
rect 14976 13744 14982 13756
rect 15197 13753 15209 13756
rect 15243 13784 15255 13787
rect 15565 13787 15623 13793
rect 15565 13784 15577 13787
rect 15243 13756 15577 13784
rect 15243 13753 15255 13756
rect 15197 13747 15255 13753
rect 15565 13753 15577 13756
rect 15611 13753 15623 13787
rect 15565 13747 15623 13753
rect 4890 13676 4896 13728
rect 4948 13676 4954 13728
rect 8757 13719 8815 13725
rect 8757 13685 8769 13719
rect 8803 13716 8815 13719
rect 9122 13716 9128 13728
rect 8803 13688 9128 13716
rect 8803 13685 8815 13688
rect 8757 13679 8815 13685
rect 9122 13676 9128 13688
rect 9180 13676 9186 13728
rect 14182 13676 14188 13728
rect 14240 13716 14246 13728
rect 14553 13719 14611 13725
rect 14553 13716 14565 13719
rect 14240 13688 14565 13716
rect 14240 13676 14246 13688
rect 14553 13685 14565 13688
rect 14599 13716 14611 13719
rect 15764 13716 15792 13815
rect 15838 13812 15844 13824
rect 15896 13812 15902 13864
rect 16960 13852 16988 13960
rect 17037 13957 17049 13991
rect 17083 13988 17095 13991
rect 20070 13988 20076 14000
rect 17083 13960 17632 13988
rect 17083 13957 17095 13960
rect 17037 13951 17095 13957
rect 17402 13880 17408 13932
rect 17460 13880 17466 13932
rect 17604 13929 17632 13960
rect 19352 13960 19840 13988
rect 19352 13932 19380 13960
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 17736 13892 18920 13920
rect 17736 13880 17742 13892
rect 18892 13864 18920 13892
rect 19242 13880 19248 13932
rect 19300 13880 19306 13932
rect 19334 13880 19340 13932
rect 19392 13880 19398 13932
rect 19426 13880 19432 13932
rect 19484 13880 19490 13932
rect 19812 13929 19840 13960
rect 19904 13960 20076 13988
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13889 19855 13923
rect 19797 13883 19855 13889
rect 16960 13824 17264 13852
rect 17236 13784 17264 13824
rect 18874 13812 18880 13864
rect 18932 13852 18938 13864
rect 19518 13852 19524 13864
rect 18932 13824 19524 13852
rect 18932 13812 18938 13824
rect 19518 13812 19524 13824
rect 19576 13812 19582 13864
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13852 19671 13855
rect 19904 13852 19932 13960
rect 20070 13948 20076 13960
rect 20128 13948 20134 14000
rect 21082 13988 21088 14000
rect 20732 13960 21088 13988
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13920 20039 13923
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 20027 13892 20361 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13920 20499 13923
rect 20530 13920 20536 13932
rect 20487 13892 20536 13920
rect 20487 13889 20499 13892
rect 20441 13883 20499 13889
rect 20530 13880 20536 13892
rect 20588 13880 20594 13932
rect 20732 13929 20760 13960
rect 21082 13948 21088 13960
rect 21140 13948 21146 14000
rect 20717 13923 20775 13929
rect 20717 13889 20729 13923
rect 20763 13889 20775 13923
rect 20717 13883 20775 13889
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13920 21051 13923
rect 21192 13920 21220 14016
rect 21039 13892 21220 13920
rect 21284 13920 21312 14016
rect 21836 13988 21864 14016
rect 22005 13991 22063 13997
rect 22005 13988 22017 13991
rect 21836 13960 22017 13988
rect 22005 13957 22017 13960
rect 22051 13957 22063 13991
rect 22005 13951 22063 13957
rect 22370 13948 22376 14000
rect 22428 13988 22434 14000
rect 22741 13991 22799 13997
rect 22741 13988 22753 13991
rect 22428 13960 22753 13988
rect 22428 13948 22434 13960
rect 22741 13957 22753 13960
rect 22787 13957 22799 13991
rect 22741 13951 22799 13957
rect 22971 13957 23029 13963
rect 22971 13954 22983 13957
rect 22956 13932 22983 13954
rect 21542 13920 21548 13932
rect 21284 13892 21548 13920
rect 21039 13889 21051 13892
rect 20993 13883 21051 13889
rect 21542 13880 21548 13892
rect 21600 13880 21606 13932
rect 22922 13880 22928 13932
rect 22980 13923 22983 13932
rect 23017 13923 23029 13957
rect 25222 13948 25228 14000
rect 25280 13948 25286 14000
rect 25608 13988 25636 14028
rect 26142 14016 26148 14028
rect 26200 14016 26206 14068
rect 26234 14016 26240 14068
rect 26292 14016 26298 14068
rect 26326 14016 26332 14068
rect 26384 14016 26390 14068
rect 26418 14016 26424 14068
rect 26476 14016 26482 14068
rect 26513 14059 26571 14065
rect 26513 14025 26525 14059
rect 26559 14025 26571 14059
rect 26513 14019 26571 14025
rect 25332 13960 25636 13988
rect 25700 13960 26004 13988
rect 22980 13917 23029 13923
rect 24949 13923 25007 13929
rect 22980 13880 22986 13917
rect 24949 13889 24961 13923
rect 24995 13920 25007 13923
rect 25332 13920 25360 13960
rect 24995 13892 25360 13920
rect 25409 13923 25467 13929
rect 24995 13889 25007 13892
rect 24949 13883 25007 13889
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25501 13923 25559 13929
rect 25501 13889 25513 13923
rect 25547 13920 25559 13923
rect 25590 13920 25596 13932
rect 25547 13892 25596 13920
rect 25547 13889 25559 13892
rect 25501 13883 25559 13889
rect 19659 13824 19932 13852
rect 20165 13855 20223 13861
rect 19659 13821 19671 13824
rect 19613 13815 19671 13821
rect 20165 13821 20177 13855
rect 20211 13852 20223 13855
rect 20625 13855 20683 13861
rect 20211 13824 20576 13852
rect 20211 13821 20223 13824
rect 20165 13815 20223 13821
rect 17236 13756 18368 13784
rect 14599 13688 15792 13716
rect 18340 13716 18368 13756
rect 18414 13744 18420 13796
rect 18472 13744 18478 13796
rect 19334 13744 19340 13796
rect 19392 13784 19398 13796
rect 19628 13784 19656 13815
rect 19392 13756 19656 13784
rect 19392 13744 19398 13756
rect 20346 13744 20352 13796
rect 20404 13744 20410 13796
rect 20548 13784 20576 13824
rect 20625 13821 20637 13855
rect 20671 13852 20683 13855
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 20671 13824 20821 13852
rect 20671 13821 20683 13824
rect 20625 13815 20683 13821
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20809 13815 20867 13821
rect 21266 13812 21272 13864
rect 21324 13852 21330 13864
rect 21453 13855 21511 13861
rect 21453 13852 21465 13855
rect 21324 13824 21465 13852
rect 21324 13812 21330 13824
rect 21453 13821 21465 13824
rect 21499 13821 21511 13855
rect 25222 13852 25228 13864
rect 21453 13815 21511 13821
rect 21560 13824 25228 13852
rect 21560 13784 21588 13824
rect 25222 13812 25228 13824
rect 25280 13812 25286 13864
rect 25424 13852 25452 13883
rect 25590 13880 25596 13892
rect 25648 13880 25654 13932
rect 25700 13929 25728 13960
rect 25685 13923 25743 13929
rect 25685 13889 25697 13923
rect 25731 13889 25743 13923
rect 25685 13883 25743 13889
rect 25774 13880 25780 13932
rect 25832 13880 25838 13932
rect 25869 13855 25927 13861
rect 25869 13852 25881 13855
rect 25424 13824 25881 13852
rect 25869 13821 25881 13824
rect 25915 13821 25927 13855
rect 25976 13852 26004 13960
rect 26050 13880 26056 13932
rect 26108 13880 26114 13932
rect 26252 13929 26280 14016
rect 26344 13929 26372 14016
rect 26237 13923 26295 13929
rect 26237 13889 26249 13923
rect 26283 13889 26295 13923
rect 26237 13883 26295 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13889 26387 13923
rect 26436 13920 26464 14016
rect 26528 13988 26556 14019
rect 27246 14016 27252 14068
rect 27304 14056 27310 14068
rect 27304 14028 27936 14056
rect 27304 14016 27310 14028
rect 26528 13960 26832 13988
rect 26697 13923 26755 13929
rect 26697 13920 26709 13923
rect 26436 13892 26709 13920
rect 26329 13883 26387 13889
rect 26697 13889 26709 13892
rect 26743 13889 26755 13923
rect 26697 13883 26755 13889
rect 26804 13852 26832 13960
rect 27172 13960 27752 13988
rect 27172 13929 27200 13960
rect 27157 13923 27215 13929
rect 27157 13889 27169 13923
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 27433 13923 27491 13929
rect 27433 13889 27445 13923
rect 27479 13920 27491 13923
rect 27522 13920 27528 13932
rect 27479 13892 27528 13920
rect 27479 13889 27491 13892
rect 27433 13883 27491 13889
rect 25976 13824 26832 13852
rect 25869 13815 25927 13821
rect 20548 13756 21588 13784
rect 25498 13744 25504 13796
rect 25556 13784 25562 13796
rect 26145 13787 26203 13793
rect 26145 13784 26157 13787
rect 25556 13756 26157 13784
rect 25556 13744 25562 13756
rect 26145 13753 26157 13756
rect 26191 13753 26203 13787
rect 26145 13747 26203 13753
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 27172 13784 27200 13883
rect 27522 13880 27528 13892
rect 27580 13880 27586 13932
rect 27724 13929 27752 13960
rect 27908 13929 27936 14028
rect 27982 14016 27988 14068
rect 28040 14016 28046 14068
rect 29270 14016 29276 14068
rect 29328 14016 29334 14068
rect 34793 14059 34851 14065
rect 34793 14025 34805 14059
rect 34839 14056 34851 14059
rect 35268 14056 35296 14232
rect 34839 14028 35296 14056
rect 34839 14025 34851 14028
rect 34793 14019 34851 14025
rect 27617 13923 27675 13929
rect 27617 13889 27629 13923
rect 27663 13889 27675 13923
rect 27617 13883 27675 13889
rect 27709 13923 27767 13929
rect 27709 13889 27721 13923
rect 27755 13889 27767 13923
rect 27709 13883 27767 13889
rect 27893 13923 27951 13929
rect 27893 13889 27905 13923
rect 27939 13889 27951 13923
rect 27893 13883 27951 13889
rect 27632 13852 27660 13883
rect 27448 13824 27660 13852
rect 27801 13855 27859 13861
rect 27448 13796 27476 13824
rect 27801 13821 27813 13855
rect 27847 13852 27859 13855
rect 28000 13852 28028 14016
rect 29288 13920 29316 14016
rect 30466 13948 30472 14000
rect 30524 13948 30530 14000
rect 31754 13988 31760 14000
rect 31588 13960 31760 13988
rect 31588 13929 31616 13960
rect 31754 13948 31760 13960
rect 31812 13948 31818 14000
rect 34054 13948 34060 14000
rect 34112 13948 34118 14000
rect 29457 13923 29515 13929
rect 29457 13920 29469 13923
rect 29288 13892 29469 13920
rect 29457 13889 29469 13892
rect 29503 13889 29515 13923
rect 31481 13923 31539 13929
rect 31481 13920 31493 13923
rect 29457 13883 29515 13889
rect 31312 13892 31493 13920
rect 27847 13824 28028 13852
rect 27847 13821 27859 13824
rect 27801 13815 27859 13821
rect 31312 13796 31340 13892
rect 31481 13889 31493 13892
rect 31527 13889 31539 13923
rect 31481 13883 31539 13889
rect 31573 13923 31631 13929
rect 31573 13889 31585 13923
rect 31619 13889 31631 13923
rect 32309 13923 32367 13929
rect 32309 13920 32321 13923
rect 31573 13883 31631 13889
rect 31726 13892 32321 13920
rect 26292 13756 27200 13784
rect 26292 13744 26298 13756
rect 27246 13744 27252 13796
rect 27304 13744 27310 13796
rect 27341 13787 27399 13793
rect 27341 13753 27353 13787
rect 27387 13753 27399 13787
rect 27341 13747 27399 13753
rect 18782 13716 18788 13728
rect 18340 13688 18788 13716
rect 14599 13685 14611 13688
rect 14553 13679 14611 13685
rect 18782 13676 18788 13688
rect 18840 13676 18846 13728
rect 20364 13716 20392 13744
rect 21177 13719 21235 13725
rect 21177 13716 21189 13719
rect 20364 13688 21189 13716
rect 21177 13685 21189 13688
rect 21223 13685 21235 13719
rect 21177 13679 21235 13685
rect 22830 13676 22836 13728
rect 22888 13716 22894 13728
rect 22925 13719 22983 13725
rect 22925 13716 22937 13719
rect 22888 13688 22937 13716
rect 22888 13676 22894 13688
rect 22925 13685 22937 13688
rect 22971 13685 22983 13719
rect 22925 13679 22983 13685
rect 25774 13676 25780 13728
rect 25832 13716 25838 13728
rect 26973 13719 27031 13725
rect 26973 13716 26985 13719
rect 25832 13688 26985 13716
rect 25832 13676 25838 13688
rect 26973 13685 26985 13688
rect 27019 13685 27031 13719
rect 27356 13716 27384 13747
rect 27430 13744 27436 13796
rect 27488 13744 27494 13796
rect 27614 13744 27620 13796
rect 27672 13744 27678 13796
rect 31294 13744 31300 13796
rect 31352 13744 31358 13796
rect 27632 13716 27660 13744
rect 27356 13688 27660 13716
rect 26973 13679 27031 13685
rect 29362 13676 29368 13728
rect 29420 13716 29426 13728
rect 29714 13719 29772 13725
rect 29714 13716 29726 13719
rect 29420 13688 29726 13716
rect 29420 13676 29426 13688
rect 29714 13685 29726 13688
rect 29760 13685 29772 13719
rect 29714 13679 29772 13685
rect 31205 13719 31263 13725
rect 31205 13685 31217 13719
rect 31251 13716 31263 13719
rect 31481 13719 31539 13725
rect 31481 13716 31493 13719
rect 31251 13688 31493 13716
rect 31251 13685 31263 13688
rect 31205 13679 31263 13685
rect 31481 13685 31493 13688
rect 31527 13716 31539 13719
rect 31726 13716 31754 13892
rect 32309 13889 32321 13892
rect 32355 13889 32367 13923
rect 32309 13883 32367 13889
rect 33042 13880 33048 13932
rect 33100 13880 33106 13932
rect 32214 13812 32220 13864
rect 32272 13812 32278 13864
rect 31849 13787 31907 13793
rect 31849 13753 31861 13787
rect 31895 13784 31907 13787
rect 31938 13784 31944 13796
rect 31895 13756 31944 13784
rect 31895 13753 31907 13756
rect 31849 13747 31907 13753
rect 31938 13744 31944 13756
rect 31996 13744 32002 13796
rect 31527 13688 31754 13716
rect 32585 13719 32643 13725
rect 31527 13685 31539 13688
rect 31481 13679 31539 13685
rect 32585 13685 32597 13719
rect 32631 13716 32643 13719
rect 33302 13719 33360 13725
rect 33302 13716 33314 13719
rect 32631 13688 33314 13716
rect 32631 13685 32643 13688
rect 32585 13679 32643 13685
rect 33302 13685 33314 13688
rect 33348 13685 33360 13719
rect 33302 13679 33360 13685
rect 1104 13626 35248 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 35248 13626
rect 1104 13552 35248 13574
rect 3145 13515 3203 13521
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 4614 13512 4620 13524
rect 3191 13484 4620 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 4798 13472 4804 13524
rect 4856 13472 4862 13524
rect 6914 13472 6920 13524
rect 6972 13472 6978 13524
rect 12161 13515 12219 13521
rect 12161 13481 12173 13515
rect 12207 13512 12219 13515
rect 12434 13512 12440 13524
rect 12207 13484 12440 13512
rect 12207 13481 12219 13484
rect 12161 13475 12219 13481
rect 12434 13472 12440 13484
rect 12492 13472 12498 13524
rect 13538 13472 13544 13524
rect 13596 13472 13602 13524
rect 13814 13472 13820 13524
rect 13872 13472 13878 13524
rect 15378 13472 15384 13524
rect 15436 13512 15442 13524
rect 15746 13512 15752 13524
rect 15436 13484 15752 13512
rect 15436 13472 15442 13484
rect 15746 13472 15752 13484
rect 15804 13512 15810 13524
rect 16206 13512 16212 13524
rect 15804 13484 16212 13512
rect 15804 13472 15810 13484
rect 16206 13472 16212 13484
rect 16264 13512 16270 13524
rect 18693 13515 18751 13521
rect 18693 13512 18705 13515
rect 16264 13484 18705 13512
rect 16264 13472 16270 13484
rect 4816 13444 4844 13472
rect 4724 13416 4844 13444
rect 1397 13379 1455 13385
rect 1397 13345 1409 13379
rect 1443 13376 1455 13379
rect 1670 13376 1676 13388
rect 1443 13348 1676 13376
rect 1443 13345 1455 13348
rect 1397 13339 1455 13345
rect 1670 13336 1676 13348
rect 1728 13376 1734 13388
rect 1728 13348 3556 13376
rect 1728 13336 1734 13348
rect 1670 13200 1676 13252
rect 1728 13200 1734 13252
rect 2314 13200 2320 13252
rect 2372 13200 2378 13252
rect 3528 13184 3556 13348
rect 4724 13317 4752 13416
rect 4801 13379 4859 13385
rect 4801 13345 4813 13379
rect 4847 13376 4859 13379
rect 4890 13376 4896 13388
rect 4847 13348 4896 13376
rect 4847 13345 4859 13348
rect 4801 13339 4859 13345
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5077 13379 5135 13385
rect 5077 13345 5089 13379
rect 5123 13345 5135 13379
rect 6932 13376 6960 13472
rect 7285 13379 7343 13385
rect 7285 13376 7297 13379
rect 6932 13348 7297 13376
rect 5077 13339 5135 13345
rect 7285 13345 7297 13348
rect 7331 13345 7343 13379
rect 7285 13339 7343 13345
rect 8757 13379 8815 13385
rect 8757 13345 8769 13379
rect 8803 13376 8815 13379
rect 10137 13379 10195 13385
rect 8803 13348 9352 13376
rect 8803 13345 8815 13348
rect 8757 13339 8815 13345
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13277 4767 13311
rect 4709 13271 4767 13277
rect 3510 13132 3516 13184
rect 3568 13132 3574 13184
rect 5092 13172 5120 13339
rect 7006 13268 7012 13320
rect 7064 13268 7070 13320
rect 9122 13268 9128 13320
rect 9180 13268 9186 13320
rect 9324 13317 9352 13348
rect 10137 13345 10149 13379
rect 10183 13376 10195 13379
rect 11974 13376 11980 13388
rect 10183 13348 11980 13376
rect 10183 13345 10195 13348
rect 10137 13339 10195 13345
rect 11974 13336 11980 13348
rect 12032 13336 12038 13388
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13277 9367 13311
rect 9309 13271 9367 13277
rect 10410 13268 10416 13320
rect 10468 13268 10474 13320
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13308 12495 13311
rect 12483 13280 12756 13308
rect 12483 13277 12495 13280
rect 12437 13271 12495 13277
rect 9033 13243 9091 13249
rect 9033 13240 9045 13243
rect 8510 13212 9045 13240
rect 9033 13209 9045 13212
rect 9079 13209 9091 13243
rect 9033 13203 9091 13209
rect 10689 13243 10747 13249
rect 10689 13209 10701 13243
rect 10735 13209 10747 13243
rect 12345 13243 12403 13249
rect 12345 13240 12357 13243
rect 11914 13212 12357 13240
rect 10689 13203 10747 13209
rect 12345 13209 12357 13212
rect 12391 13209 12403 13243
rect 12345 13203 12403 13209
rect 10704 13172 10732 13203
rect 12728 13184 12756 13280
rect 13556 13240 13584 13472
rect 13832 13308 13860 13472
rect 15105 13447 15163 13453
rect 15105 13413 15117 13447
rect 15151 13444 15163 13447
rect 15151 13416 15884 13444
rect 15151 13413 15163 13416
rect 15105 13407 15163 13413
rect 15856 13388 15884 13416
rect 17586 13404 17592 13456
rect 17644 13404 17650 13456
rect 14918 13376 14924 13388
rect 14200 13348 14924 13376
rect 14200 13317 14228 13348
rect 14918 13336 14924 13348
rect 14976 13376 14982 13388
rect 15381 13379 15439 13385
rect 15381 13376 15393 13379
rect 14976 13348 15393 13376
rect 14976 13336 14982 13348
rect 15381 13345 15393 13348
rect 15427 13345 15439 13379
rect 15381 13339 15439 13345
rect 14185 13311 14243 13317
rect 14185 13308 14197 13311
rect 13832 13280 14197 13308
rect 14185 13277 14197 13280
rect 14231 13277 14243 13311
rect 14185 13271 14243 13277
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 15396 13308 15424 13339
rect 15838 13336 15844 13388
rect 15896 13376 15902 13388
rect 16209 13379 16267 13385
rect 16209 13376 16221 13379
rect 15896 13348 16221 13376
rect 15896 13336 15902 13348
rect 16209 13345 16221 13348
rect 16255 13376 16267 13379
rect 16255 13348 17724 13376
rect 16255 13345 16267 13348
rect 16209 13339 16267 13345
rect 16298 13308 16304 13320
rect 15396 13280 16304 13308
rect 14369 13271 14427 13277
rect 14274 13240 14280 13252
rect 13556 13212 14280 13240
rect 14274 13200 14280 13212
rect 14332 13240 14338 13252
rect 14384 13240 14412 13271
rect 16298 13268 16304 13280
rect 16356 13268 16362 13320
rect 16960 13317 16988 13348
rect 17696 13320 17724 13348
rect 16669 13311 16727 13317
rect 16669 13277 16681 13311
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13277 17003 13311
rect 16945 13271 17003 13277
rect 14332 13212 14412 13240
rect 14332 13200 14338 13212
rect 14550 13200 14556 13252
rect 14608 13200 14614 13252
rect 16684 13240 16712 13271
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 17092 13280 17233 13308
rect 17092 13268 17098 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 17678 13268 17684 13320
rect 17736 13308 17742 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17736 13280 17785 13308
rect 17736 13268 17742 13280
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18156 13308 18184 13484
rect 18693 13481 18705 13484
rect 18739 13481 18751 13515
rect 18693 13475 18751 13481
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19242 13512 19248 13524
rect 19015 13484 19248 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 18708 13444 18736 13475
rect 19242 13472 19248 13484
rect 19300 13512 19306 13524
rect 19613 13515 19671 13521
rect 19613 13512 19625 13515
rect 19300 13484 19625 13512
rect 19300 13472 19306 13484
rect 19613 13481 19625 13484
rect 19659 13481 19671 13515
rect 19613 13475 19671 13481
rect 19705 13515 19763 13521
rect 19705 13481 19717 13515
rect 19751 13512 19763 13515
rect 19978 13512 19984 13524
rect 19751 13484 19984 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 21542 13472 21548 13524
rect 21600 13512 21606 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21600 13484 21833 13512
rect 21600 13472 21606 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 21821 13475 21879 13481
rect 22649 13515 22707 13521
rect 22649 13481 22661 13515
rect 22695 13512 22707 13515
rect 23106 13512 23112 13524
rect 22695 13484 23112 13512
rect 22695 13481 22707 13484
rect 22649 13475 22707 13481
rect 23106 13472 23112 13484
rect 23164 13472 23170 13524
rect 26326 13472 26332 13524
rect 26384 13472 26390 13524
rect 28261 13515 28319 13521
rect 28261 13481 28273 13515
rect 28307 13512 28319 13515
rect 29362 13512 29368 13524
rect 28307 13484 29368 13512
rect 28307 13481 28319 13484
rect 28261 13475 28319 13481
rect 29362 13472 29368 13484
rect 29420 13472 29426 13524
rect 30374 13472 30380 13524
rect 30432 13472 30438 13524
rect 30466 13472 30472 13524
rect 30524 13512 30530 13524
rect 30561 13515 30619 13521
rect 30561 13512 30573 13515
rect 30524 13484 30573 13512
rect 30524 13472 30530 13484
rect 30561 13481 30573 13484
rect 30607 13481 30619 13515
rect 30561 13475 30619 13481
rect 34054 13472 34060 13524
rect 34112 13512 34118 13524
rect 34149 13515 34207 13521
rect 34149 13512 34161 13515
rect 34112 13484 34161 13512
rect 34112 13472 34118 13484
rect 34149 13481 34161 13484
rect 34195 13481 34207 13515
rect 34149 13475 34207 13481
rect 19334 13444 19340 13456
rect 18708 13416 19340 13444
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 20809 13447 20867 13453
rect 20809 13413 20821 13447
rect 20855 13413 20867 13447
rect 25038 13444 25044 13456
rect 20809 13407 20867 13413
rect 24688 13416 25044 13444
rect 18506 13336 18512 13388
rect 18564 13376 18570 13388
rect 19521 13379 19579 13385
rect 19521 13376 19533 13379
rect 18564 13348 19533 13376
rect 18564 13336 18570 13348
rect 19521 13345 19533 13348
rect 19567 13376 19579 13379
rect 19567 13348 20576 13376
rect 19567 13345 19579 13348
rect 19521 13339 19579 13345
rect 20548 13320 20576 13348
rect 18003 13280 18184 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18874 13268 18880 13320
rect 18932 13268 18938 13320
rect 19058 13268 19064 13320
rect 19116 13268 19122 13320
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 18322 13240 18328 13252
rect 16684 13212 18328 13240
rect 18322 13200 18328 13212
rect 18380 13240 18386 13252
rect 19260 13240 19288 13271
rect 19426 13268 19432 13320
rect 19484 13308 19490 13320
rect 20070 13308 20076 13320
rect 19484 13280 20076 13308
rect 19484 13268 19490 13280
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 20438 13268 20444 13320
rect 20496 13268 20502 13320
rect 20530 13268 20536 13320
rect 20588 13268 20594 13320
rect 20717 13311 20775 13317
rect 20717 13277 20729 13311
rect 20763 13308 20775 13311
rect 20824 13308 20852 13407
rect 20898 13336 20904 13388
rect 20956 13376 20962 13388
rect 21082 13376 21088 13388
rect 20956 13348 21088 13376
rect 20956 13336 20962 13348
rect 21082 13336 21088 13348
rect 21140 13376 21146 13388
rect 21361 13379 21419 13385
rect 21361 13376 21373 13379
rect 21140 13348 21373 13376
rect 21140 13336 21146 13348
rect 21361 13345 21373 13348
rect 21407 13345 21419 13379
rect 21361 13339 21419 13345
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13376 23351 13379
rect 23339 13348 23888 13376
rect 23339 13345 23351 13348
rect 23293 13339 23351 13345
rect 23860 13320 23888 13348
rect 20763 13280 20852 13308
rect 21177 13311 21235 13317
rect 20763 13277 20775 13280
rect 20717 13271 20775 13277
rect 21177 13277 21189 13311
rect 21223 13308 21235 13311
rect 21266 13308 21272 13320
rect 21223 13280 21272 13308
rect 21223 13277 21235 13280
rect 21177 13271 21235 13277
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 22922 13268 22928 13320
rect 22980 13268 22986 13320
rect 23198 13308 23204 13320
rect 23124 13280 23204 13308
rect 21358 13240 21364 13252
rect 18380 13212 19288 13240
rect 19996 13212 21364 13240
rect 18380 13200 18386 13212
rect 5092 13144 10732 13172
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 13173 13175 13231 13181
rect 13173 13141 13185 13175
rect 13219 13172 13231 13175
rect 13538 13172 13544 13184
rect 13219 13144 13544 13172
rect 13219 13141 13231 13144
rect 13173 13135 13231 13141
rect 13538 13132 13544 13144
rect 13596 13172 13602 13184
rect 14182 13172 14188 13184
rect 13596 13144 14188 13172
rect 13596 13132 13602 13144
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 17402 13132 17408 13184
rect 17460 13132 17466 13184
rect 17494 13132 17500 13184
rect 17552 13172 17558 13184
rect 17865 13175 17923 13181
rect 17865 13172 17877 13175
rect 17552 13144 17877 13172
rect 17552 13132 17558 13144
rect 17865 13141 17877 13144
rect 17911 13141 17923 13175
rect 17865 13135 17923 13141
rect 17954 13132 17960 13184
rect 18012 13172 18018 13184
rect 18141 13175 18199 13181
rect 18141 13172 18153 13175
rect 18012 13144 18153 13172
rect 18012 13132 18018 13144
rect 18141 13141 18153 13144
rect 18187 13172 18199 13175
rect 18506 13172 18512 13184
rect 18187 13144 18512 13172
rect 18187 13141 18199 13144
rect 18141 13135 18199 13141
rect 18506 13132 18512 13144
rect 18564 13132 18570 13184
rect 18782 13132 18788 13184
rect 18840 13172 18846 13184
rect 19150 13172 19156 13184
rect 18840 13144 19156 13172
rect 18840 13132 18846 13144
rect 19150 13132 19156 13144
rect 19208 13172 19214 13184
rect 19996 13181 20024 13212
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 23124 13249 23152 13280
rect 23198 13268 23204 13280
rect 23256 13268 23262 13320
rect 23382 13268 23388 13320
rect 23440 13268 23446 13320
rect 23842 13268 23848 13320
rect 23900 13268 23906 13320
rect 24688 13317 24716 13416
rect 25038 13404 25044 13416
rect 25096 13404 25102 13456
rect 25685 13447 25743 13453
rect 25685 13413 25697 13447
rect 25731 13413 25743 13447
rect 25685 13407 25743 13413
rect 26237 13447 26295 13453
rect 26237 13413 26249 13447
rect 26283 13413 26295 13447
rect 26237 13407 26295 13413
rect 27525 13447 27583 13453
rect 27525 13413 27537 13447
rect 27571 13444 27583 13447
rect 27571 13416 27936 13444
rect 27571 13413 27583 13416
rect 27525 13407 27583 13413
rect 25590 13376 25596 13388
rect 24780 13348 25596 13376
rect 24673 13311 24731 13317
rect 24673 13277 24685 13311
rect 24719 13277 24731 13311
rect 24673 13271 24731 13277
rect 23109 13243 23167 13249
rect 23109 13209 23121 13243
rect 23155 13209 23167 13243
rect 24780 13240 24808 13348
rect 25590 13336 25596 13348
rect 25648 13336 25654 13388
rect 24949 13311 25007 13317
rect 24949 13308 24961 13311
rect 23109 13203 23167 13209
rect 23768 13212 24808 13240
rect 24872 13280 24961 13308
rect 23768 13184 23796 13212
rect 19337 13175 19395 13181
rect 19337 13172 19349 13175
rect 19208 13144 19349 13172
rect 19208 13132 19214 13144
rect 19337 13141 19349 13144
rect 19383 13141 19395 13175
rect 19337 13135 19395 13141
rect 19981 13175 20039 13181
rect 19981 13141 19993 13175
rect 20027 13141 20039 13175
rect 19981 13135 20039 13141
rect 20254 13132 20260 13184
rect 20312 13132 20318 13184
rect 20622 13132 20628 13184
rect 20680 13132 20686 13184
rect 20806 13132 20812 13184
rect 20864 13172 20870 13184
rect 21269 13175 21327 13181
rect 21269 13172 21281 13175
rect 20864 13144 21281 13172
rect 20864 13132 20870 13144
rect 21269 13141 21281 13144
rect 21315 13141 21327 13175
rect 21269 13135 21327 13141
rect 23014 13132 23020 13184
rect 23072 13132 23078 13184
rect 23750 13132 23756 13184
rect 23808 13132 23814 13184
rect 24872 13181 24900 13280
rect 24949 13277 24961 13280
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25222 13268 25228 13320
rect 25280 13268 25286 13320
rect 25501 13311 25559 13317
rect 25501 13277 25513 13311
rect 25547 13277 25559 13311
rect 25501 13271 25559 13277
rect 25516 13240 25544 13271
rect 25148 13212 25544 13240
rect 25608 13240 25636 13336
rect 25700 13308 25728 13407
rect 25884 13348 26188 13376
rect 25777 13311 25835 13317
rect 25777 13308 25789 13311
rect 25700 13280 25789 13308
rect 25777 13277 25789 13280
rect 25823 13277 25835 13311
rect 25777 13271 25835 13277
rect 25884 13240 25912 13348
rect 26053 13311 26111 13317
rect 26053 13308 26065 13311
rect 25608 13212 25912 13240
rect 25976 13280 26065 13308
rect 25148 13181 25176 13212
rect 24857 13175 24915 13181
rect 24857 13141 24869 13175
rect 24903 13141 24915 13175
rect 24857 13135 24915 13141
rect 25133 13175 25191 13181
rect 25133 13141 25145 13175
rect 25179 13141 25191 13175
rect 25133 13135 25191 13141
rect 25406 13132 25412 13184
rect 25464 13132 25470 13184
rect 25976 13181 26004 13280
rect 26053 13277 26065 13280
rect 26099 13277 26111 13311
rect 26053 13271 26111 13277
rect 26160 13240 26188 13348
rect 26252 13308 26280 13407
rect 27249 13379 27307 13385
rect 27249 13345 27261 13379
rect 27295 13376 27307 13379
rect 27430 13376 27436 13388
rect 27295 13348 27436 13376
rect 27295 13345 27307 13348
rect 27249 13339 27307 13345
rect 27430 13336 27436 13348
rect 27488 13336 27494 13388
rect 27908 13385 27936 13416
rect 27893 13379 27951 13385
rect 27893 13345 27905 13379
rect 27939 13345 27951 13379
rect 27893 13339 27951 13345
rect 26513 13311 26571 13317
rect 26513 13308 26525 13311
rect 26252 13280 26525 13308
rect 26513 13277 26525 13280
rect 26559 13277 26571 13311
rect 26513 13271 26571 13277
rect 27157 13311 27215 13317
rect 27157 13277 27169 13311
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 27172 13240 27200 13271
rect 27982 13268 27988 13320
rect 28040 13268 28046 13320
rect 30392 13308 30420 13472
rect 32125 13379 32183 13385
rect 32125 13345 32137 13379
rect 32171 13376 32183 13379
rect 32585 13379 32643 13385
rect 32585 13376 32597 13379
rect 32171 13348 32597 13376
rect 32171 13345 32183 13348
rect 32125 13339 32183 13345
rect 32585 13345 32597 13348
rect 32631 13345 32643 13379
rect 32585 13339 32643 13345
rect 30469 13311 30527 13317
rect 30469 13308 30481 13311
rect 30392 13280 30481 13308
rect 30469 13277 30481 13280
rect 30515 13277 30527 13311
rect 30469 13271 30527 13277
rect 31754 13268 31760 13320
rect 31812 13308 31818 13320
rect 32033 13311 32091 13317
rect 32033 13308 32045 13311
rect 31812 13280 32045 13308
rect 31812 13268 31818 13280
rect 32033 13277 32045 13280
rect 32079 13277 32091 13311
rect 32033 13271 32091 13277
rect 32493 13311 32551 13317
rect 32493 13277 32505 13311
rect 32539 13277 32551 13311
rect 32493 13271 32551 13277
rect 26160 13212 27200 13240
rect 31294 13200 31300 13252
rect 31352 13240 31358 13252
rect 32508 13240 32536 13271
rect 32674 13268 32680 13320
rect 32732 13308 32738 13320
rect 32953 13311 33011 13317
rect 32953 13308 32965 13311
rect 32732 13280 32965 13308
rect 32732 13268 32738 13280
rect 32953 13277 32965 13280
rect 32999 13277 33011 13311
rect 32953 13271 33011 13277
rect 34057 13311 34115 13317
rect 34057 13277 34069 13311
rect 34103 13308 34115 13311
rect 34517 13311 34575 13317
rect 34103 13280 34137 13308
rect 34103 13277 34115 13280
rect 34057 13271 34115 13277
rect 34517 13277 34529 13311
rect 34563 13308 34575 13311
rect 34563 13280 34597 13308
rect 34563 13277 34575 13280
rect 34517 13271 34575 13277
rect 31352 13212 32536 13240
rect 33597 13243 33655 13249
rect 31352 13200 31358 13212
rect 33597 13209 33609 13243
rect 33643 13240 33655 13243
rect 33870 13240 33876 13252
rect 33643 13212 33876 13240
rect 33643 13209 33655 13212
rect 33597 13203 33655 13209
rect 33870 13200 33876 13212
rect 33928 13240 33934 13252
rect 34072 13240 34100 13271
rect 34532 13240 34560 13271
rect 33928 13212 34560 13240
rect 33928 13200 33934 13212
rect 34532 13184 34560 13212
rect 25961 13175 26019 13181
rect 25961 13141 25973 13175
rect 26007 13141 26019 13175
rect 25961 13135 26019 13141
rect 26418 13132 26424 13184
rect 26476 13172 26482 13184
rect 27246 13172 27252 13184
rect 26476 13144 27252 13172
rect 26476 13132 26482 13144
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 32398 13132 32404 13184
rect 32456 13132 32462 13184
rect 34422 13132 34428 13184
rect 34480 13132 34486 13184
rect 34514 13132 34520 13184
rect 34572 13132 34578 13184
rect 1104 13082 35236 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 35236 13082
rect 1104 13008 35236 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12937 1639 12971
rect 1581 12931 1639 12937
rect 1596 12900 1624 12931
rect 2314 12928 2320 12980
rect 2372 12928 2378 12980
rect 4525 12971 4583 12977
rect 2700 12940 3096 12968
rect 2700 12900 2728 12940
rect 3068 12909 3096 12940
rect 4525 12937 4537 12971
rect 4571 12968 4583 12971
rect 5258 12968 5264 12980
rect 4571 12940 5264 12968
rect 4571 12937 4583 12940
rect 4525 12931 4583 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 5534 12928 5540 12980
rect 5592 12968 5598 12980
rect 5645 12971 5703 12977
rect 5645 12968 5657 12971
rect 5592 12940 5657 12968
rect 5592 12928 5598 12940
rect 5645 12937 5657 12940
rect 5691 12937 5703 12971
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 5645 12931 5703 12937
rect 9646 12940 10333 12968
rect 1596 12872 2728 12900
rect 3053 12903 3111 12909
rect 3053 12869 3065 12903
rect 3099 12869 3111 12903
rect 4709 12903 4767 12909
rect 4709 12900 4721 12903
rect 4278 12872 4721 12900
rect 3053 12863 3111 12869
rect 4709 12869 4721 12872
rect 4755 12869 4767 12903
rect 4709 12863 4767 12869
rect 4982 12860 4988 12912
rect 5040 12900 5046 12912
rect 5077 12903 5135 12909
rect 5077 12900 5089 12903
rect 5040 12872 5089 12900
rect 5040 12860 5046 12872
rect 5077 12869 5089 12872
rect 5123 12869 5135 12903
rect 5077 12863 5135 12869
rect 5442 12860 5448 12912
rect 5500 12860 5506 12912
rect 934 12792 940 12844
rect 992 12832 998 12844
rect 1397 12835 1455 12841
rect 1397 12832 1409 12835
rect 992 12804 1409 12832
rect 992 12792 998 12804
rect 1397 12801 1409 12804
rect 1443 12801 1455 12835
rect 2225 12835 2283 12841
rect 2225 12832 2237 12835
rect 1397 12795 1455 12801
rect 2148 12804 2237 12832
rect 2148 12640 2176 12804
rect 2225 12801 2237 12804
rect 2271 12801 2283 12835
rect 2225 12795 2283 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 5000 12832 5028 12860
rect 4847 12804 5028 12832
rect 8021 12835 8079 12841
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 8021 12801 8033 12835
rect 8067 12832 8079 12835
rect 8067 12804 8616 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 2777 12767 2835 12773
rect 2777 12733 2789 12767
rect 2823 12733 2835 12767
rect 2777 12727 2835 12733
rect 2130 12588 2136 12640
rect 2188 12588 2194 12640
rect 2792 12628 2820 12727
rect 3510 12628 3516 12640
rect 2792 12600 3516 12628
rect 3510 12588 3516 12600
rect 3568 12588 3574 12640
rect 5626 12588 5632 12640
rect 5684 12588 5690 12640
rect 5810 12588 5816 12640
rect 5868 12588 5874 12640
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8294 12628 8300 12640
rect 8159 12600 8300 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8588 12637 8616 12804
rect 8754 12656 8760 12708
rect 8812 12696 8818 12708
rect 8849 12699 8907 12705
rect 8849 12696 8861 12699
rect 8812 12668 8861 12696
rect 8812 12656 8818 12668
rect 8849 12665 8861 12668
rect 8895 12696 8907 12699
rect 9646 12696 9674 12940
rect 10321 12937 10333 12940
rect 10367 12968 10379 12971
rect 10410 12968 10416 12980
rect 10367 12940 10416 12968
rect 10367 12937 10379 12940
rect 10321 12931 10379 12937
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 12437 12971 12495 12977
rect 12437 12937 12449 12971
rect 12483 12968 12495 12971
rect 12986 12968 12992 12980
rect 12483 12940 12992 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 12636 12844 12664 12940
rect 12986 12928 12992 12940
rect 13044 12928 13050 12980
rect 13814 12928 13820 12980
rect 13872 12928 13878 12980
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12968 14151 12971
rect 14182 12968 14188 12980
rect 14139 12940 14188 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 14182 12928 14188 12940
rect 14240 12928 14246 12980
rect 14550 12928 14556 12980
rect 14608 12928 14614 12980
rect 16298 12928 16304 12980
rect 16356 12968 16362 12980
rect 17405 12971 17463 12977
rect 17405 12968 17417 12971
rect 16356 12940 17417 12968
rect 16356 12928 16362 12940
rect 17405 12937 17417 12940
rect 17451 12968 17463 12971
rect 17494 12968 17500 12980
rect 17451 12940 17500 12968
rect 17451 12937 17463 12940
rect 17405 12931 17463 12937
rect 17494 12928 17500 12940
rect 17552 12928 17558 12980
rect 18693 12971 18751 12977
rect 18693 12968 18705 12971
rect 17788 12940 18705 12968
rect 14568 12900 14596 12928
rect 14568 12872 14780 12900
rect 12618 12792 12624 12844
rect 12676 12792 12682 12844
rect 12802 12792 12808 12844
rect 12860 12792 12866 12844
rect 13906 12832 13912 12844
rect 13464 12804 13912 12832
rect 8895 12668 9674 12696
rect 8895 12665 8907 12668
rect 8849 12659 8907 12665
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 13464 12705 13492 12804
rect 13906 12792 13912 12804
rect 13964 12832 13970 12844
rect 14001 12835 14059 12841
rect 14001 12832 14013 12835
rect 13964 12804 14013 12832
rect 13964 12792 13970 12804
rect 14001 12801 14013 12804
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 13449 12699 13507 12705
rect 13449 12696 13461 12699
rect 11020 12668 13461 12696
rect 11020 12656 11026 12668
rect 13449 12665 13461 12668
rect 13495 12665 13507 12699
rect 14016 12696 14044 12795
rect 14274 12792 14280 12844
rect 14332 12792 14338 12844
rect 14752 12841 14780 12872
rect 15654 12860 15660 12912
rect 15712 12900 15718 12912
rect 16666 12900 16672 12912
rect 15712 12872 16672 12900
rect 15712 12860 15718 12872
rect 16666 12860 16672 12872
rect 16724 12900 16730 12912
rect 16724 12872 17080 12900
rect 16724 12860 16730 12872
rect 14461 12835 14519 12841
rect 14461 12801 14473 12835
rect 14507 12832 14519 12835
rect 14553 12835 14611 12841
rect 14553 12832 14565 12835
rect 14507 12804 14565 12832
rect 14507 12801 14519 12804
rect 14461 12795 14519 12801
rect 14553 12801 14565 12804
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12801 14795 12835
rect 14737 12795 14795 12801
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15105 12835 15163 12841
rect 15105 12801 15117 12835
rect 15151 12832 15163 12835
rect 15930 12832 15936 12844
rect 15151 12804 15936 12832
rect 15151 12801 15163 12804
rect 15105 12795 15163 12801
rect 14826 12724 14832 12776
rect 14884 12724 14890 12776
rect 15120 12696 15148 12795
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 16117 12835 16175 12841
rect 16117 12801 16129 12835
rect 16163 12801 16175 12835
rect 16117 12795 16175 12801
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 16132 12764 16160 12795
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 16776 12841 16804 12872
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 16264 12804 16313 12832
rect 16264 12792 16270 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 16945 12835 17003 12841
rect 16945 12832 16957 12835
rect 16908 12804 16957 12832
rect 16908 12792 16914 12804
rect 16945 12801 16957 12804
rect 16991 12801 17003 12835
rect 17052 12832 17080 12872
rect 17788 12832 17816 12940
rect 18693 12937 18705 12940
rect 18739 12968 18751 12971
rect 19058 12968 19064 12980
rect 18739 12940 19064 12968
rect 18739 12937 18751 12940
rect 18693 12931 18751 12937
rect 19058 12928 19064 12940
rect 19116 12928 19122 12980
rect 19150 12928 19156 12980
rect 19208 12968 19214 12980
rect 19208 12940 19472 12968
rect 19208 12928 19214 12940
rect 18966 12900 18972 12912
rect 17052 12804 17816 12832
rect 17866 12872 18972 12900
rect 16945 12795 17003 12801
rect 15620 12736 16988 12764
rect 15620 12724 15626 12736
rect 15654 12696 15660 12708
rect 14016 12668 15148 12696
rect 15212 12668 15660 12696
rect 13449 12659 13507 12665
rect 8573 12631 8631 12637
rect 8573 12597 8585 12631
rect 8619 12628 8631 12631
rect 8662 12628 8668 12640
rect 8619 12600 8668 12628
rect 8619 12597 8631 12600
rect 8573 12591 8631 12597
rect 8662 12588 8668 12600
rect 8720 12628 8726 12640
rect 9122 12628 9128 12640
rect 8720 12600 9128 12628
rect 8720 12588 8726 12600
rect 9122 12588 9128 12600
rect 9180 12628 9186 12640
rect 9217 12631 9275 12637
rect 9217 12628 9229 12631
rect 9180 12600 9229 12628
rect 9180 12588 9186 12600
rect 9217 12597 9229 12600
rect 9263 12597 9275 12631
rect 9217 12591 9275 12597
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12621 12631 12679 12637
rect 12621 12628 12633 12631
rect 12492 12600 12633 12628
rect 12492 12588 12498 12600
rect 12621 12597 12633 12600
rect 12667 12597 12679 12631
rect 12621 12591 12679 12597
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 15102 12628 15108 12640
rect 14332 12600 15108 12628
rect 14332 12588 14338 12600
rect 15102 12588 15108 12600
rect 15160 12628 15166 12640
rect 15212 12628 15240 12668
rect 15654 12656 15660 12668
rect 15712 12656 15718 12708
rect 15930 12656 15936 12708
rect 15988 12696 15994 12708
rect 16850 12696 16856 12708
rect 15988 12668 16856 12696
rect 15988 12656 15994 12668
rect 16850 12656 16856 12668
rect 16908 12656 16914 12708
rect 16960 12696 16988 12736
rect 17494 12724 17500 12776
rect 17552 12764 17558 12776
rect 17866 12764 17894 12872
rect 18966 12860 18972 12872
rect 19024 12900 19030 12912
rect 19334 12900 19340 12912
rect 19024 12872 19340 12900
rect 19024 12860 19030 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 19444 12900 19472 12940
rect 19518 12928 19524 12980
rect 19576 12977 19582 12980
rect 19576 12971 19595 12977
rect 19583 12937 19595 12971
rect 19576 12931 19595 12937
rect 19705 12971 19763 12977
rect 19705 12937 19717 12971
rect 19751 12968 19763 12971
rect 20438 12968 20444 12980
rect 19751 12940 20444 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 19576 12928 19582 12931
rect 20438 12928 20444 12940
rect 20496 12928 20502 12980
rect 23658 12928 23664 12980
rect 23716 12968 23722 12980
rect 23845 12971 23903 12977
rect 23845 12968 23857 12971
rect 23716 12940 23857 12968
rect 23716 12928 23722 12940
rect 23845 12937 23857 12940
rect 23891 12937 23903 12971
rect 23845 12931 23903 12937
rect 24489 12971 24547 12977
rect 24489 12937 24501 12971
rect 24535 12968 24547 12971
rect 24578 12968 24584 12980
rect 24535 12940 24584 12968
rect 24535 12937 24547 12940
rect 24489 12931 24547 12937
rect 24578 12928 24584 12940
rect 24636 12928 24642 12980
rect 24670 12928 24676 12980
rect 24728 12968 24734 12980
rect 24765 12971 24823 12977
rect 24765 12968 24777 12971
rect 24728 12940 24777 12968
rect 24728 12928 24734 12940
rect 24765 12937 24777 12940
rect 24811 12937 24823 12971
rect 24765 12931 24823 12937
rect 25038 12928 25044 12980
rect 25096 12928 25102 12980
rect 25133 12971 25191 12977
rect 25133 12937 25145 12971
rect 25179 12968 25191 12971
rect 25222 12968 25228 12980
rect 25179 12940 25228 12968
rect 25179 12937 25191 12940
rect 25133 12931 25191 12937
rect 25222 12928 25228 12940
rect 25280 12928 25286 12980
rect 25314 12928 25320 12980
rect 25372 12968 25378 12980
rect 25685 12971 25743 12977
rect 25685 12968 25697 12971
rect 25372 12940 25697 12968
rect 25372 12928 25378 12940
rect 25685 12937 25697 12940
rect 25731 12937 25743 12971
rect 25685 12931 25743 12937
rect 25961 12971 26019 12977
rect 25961 12937 25973 12971
rect 26007 12937 26019 12971
rect 27614 12968 27620 12980
rect 25961 12931 26019 12937
rect 26712 12940 27620 12968
rect 19981 12903 20039 12909
rect 19981 12900 19993 12903
rect 19444 12872 19993 12900
rect 19981 12869 19993 12872
rect 20027 12900 20039 12903
rect 20533 12903 20591 12909
rect 20533 12900 20545 12903
rect 20027 12872 20545 12900
rect 20027 12869 20039 12872
rect 19981 12863 20039 12869
rect 20533 12869 20545 12872
rect 20579 12900 20591 12903
rect 20898 12900 20904 12912
rect 20579 12872 20904 12900
rect 20579 12869 20591 12872
rect 20533 12863 20591 12869
rect 20898 12860 20904 12872
rect 20956 12860 20962 12912
rect 24596 12900 24624 12928
rect 25056 12900 25084 12928
rect 25976 12900 26004 12931
rect 24596 12872 24716 12900
rect 25056 12872 26004 12900
rect 18414 12792 18420 12844
rect 18472 12832 18478 12844
rect 20162 12832 20168 12844
rect 18472 12804 20168 12832
rect 18472 12792 18478 12804
rect 20162 12792 20168 12804
rect 20220 12832 20226 12844
rect 23382 12832 23388 12844
rect 20220 12804 23388 12832
rect 20220 12792 20226 12804
rect 23382 12792 23388 12804
rect 23440 12832 23446 12844
rect 24394 12832 24400 12844
rect 23440 12804 24400 12832
rect 23440 12792 23446 12804
rect 24394 12792 24400 12804
rect 24452 12792 24458 12844
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24544 12804 24593 12832
rect 24544 12792 24550 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24688 12832 24716 12872
rect 24857 12835 24915 12841
rect 24857 12832 24869 12835
rect 24688 12804 24869 12832
rect 24581 12795 24639 12801
rect 24857 12801 24869 12804
rect 24903 12801 24915 12835
rect 24857 12795 24915 12801
rect 24946 12792 24952 12844
rect 25004 12792 25010 12844
rect 25593 12835 25651 12841
rect 25593 12801 25605 12835
rect 25639 12801 25651 12835
rect 25593 12795 25651 12801
rect 17552 12736 17894 12764
rect 17552 12724 17558 12736
rect 19334 12724 19340 12776
rect 19392 12764 19398 12776
rect 19518 12764 19524 12776
rect 19392 12736 19524 12764
rect 19392 12724 19398 12736
rect 19518 12724 19524 12736
rect 19576 12764 19582 12776
rect 20806 12764 20812 12776
rect 19576 12736 20812 12764
rect 19576 12724 19582 12736
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 23293 12767 23351 12773
rect 23293 12733 23305 12767
rect 23339 12764 23351 12767
rect 23842 12764 23848 12776
rect 23339 12736 23848 12764
rect 23339 12733 23351 12736
rect 23293 12727 23351 12733
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 24118 12724 24124 12776
rect 24176 12724 24182 12776
rect 24302 12724 24308 12776
rect 24360 12764 24366 12776
rect 24964 12764 24992 12792
rect 24360 12736 24992 12764
rect 24360 12724 24366 12736
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 25498 12764 25504 12776
rect 25096 12736 25504 12764
rect 25096 12724 25102 12736
rect 25498 12724 25504 12736
rect 25556 12724 25562 12776
rect 25608 12764 25636 12795
rect 25774 12792 25780 12844
rect 25832 12792 25838 12844
rect 25866 12792 25872 12844
rect 25924 12792 25930 12844
rect 26142 12792 26148 12844
rect 26200 12792 26206 12844
rect 26418 12792 26424 12844
rect 26476 12792 26482 12844
rect 26605 12835 26663 12841
rect 26605 12801 26617 12835
rect 26651 12801 26663 12835
rect 26712 12832 26740 12940
rect 27614 12928 27620 12940
rect 27672 12928 27678 12980
rect 27801 12971 27859 12977
rect 27801 12937 27813 12971
rect 27847 12968 27859 12971
rect 27982 12968 27988 12980
rect 27847 12940 27988 12968
rect 27847 12937 27859 12940
rect 27801 12931 27859 12937
rect 27982 12928 27988 12940
rect 28040 12928 28046 12980
rect 28537 12971 28595 12977
rect 28537 12937 28549 12971
rect 28583 12968 28595 12971
rect 29270 12968 29276 12980
rect 28583 12940 29276 12968
rect 28583 12937 28595 12940
rect 28537 12931 28595 12937
rect 26789 12903 26847 12909
rect 26789 12869 26801 12903
rect 26835 12900 26847 12903
rect 27065 12903 27123 12909
rect 27065 12900 27077 12903
rect 26835 12872 27077 12900
rect 26835 12869 26847 12872
rect 26789 12863 26847 12869
rect 27065 12869 27077 12872
rect 27111 12900 27123 12903
rect 27111 12872 27568 12900
rect 27111 12869 27123 12872
rect 27065 12863 27123 12869
rect 26973 12835 27031 12841
rect 26973 12832 26985 12835
rect 26712 12804 26985 12832
rect 26605 12795 26663 12801
rect 26973 12801 26985 12804
rect 27019 12801 27031 12835
rect 26973 12795 27031 12801
rect 25792 12764 25820 12792
rect 26050 12764 26056 12776
rect 25608 12736 25728 12764
rect 25792 12736 26056 12764
rect 17586 12696 17592 12708
rect 16960 12668 17592 12696
rect 17586 12656 17592 12668
rect 17644 12696 17650 12708
rect 17865 12699 17923 12705
rect 17865 12696 17877 12699
rect 17644 12668 17877 12696
rect 17644 12656 17650 12668
rect 17865 12665 17877 12668
rect 17911 12665 17923 12699
rect 17865 12659 17923 12665
rect 19058 12656 19064 12708
rect 19116 12696 19122 12708
rect 21177 12699 21235 12705
rect 21177 12696 21189 12699
rect 19116 12668 21189 12696
rect 19116 12656 19122 12668
rect 21177 12665 21189 12668
rect 21223 12696 21235 12699
rect 21542 12696 21548 12708
rect 21223 12668 21548 12696
rect 21223 12665 21235 12668
rect 21177 12659 21235 12665
rect 21542 12656 21548 12668
rect 21600 12656 21606 12708
rect 23750 12656 23756 12708
rect 23808 12656 23814 12708
rect 24136 12696 24164 12724
rect 24136 12668 24716 12696
rect 15160 12600 15240 12628
rect 15160 12588 15166 12600
rect 15286 12588 15292 12640
rect 15344 12588 15350 12640
rect 16206 12588 16212 12640
rect 16264 12588 16270 12640
rect 16945 12631 17003 12637
rect 16945 12597 16957 12631
rect 16991 12628 17003 12631
rect 17218 12628 17224 12640
rect 16991 12600 17224 12628
rect 16991 12597 17003 12600
rect 16945 12591 17003 12597
rect 17218 12588 17224 12600
rect 17276 12588 17282 12640
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18325 12631 18383 12637
rect 18325 12628 18337 12631
rect 18012 12600 18337 12628
rect 18012 12588 18018 12600
rect 18325 12597 18337 12600
rect 18371 12628 18383 12631
rect 18874 12628 18880 12640
rect 18371 12600 18880 12628
rect 18371 12597 18383 12600
rect 18325 12591 18383 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 19334 12588 19340 12640
rect 19392 12628 19398 12640
rect 19521 12631 19579 12637
rect 19521 12628 19533 12631
rect 19392 12600 19533 12628
rect 19392 12588 19398 12600
rect 19521 12597 19533 12600
rect 19567 12628 19579 12631
rect 20070 12628 20076 12640
rect 19567 12600 20076 12628
rect 19567 12597 19579 12600
rect 19521 12591 19579 12597
rect 20070 12588 20076 12600
rect 20128 12628 20134 12640
rect 20438 12628 20444 12640
rect 20128 12600 20444 12628
rect 20128 12588 20134 12600
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 24210 12588 24216 12640
rect 24268 12588 24274 12640
rect 24302 12588 24308 12640
rect 24360 12588 24366 12640
rect 24688 12628 24716 12668
rect 24854 12656 24860 12708
rect 24912 12696 24918 12708
rect 25314 12696 25320 12708
rect 24912 12668 25320 12696
rect 24912 12656 24918 12668
rect 25314 12656 25320 12668
rect 25372 12656 25378 12708
rect 25409 12699 25467 12705
rect 25409 12665 25421 12699
rect 25455 12696 25467 12699
rect 25590 12696 25596 12708
rect 25455 12668 25596 12696
rect 25455 12665 25467 12668
rect 25409 12659 25467 12665
rect 25590 12656 25596 12668
rect 25648 12656 25654 12708
rect 25700 12696 25728 12736
rect 26050 12724 26056 12736
rect 26108 12764 26114 12776
rect 26620 12764 26648 12795
rect 27154 12792 27160 12844
rect 27212 12832 27218 12844
rect 27540 12841 27568 12872
rect 27632 12841 27660 12928
rect 28644 12844 28672 12940
rect 29270 12928 29276 12940
rect 29328 12928 29334 12980
rect 32398 12928 32404 12980
rect 32456 12928 32462 12980
rect 32953 12971 33011 12977
rect 32953 12937 32965 12971
rect 32999 12968 33011 12971
rect 33042 12968 33048 12980
rect 32999 12940 33048 12968
rect 32999 12937 33011 12940
rect 32953 12931 33011 12937
rect 33042 12928 33048 12940
rect 33100 12928 33106 12980
rect 29638 12860 29644 12912
rect 29696 12860 29702 12912
rect 32416 12900 32444 12928
rect 33321 12903 33379 12909
rect 33321 12900 33333 12903
rect 32416 12872 33333 12900
rect 33321 12869 33333 12872
rect 33367 12869 33379 12903
rect 33321 12863 33379 12869
rect 27249 12835 27307 12841
rect 27249 12832 27261 12835
rect 27212 12804 27261 12832
rect 27212 12792 27218 12804
rect 27249 12801 27261 12804
rect 27295 12801 27307 12835
rect 27249 12795 27307 12801
rect 27525 12835 27583 12841
rect 27525 12801 27537 12835
rect 27571 12801 27583 12835
rect 27525 12795 27583 12801
rect 27617 12835 27675 12841
rect 27617 12801 27629 12835
rect 27663 12801 27675 12835
rect 27617 12795 27675 12801
rect 26108 12736 26648 12764
rect 26108 12724 26114 12736
rect 25774 12696 25780 12708
rect 25700 12668 25780 12696
rect 25774 12656 25780 12668
rect 25832 12656 25838 12708
rect 25133 12631 25191 12637
rect 25133 12628 25145 12631
rect 24688 12600 25145 12628
rect 25133 12597 25145 12600
rect 25179 12628 25191 12631
rect 27264 12628 27292 12795
rect 27706 12792 27712 12844
rect 27764 12832 27770 12844
rect 27764 12804 27936 12832
rect 27764 12792 27770 12804
rect 27433 12767 27491 12773
rect 27433 12733 27445 12767
rect 27479 12764 27491 12767
rect 27801 12767 27859 12773
rect 27801 12764 27813 12767
rect 27479 12736 27813 12764
rect 27479 12733 27491 12736
rect 27433 12727 27491 12733
rect 27801 12733 27813 12736
rect 27847 12733 27859 12767
rect 27908 12764 27936 12804
rect 28626 12792 28632 12844
rect 28684 12792 28690 12844
rect 33042 12792 33048 12844
rect 33100 12792 33106 12844
rect 34422 12792 34428 12844
rect 34480 12792 34486 12844
rect 28905 12767 28963 12773
rect 28905 12764 28917 12767
rect 27908 12736 28917 12764
rect 27801 12727 27859 12733
rect 28905 12733 28917 12736
rect 28951 12733 28963 12767
rect 28905 12727 28963 12733
rect 25179 12600 27292 12628
rect 30377 12631 30435 12637
rect 25179 12597 25191 12600
rect 25133 12591 25191 12597
rect 30377 12597 30389 12631
rect 30423 12628 30435 12631
rect 30834 12628 30840 12640
rect 30423 12600 30840 12628
rect 30423 12597 30435 12600
rect 30377 12591 30435 12597
rect 30834 12588 30840 12600
rect 30892 12588 30898 12640
rect 34422 12588 34428 12640
rect 34480 12628 34486 12640
rect 34793 12631 34851 12637
rect 34793 12628 34805 12631
rect 34480 12600 34805 12628
rect 34480 12588 34486 12600
rect 34793 12597 34805 12600
rect 34839 12597 34851 12631
rect 34793 12591 34851 12597
rect 1104 12538 35248 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 35248 12538
rect 1104 12464 35248 12486
rect 3510 12384 3516 12436
rect 3568 12424 3574 12436
rect 4617 12427 4675 12433
rect 4617 12424 4629 12427
rect 3568 12396 4629 12424
rect 3568 12384 3574 12396
rect 4617 12393 4629 12396
rect 4663 12424 4675 12427
rect 5350 12424 5356 12436
rect 4663 12396 5356 12424
rect 4663 12393 4675 12396
rect 4617 12387 4675 12393
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 17865 12427 17923 12433
rect 17865 12424 17877 12427
rect 17328 12396 17877 12424
rect 12802 12316 12808 12368
rect 12860 12356 12866 12368
rect 16117 12359 16175 12365
rect 16117 12356 16129 12359
rect 12860 12328 16129 12356
rect 12860 12316 12866 12328
rect 16117 12325 16129 12328
rect 16163 12325 16175 12359
rect 16117 12319 16175 12325
rect 5810 12248 5816 12300
rect 5868 12248 5874 12300
rect 6273 12291 6331 12297
rect 6273 12257 6285 12291
rect 6319 12288 6331 12291
rect 7285 12291 7343 12297
rect 7285 12288 7297 12291
rect 6319 12260 7297 12288
rect 6319 12257 6331 12260
rect 6273 12251 6331 12257
rect 7285 12257 7297 12260
rect 7331 12257 7343 12291
rect 7285 12251 7343 12257
rect 8757 12291 8815 12297
rect 8757 12257 8769 12291
rect 8803 12288 8815 12291
rect 10965 12291 11023 12297
rect 8803 12260 10456 12288
rect 8803 12257 8815 12260
rect 8757 12251 8815 12257
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 5166 12220 5172 12232
rect 4672 12192 5172 12220
rect 4672 12180 4678 12192
rect 5166 12180 5172 12192
rect 5224 12220 5230 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5224 12192 5917 12220
rect 5224 12180 5230 12192
rect 5905 12189 5917 12192
rect 5951 12189 5963 12223
rect 5905 12183 5963 12189
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 7006 12220 7012 12232
rect 6733 12183 6791 12189
rect 6840 12192 7012 12220
rect 5350 12112 5356 12164
rect 5408 12112 5414 12164
rect 5534 12112 5540 12164
rect 5592 12152 5598 12164
rect 6748 12152 6776 12183
rect 5592 12124 6776 12152
rect 6840 12152 6868 12192
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 10428 12229 10456 12260
rect 10965 12257 10977 12291
rect 11011 12288 11023 12291
rect 11514 12288 11520 12300
rect 11011 12260 11520 12288
rect 11011 12257 11023 12260
rect 10965 12251 11023 12257
rect 11514 12248 11520 12260
rect 11572 12248 11578 12300
rect 15654 12248 15660 12300
rect 15712 12288 15718 12300
rect 16132 12288 16160 12319
rect 17328 12288 17356 12396
rect 17865 12393 17877 12396
rect 17911 12424 17923 12427
rect 17954 12424 17960 12436
rect 17911 12396 17960 12424
rect 17911 12393 17923 12396
rect 17865 12387 17923 12393
rect 17954 12384 17960 12396
rect 18012 12424 18018 12436
rect 18012 12396 19334 12424
rect 18012 12384 18018 12396
rect 17494 12316 17500 12368
rect 17552 12316 17558 12368
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 19306 12356 19334 12396
rect 19518 12384 19524 12436
rect 19576 12384 19582 12436
rect 19978 12384 19984 12436
rect 20036 12384 20042 12436
rect 20717 12427 20775 12433
rect 20717 12393 20729 12427
rect 20763 12424 20775 12427
rect 25225 12427 25283 12433
rect 20763 12396 22048 12424
rect 20763 12393 20775 12396
rect 20717 12387 20775 12393
rect 20993 12359 21051 12365
rect 20993 12356 21005 12359
rect 17828 12328 18920 12356
rect 19306 12328 21005 12356
rect 17828 12316 17834 12328
rect 15712 12260 15792 12288
rect 16132 12260 16988 12288
rect 15712 12248 15718 12260
rect 10413 12223 10471 12229
rect 10413 12189 10425 12223
rect 10459 12189 10471 12223
rect 10413 12183 10471 12189
rect 12434 12180 12440 12232
rect 12492 12180 12498 12232
rect 12802 12180 12808 12232
rect 12860 12180 12866 12232
rect 14550 12180 14556 12232
rect 14608 12180 14614 12232
rect 14826 12180 14832 12232
rect 14884 12180 14890 12232
rect 15764 12220 15792 12260
rect 16960 12229 16988 12260
rect 17052 12260 17356 12288
rect 16301 12223 16359 12229
rect 16301 12220 16313 12223
rect 15764 12192 16313 12220
rect 16301 12189 16313 12192
rect 16347 12189 16359 12223
rect 16761 12223 16819 12229
rect 16761 12220 16773 12223
rect 16301 12183 16359 12189
rect 16500 12192 16773 12220
rect 15660 12164 15712 12170
rect 6840 12124 7696 12152
rect 5592 12112 5598 12124
rect 5368 12084 5396 12112
rect 6840 12084 6868 12124
rect 5368 12056 6868 12084
rect 6917 12087 6975 12093
rect 6917 12053 6929 12087
rect 6963 12084 6975 12087
rect 7558 12084 7564 12096
rect 6963 12056 7564 12084
rect 6963 12053 6975 12056
rect 6917 12047 6975 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 7668 12084 7696 12124
rect 8294 12112 8300 12164
rect 8352 12112 8358 12164
rect 13570 12124 15056 12152
rect 8202 12084 8208 12096
rect 7668 12056 8208 12084
rect 8202 12044 8208 12056
rect 8260 12084 8266 12096
rect 8754 12084 8760 12096
rect 8260 12056 8760 12084
rect 8260 12044 8266 12056
rect 8754 12044 8760 12056
rect 8812 12084 8818 12096
rect 9030 12084 9036 12096
rect 8812 12056 9036 12084
rect 8812 12044 8818 12056
rect 9030 12044 9036 12056
rect 9088 12084 9094 12096
rect 9125 12087 9183 12093
rect 9125 12084 9137 12087
rect 9088 12056 9137 12084
rect 9088 12044 9094 12056
rect 9125 12053 9137 12056
rect 9171 12053 9183 12087
rect 15028 12084 15056 12124
rect 16500 12161 16528 12192
rect 16761 12189 16773 12192
rect 16807 12189 16819 12223
rect 16761 12183 16819 12189
rect 16945 12223 17003 12229
rect 16945 12189 16957 12223
rect 16991 12189 17003 12223
rect 16945 12183 17003 12189
rect 16485 12155 16543 12161
rect 16485 12152 16497 12155
rect 15660 12106 15712 12112
rect 15856 12124 16497 12152
rect 15856 12096 15884 12124
rect 16485 12121 16497 12124
rect 16531 12121 16543 12155
rect 16776 12152 16804 12183
rect 17052 12152 17080 12260
rect 17402 12248 17408 12300
rect 17460 12288 17466 12300
rect 18046 12288 18052 12300
rect 17460 12260 18052 12288
rect 17460 12248 17466 12260
rect 18046 12248 18052 12260
rect 18104 12288 18110 12300
rect 18104 12260 18828 12288
rect 18104 12248 18110 12260
rect 17218 12180 17224 12232
rect 17276 12180 17282 12232
rect 17313 12223 17371 12229
rect 17313 12189 17325 12223
rect 17359 12220 17371 12223
rect 17420 12220 17448 12248
rect 18141 12223 18199 12229
rect 18141 12220 18153 12223
rect 17359 12192 17448 12220
rect 18064 12192 18153 12220
rect 17359 12189 17371 12192
rect 17313 12183 17371 12189
rect 16776 12124 17080 12152
rect 17129 12155 17187 12161
rect 16485 12115 16543 12121
rect 17129 12121 17141 12155
rect 17175 12152 17187 12155
rect 17497 12155 17555 12161
rect 17497 12152 17509 12155
rect 17175 12124 17509 12152
rect 17175 12121 17187 12124
rect 17129 12115 17187 12121
rect 17497 12121 17509 12124
rect 17543 12152 17555 12155
rect 17678 12152 17684 12164
rect 17543 12124 17684 12152
rect 17543 12121 17555 12124
rect 17497 12115 17555 12121
rect 17678 12112 17684 12124
rect 17736 12112 17742 12164
rect 15194 12084 15200 12096
rect 15028 12056 15200 12084
rect 9125 12047 9183 12053
rect 15194 12044 15200 12056
rect 15252 12044 15258 12096
rect 15838 12044 15844 12096
rect 15896 12044 15902 12096
rect 15930 12044 15936 12096
rect 15988 12084 15994 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 15988 12056 16405 12084
rect 15988 12044 15994 12056
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 16669 12087 16727 12093
rect 16669 12053 16681 12087
rect 16715 12084 16727 12087
rect 16942 12084 16948 12096
rect 16715 12056 16948 12084
rect 16715 12053 16727 12056
rect 16669 12047 16727 12053
rect 16942 12044 16948 12056
rect 17000 12084 17006 12096
rect 17770 12084 17776 12096
rect 17000 12056 17776 12084
rect 17000 12044 17006 12056
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 17954 12044 17960 12096
rect 18012 12044 18018 12096
rect 18064 12084 18092 12192
rect 18141 12189 18153 12192
rect 18187 12189 18199 12223
rect 18141 12183 18199 12189
rect 18230 12180 18236 12232
rect 18288 12180 18294 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18340 12192 18705 12220
rect 18340 12084 18368 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18417 12087 18475 12093
rect 18417 12084 18429 12087
rect 18064 12056 18429 12084
rect 18417 12053 18429 12056
rect 18463 12053 18475 12087
rect 18417 12047 18475 12053
rect 18506 12044 18512 12096
rect 18564 12044 18570 12096
rect 18800 12084 18828 12260
rect 18892 12152 18920 12328
rect 20993 12325 21005 12328
rect 21039 12325 21051 12359
rect 20993 12319 21051 12325
rect 19978 12248 19984 12300
rect 20036 12288 20042 12300
rect 20073 12291 20131 12297
rect 20073 12288 20085 12291
rect 20036 12260 20085 12288
rect 20036 12248 20042 12260
rect 20073 12257 20085 12260
rect 20119 12257 20131 12291
rect 20254 12288 20260 12300
rect 20073 12251 20131 12257
rect 20246 12248 20260 12288
rect 20312 12248 20318 12300
rect 20622 12248 20628 12300
rect 20680 12248 20686 12300
rect 21008 12288 21036 12319
rect 21818 12288 21824 12300
rect 21008 12260 21824 12288
rect 20246 12229 20274 12248
rect 20211 12223 20274 12229
rect 20211 12189 20223 12223
rect 20257 12192 20274 12223
rect 20257 12189 20269 12192
rect 20211 12183 20269 12189
rect 20346 12180 20352 12232
rect 20404 12180 20410 12232
rect 20438 12180 20444 12232
rect 20496 12180 20502 12232
rect 20533 12223 20591 12229
rect 20533 12189 20545 12223
rect 20579 12220 20591 12223
rect 20640 12220 20668 12248
rect 21376 12229 21404 12260
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 22020 12297 22048 12396
rect 25225 12393 25237 12427
rect 25271 12424 25283 12427
rect 25866 12424 25872 12436
rect 25271 12396 25872 12424
rect 25271 12393 25283 12396
rect 25225 12387 25283 12393
rect 25866 12384 25872 12396
rect 25924 12384 25930 12436
rect 29638 12384 29644 12436
rect 29696 12424 29702 12436
rect 29733 12427 29791 12433
rect 29733 12424 29745 12427
rect 29696 12396 29745 12424
rect 29696 12384 29702 12396
rect 29733 12393 29745 12396
rect 29779 12393 29791 12427
rect 29733 12387 29791 12393
rect 30193 12427 30251 12433
rect 30193 12393 30205 12427
rect 30239 12424 30251 12427
rect 30282 12424 30288 12436
rect 30239 12396 30288 12424
rect 30239 12393 30251 12396
rect 30193 12387 30251 12393
rect 25038 12356 25044 12368
rect 22296 12328 25044 12356
rect 22296 12297 22324 12328
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 25317 12359 25375 12365
rect 25317 12325 25329 12359
rect 25363 12325 25375 12359
rect 25317 12319 25375 12325
rect 22005 12291 22063 12297
rect 22005 12257 22017 12291
rect 22051 12257 22063 12291
rect 22005 12251 22063 12257
rect 22281 12291 22339 12297
rect 22281 12257 22293 12291
rect 22327 12257 22339 12291
rect 25222 12288 25228 12300
rect 22281 12251 22339 12257
rect 24044 12260 25228 12288
rect 21177 12223 21235 12229
rect 21177 12220 21189 12223
rect 20579 12192 21189 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 21177 12189 21189 12192
rect 21223 12189 21235 12223
rect 21177 12183 21235 12189
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21542 12180 21548 12232
rect 21600 12180 21606 12232
rect 21634 12180 21640 12232
rect 21692 12220 21698 12232
rect 24044 12229 24072 12260
rect 25222 12248 25228 12260
rect 25280 12248 25286 12300
rect 21913 12223 21971 12229
rect 21913 12220 21925 12223
rect 21692 12192 21925 12220
rect 21692 12180 21698 12192
rect 21913 12189 21925 12192
rect 21959 12189 21971 12223
rect 21913 12183 21971 12189
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12189 24087 12223
rect 24489 12223 24547 12229
rect 24489 12220 24501 12223
rect 24029 12183 24087 12189
rect 24228 12192 24501 12220
rect 20070 12152 20076 12164
rect 18892 12124 20076 12152
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 19334 12084 19340 12096
rect 18800 12056 19340 12084
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 19426 12044 19432 12096
rect 19484 12084 19490 12096
rect 22370 12084 22376 12096
rect 19484 12056 22376 12084
rect 19484 12044 19490 12056
rect 22370 12044 22376 12056
rect 22428 12044 22434 12096
rect 24228 12093 24256 12192
rect 24489 12189 24501 12192
rect 24535 12189 24547 12223
rect 24489 12183 24547 12189
rect 24765 12223 24823 12229
rect 24765 12189 24777 12223
rect 24811 12220 24823 12223
rect 24854 12220 24860 12232
rect 24811 12192 24860 12220
rect 24811 12189 24823 12192
rect 24765 12183 24823 12189
rect 24854 12180 24860 12192
rect 24912 12180 24918 12232
rect 25041 12223 25099 12229
rect 25041 12189 25053 12223
rect 25087 12220 25099 12223
rect 25332 12220 25360 12319
rect 25087 12192 25360 12220
rect 25087 12189 25099 12192
rect 25041 12183 25099 12189
rect 25498 12180 25504 12232
rect 25556 12180 25562 12232
rect 26142 12180 26148 12232
rect 26200 12180 26206 12232
rect 27801 12223 27859 12229
rect 27801 12189 27813 12223
rect 27847 12220 27859 12223
rect 28353 12223 28411 12229
rect 28353 12220 28365 12223
rect 27847 12192 28365 12220
rect 27847 12189 27859 12192
rect 27801 12183 27859 12189
rect 28353 12189 28365 12192
rect 28399 12220 28411 12223
rect 28994 12220 29000 12232
rect 28399 12192 29000 12220
rect 28399 12189 28411 12192
rect 28353 12183 28411 12189
rect 28994 12180 29000 12192
rect 29052 12220 29058 12232
rect 29641 12223 29699 12229
rect 29641 12220 29653 12223
rect 29052 12192 29653 12220
rect 29052 12180 29058 12192
rect 29641 12189 29653 12192
rect 29687 12220 29699 12223
rect 29822 12220 29828 12232
rect 29687 12192 29828 12220
rect 29687 12189 29699 12192
rect 29641 12183 29699 12189
rect 29822 12180 29828 12192
rect 29880 12220 29886 12232
rect 30208 12220 30236 12387
rect 30282 12384 30288 12396
rect 30340 12384 30346 12436
rect 31665 12427 31723 12433
rect 31665 12424 31677 12427
rect 31404 12396 31677 12424
rect 31404 12297 31432 12396
rect 31665 12393 31677 12396
rect 31711 12424 31723 12427
rect 31754 12424 31760 12436
rect 31711 12396 31760 12424
rect 31711 12393 31723 12396
rect 31665 12387 31723 12393
rect 31754 12384 31760 12396
rect 31812 12424 31818 12436
rect 32674 12424 32680 12436
rect 31812 12396 32680 12424
rect 31812 12384 31818 12396
rect 32674 12384 32680 12396
rect 32732 12384 32738 12436
rect 31021 12291 31079 12297
rect 31021 12257 31033 12291
rect 31067 12288 31079 12291
rect 31389 12291 31447 12297
rect 31389 12288 31401 12291
rect 31067 12260 31401 12288
rect 31067 12257 31079 12260
rect 31021 12251 31079 12257
rect 31389 12257 31401 12260
rect 31435 12257 31447 12291
rect 31389 12251 31447 12257
rect 34057 12291 34115 12297
rect 34057 12257 34069 12291
rect 34103 12288 34115 12291
rect 34103 12260 34652 12288
rect 34103 12257 34115 12260
rect 34057 12251 34115 12257
rect 29880 12192 30236 12220
rect 29880 12180 29886 12192
rect 31110 12180 31116 12232
rect 31168 12180 31174 12232
rect 31202 12180 31208 12232
rect 31260 12180 31266 12232
rect 34422 12180 34428 12232
rect 34480 12180 34486 12232
rect 26160 12152 26188 12180
rect 34624 12164 34652 12260
rect 24688 12124 26188 12152
rect 24688 12093 24716 12124
rect 34606 12112 34612 12164
rect 34664 12112 34670 12164
rect 24213 12087 24271 12093
rect 24213 12053 24225 12087
rect 24259 12053 24271 12087
rect 24213 12047 24271 12053
rect 24673 12087 24731 12093
rect 24673 12053 24685 12087
rect 24719 12053 24731 12087
rect 24673 12047 24731 12053
rect 24949 12087 25007 12093
rect 24949 12053 24961 12087
rect 24995 12084 25007 12087
rect 25774 12084 25780 12096
rect 24995 12056 25780 12084
rect 24995 12053 25007 12056
rect 24949 12047 25007 12053
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 27798 12044 27804 12096
rect 27856 12084 27862 12096
rect 27893 12087 27951 12093
rect 27893 12084 27905 12087
rect 27856 12056 27905 12084
rect 27856 12044 27862 12056
rect 27893 12053 27905 12056
rect 27939 12053 27951 12087
rect 27893 12047 27951 12053
rect 28626 12044 28632 12096
rect 28684 12044 28690 12096
rect 31386 12044 31392 12096
rect 31444 12044 31450 12096
rect 1104 11994 35236 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 35236 11994
rect 1104 11920 35236 11942
rect 4614 11840 4620 11892
rect 4672 11840 4678 11892
rect 4982 11840 4988 11892
rect 5040 11880 5046 11892
rect 5169 11883 5227 11889
rect 5169 11880 5181 11883
rect 5040 11852 5181 11880
rect 5040 11840 5046 11852
rect 5169 11849 5181 11852
rect 5215 11880 5227 11883
rect 5215 11852 7512 11880
rect 5215 11849 5227 11852
rect 5169 11843 5227 11849
rect 2866 11772 2872 11824
rect 2924 11812 2930 11824
rect 3145 11815 3203 11821
rect 3145 11812 3157 11815
rect 2924 11784 3157 11812
rect 2924 11772 2930 11784
rect 3145 11781 3157 11784
rect 3191 11781 3203 11815
rect 4801 11815 4859 11821
rect 4801 11812 4813 11815
rect 4370 11784 4813 11812
rect 3145 11775 3203 11781
rect 4801 11781 4813 11784
rect 4847 11781 4859 11815
rect 4801 11775 4859 11781
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 4893 11747 4951 11753
rect 2188 11716 2728 11744
rect 2188 11704 2194 11716
rect 2700 11620 2728 11716
rect 4893 11713 4905 11747
rect 4939 11744 4951 11747
rect 5000 11744 5028 11840
rect 5350 11772 5356 11824
rect 5408 11812 5414 11824
rect 5537 11815 5595 11821
rect 5537 11812 5549 11815
rect 5408 11784 5549 11812
rect 5408 11772 5414 11784
rect 5537 11781 5549 11784
rect 5583 11781 5595 11815
rect 5537 11775 5595 11781
rect 4939 11716 5028 11744
rect 4939 11713 4951 11716
rect 4893 11707 4951 11713
rect 5994 11704 6000 11756
rect 6052 11704 6058 11756
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11744 6423 11747
rect 6454 11744 6460 11756
rect 6411 11716 6460 11744
rect 6411 11713 6423 11716
rect 6365 11707 6423 11713
rect 2774 11636 2780 11688
rect 2832 11676 2838 11688
rect 2869 11679 2927 11685
rect 2869 11676 2881 11679
rect 2832 11648 2881 11676
rect 2832 11636 2838 11648
rect 2869 11645 2881 11648
rect 2915 11645 2927 11679
rect 3786 11676 3792 11688
rect 2869 11639 2927 11645
rect 2976 11648 3792 11676
rect 2682 11568 2688 11620
rect 2740 11608 2746 11620
rect 2976 11608 3004 11648
rect 3786 11636 3792 11648
rect 3844 11676 3850 11688
rect 6380 11676 6408 11707
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 3844 11648 6408 11676
rect 7484 11676 7512 11852
rect 7558 11840 7564 11892
rect 7616 11840 7622 11892
rect 8202 11840 8208 11892
rect 8260 11840 8266 11892
rect 8389 11883 8447 11889
rect 8389 11849 8401 11883
rect 8435 11880 8447 11883
rect 8435 11852 8800 11880
rect 8435 11849 8447 11852
rect 8389 11843 8447 11849
rect 7576 11744 7604 11840
rect 8220 11812 8248 11840
rect 8772 11821 8800 11852
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 8904 11852 10548 11880
rect 8904 11840 8910 11852
rect 8757 11815 8815 11821
rect 8220 11784 8524 11812
rect 8496 11753 8524 11784
rect 8757 11781 8769 11815
rect 8803 11781 8815 11815
rect 10413 11815 10471 11821
rect 10413 11812 10425 11815
rect 9982 11784 10425 11812
rect 8757 11775 8815 11781
rect 10413 11781 10425 11784
rect 10459 11781 10471 11815
rect 10413 11775 10471 11781
rect 10520 11753 10548 11852
rect 11974 11840 11980 11892
rect 12032 11880 12038 11892
rect 12529 11883 12587 11889
rect 12529 11880 12541 11883
rect 12032 11852 12541 11880
rect 12032 11840 12038 11852
rect 12529 11849 12541 11852
rect 12575 11849 12587 11883
rect 12529 11843 12587 11849
rect 8205 11747 8263 11753
rect 8205 11744 8217 11747
rect 7576 11716 8217 11744
rect 8205 11713 8217 11716
rect 8251 11713 8263 11747
rect 8205 11707 8263 11713
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 8481 11707 8539 11713
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11744 10563 11747
rect 10594 11744 10600 11756
rect 10551 11716 10600 11744
rect 10551 11713 10563 11716
rect 10505 11707 10563 11713
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 10689 11747 10747 11753
rect 10689 11713 10701 11747
rect 10735 11713 10747 11747
rect 12544 11744 12572 11843
rect 12802 11840 12808 11892
rect 12860 11840 12866 11892
rect 13538 11840 13544 11892
rect 13596 11840 13602 11892
rect 13906 11840 13912 11892
rect 13964 11880 13970 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 13964 11852 14289 11880
rect 13964 11840 13970 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 15102 11840 15108 11892
rect 15160 11880 15166 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 15160 11852 15209 11880
rect 15160 11840 15166 11852
rect 15197 11849 15209 11852
rect 15243 11849 15255 11883
rect 15197 11843 15255 11849
rect 15562 11840 15568 11892
rect 15620 11840 15626 11892
rect 16114 11840 16120 11892
rect 16172 11840 16178 11892
rect 18506 11880 18512 11892
rect 17328 11852 18512 11880
rect 12713 11815 12771 11821
rect 12713 11781 12725 11815
rect 12759 11812 12771 11815
rect 12820 11812 12848 11840
rect 12759 11784 12848 11812
rect 13556 11812 13584 11840
rect 13556 11784 14688 11812
rect 12759 11781 12771 11784
rect 12713 11775 12771 11781
rect 12805 11747 12863 11753
rect 12805 11744 12817 11747
rect 12544 11716 12817 11744
rect 10689 11707 10747 11713
rect 12805 11713 12817 11716
rect 12851 11713 12863 11747
rect 12805 11707 12863 11713
rect 8110 11676 8116 11688
rect 7484 11648 8116 11676
rect 3844 11636 3850 11648
rect 8110 11636 8116 11648
rect 8168 11636 8174 11688
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11676 10287 11679
rect 10704 11676 10732 11707
rect 12986 11704 12992 11756
rect 13044 11704 13050 11756
rect 10275 11648 10732 11676
rect 11241 11679 11299 11685
rect 10275 11645 10287 11648
rect 10229 11639 10287 11645
rect 11241 11645 11253 11679
rect 11287 11676 11299 11679
rect 13556 11676 13584 11784
rect 13906 11704 13912 11756
rect 13964 11744 13970 11756
rect 14660 11753 14688 11784
rect 14826 11772 14832 11824
rect 14884 11772 14890 11824
rect 16132 11812 16160 11840
rect 15856 11784 17172 11812
rect 14461 11747 14519 11753
rect 14461 11744 14473 11747
rect 13964 11716 14473 11744
rect 13964 11704 13970 11716
rect 14461 11713 14473 11716
rect 14507 11713 14519 11747
rect 14461 11707 14519 11713
rect 14645 11747 14703 11753
rect 14645 11713 14657 11747
rect 14691 11713 14703 11747
rect 14645 11707 14703 11713
rect 15194 11704 15200 11756
rect 15252 11704 15258 11756
rect 15286 11704 15292 11756
rect 15344 11744 15350 11756
rect 15856 11753 15884 11784
rect 15749 11747 15807 11753
rect 15749 11744 15761 11747
rect 15344 11716 15761 11744
rect 15344 11704 15350 11716
rect 15749 11713 15761 11716
rect 15795 11713 15807 11747
rect 15749 11707 15807 11713
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11713 15899 11747
rect 15841 11707 15899 11713
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 11287 11648 13584 11676
rect 15212 11676 15240 11704
rect 16040 11676 16068 11707
rect 16114 11704 16120 11756
rect 16172 11744 16178 11756
rect 16574 11744 16580 11756
rect 16172 11716 16580 11744
rect 16172 11704 16178 11716
rect 16574 11704 16580 11716
rect 16632 11704 16638 11756
rect 16850 11704 16856 11756
rect 16908 11704 16914 11756
rect 17144 11753 17172 11784
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 17129 11747 17187 11753
rect 17129 11713 17141 11747
rect 17175 11744 17187 11747
rect 17218 11744 17224 11756
rect 17175 11716 17224 11744
rect 17175 11713 17187 11716
rect 17129 11707 17187 11713
rect 16482 11676 16488 11688
rect 15212 11648 16488 11676
rect 11287 11645 11299 11648
rect 11241 11639 11299 11645
rect 16482 11636 16488 11648
rect 16540 11636 16546 11688
rect 17052 11676 17080 11707
rect 17218 11704 17224 11716
rect 17276 11704 17282 11756
rect 17328 11753 17356 11852
rect 18506 11840 18512 11852
rect 18564 11840 18570 11892
rect 18874 11880 18880 11892
rect 18708 11852 18880 11880
rect 18138 11772 18144 11824
rect 18196 11812 18202 11824
rect 18196 11784 18276 11812
rect 18196 11772 18202 11784
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11744 17463 11747
rect 17770 11744 17776 11756
rect 17451 11716 17776 11744
rect 17451 11713 17463 11716
rect 17405 11707 17463 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 18248 11746 18276 11784
rect 18708 11753 18736 11852
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 19058 11840 19064 11892
rect 19116 11880 19122 11892
rect 19116 11852 19334 11880
rect 19116 11840 19122 11852
rect 19306 11812 19334 11852
rect 19426 11840 19432 11892
rect 19484 11840 19490 11892
rect 20272 11852 20484 11880
rect 20272 11812 20300 11852
rect 18800 11784 19012 11812
rect 19306 11784 20300 11812
rect 18325 11747 18383 11753
rect 18325 11746 18337 11747
rect 18248 11718 18337 11746
rect 18325 11713 18337 11718
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 18693 11747 18751 11753
rect 18693 11713 18705 11747
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 18141 11679 18199 11685
rect 17052 11648 17632 11676
rect 2740 11580 3004 11608
rect 2740 11568 2746 11580
rect 9858 11568 9864 11620
rect 9916 11568 9922 11620
rect 2222 11500 2228 11552
rect 2280 11500 2286 11552
rect 6178 11500 6184 11552
rect 6236 11500 6242 11552
rect 9876 11540 9904 11568
rect 17604 11552 17632 11648
rect 18141 11645 18153 11679
rect 18187 11645 18199 11679
rect 18141 11639 18199 11645
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 18417 11679 18475 11685
rect 18417 11645 18429 11679
rect 18463 11676 18475 11679
rect 18506 11676 18512 11688
rect 18463 11648 18512 11676
rect 18463 11645 18475 11648
rect 18417 11639 18475 11645
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 9876 11512 12173 11540
rect 12161 11509 12173 11512
rect 12207 11540 12219 11543
rect 12986 11540 12992 11552
rect 12207 11512 12992 11540
rect 12207 11509 12219 11512
rect 12161 11503 12219 11509
rect 12986 11500 12992 11512
rect 13044 11500 13050 11552
rect 16298 11500 16304 11552
rect 16356 11500 16362 11552
rect 17586 11500 17592 11552
rect 17644 11500 17650 11552
rect 18156 11540 18184 11639
rect 18248 11608 18276 11639
rect 18506 11636 18512 11648
rect 18564 11636 18570 11688
rect 18601 11679 18659 11685
rect 18601 11645 18613 11679
rect 18647 11676 18659 11679
rect 18800 11676 18828 11784
rect 18874 11704 18880 11756
rect 18932 11704 18938 11756
rect 18984 11753 19012 11784
rect 18969 11747 19027 11753
rect 18969 11713 18981 11747
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 19061 11747 19119 11753
rect 19061 11713 19073 11747
rect 19107 11744 19119 11747
rect 19107 11716 19196 11744
rect 19107 11713 19119 11716
rect 19061 11707 19119 11713
rect 18647 11648 18828 11676
rect 18647 11645 18659 11648
rect 18601 11639 18659 11645
rect 18966 11608 18972 11620
rect 18248 11580 18972 11608
rect 18966 11568 18972 11580
rect 19024 11568 19030 11620
rect 19168 11608 19196 11716
rect 19242 11704 19248 11756
rect 19300 11704 19306 11756
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 19392 11716 19717 11744
rect 19392 11704 19398 11716
rect 19705 11713 19717 11716
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 19794 11704 19800 11756
rect 19852 11704 19858 11756
rect 19886 11704 19892 11756
rect 19944 11753 19950 11756
rect 19944 11747 19993 11753
rect 19944 11713 19947 11747
rect 19981 11713 19993 11747
rect 19944 11707 19993 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 19944 11704 19950 11707
rect 19521 11611 19579 11617
rect 19521 11608 19533 11611
rect 19168 11580 19533 11608
rect 19521 11577 19533 11580
rect 19567 11577 19579 11611
rect 19521 11571 19579 11577
rect 20088 11552 20116 11707
rect 20162 11704 20168 11756
rect 20220 11704 20226 11756
rect 20349 11747 20407 11753
rect 20349 11713 20361 11747
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 20364 11676 20392 11707
rect 20180 11648 20392 11676
rect 20180 11620 20208 11648
rect 20162 11568 20168 11620
rect 20220 11568 20226 11620
rect 20456 11608 20484 11852
rect 20622 11840 20628 11892
rect 20680 11840 20686 11892
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 21634 11880 21640 11892
rect 21048 11852 21640 11880
rect 21048 11840 21054 11852
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 23566 11840 23572 11892
rect 23624 11880 23630 11892
rect 23661 11883 23719 11889
rect 23661 11880 23673 11883
rect 23624 11852 23673 11880
rect 23624 11840 23630 11852
rect 23661 11849 23673 11852
rect 23707 11849 23719 11883
rect 23661 11843 23719 11849
rect 23845 11883 23903 11889
rect 23845 11849 23857 11883
rect 23891 11880 23903 11883
rect 24210 11880 24216 11892
rect 23891 11852 24216 11880
rect 23891 11849 23903 11852
rect 23845 11843 23903 11849
rect 24210 11840 24216 11852
rect 24268 11840 24274 11892
rect 24486 11840 24492 11892
rect 24544 11840 24550 11892
rect 24578 11840 24584 11892
rect 24636 11840 24642 11892
rect 25590 11840 25596 11892
rect 25648 11840 25654 11892
rect 28994 11840 29000 11892
rect 29052 11840 29058 11892
rect 32401 11883 32459 11889
rect 32401 11849 32413 11883
rect 32447 11880 32459 11883
rect 33042 11880 33048 11892
rect 32447 11852 33048 11880
rect 32447 11849 32459 11852
rect 32401 11843 32459 11849
rect 20640 11812 20668 11840
rect 20640 11784 21496 11812
rect 20530 11704 20536 11756
rect 20588 11744 20594 11756
rect 20625 11747 20683 11753
rect 20625 11744 20637 11747
rect 20588 11716 20637 11744
rect 20588 11704 20594 11716
rect 20625 11713 20637 11716
rect 20671 11713 20683 11747
rect 20625 11707 20683 11713
rect 20640 11676 20668 11707
rect 20990 11704 20996 11756
rect 21048 11704 21054 11756
rect 21174 11704 21180 11756
rect 21232 11704 21238 11756
rect 21468 11753 21496 11784
rect 23106 11772 23112 11824
rect 23164 11812 23170 11824
rect 23477 11815 23535 11821
rect 23477 11812 23489 11815
rect 23164 11784 23489 11812
rect 23164 11772 23170 11784
rect 23477 11781 23489 11784
rect 23523 11781 23535 11815
rect 24673 11815 24731 11821
rect 24673 11812 24685 11815
rect 23477 11775 23535 11781
rect 24136 11784 24685 11812
rect 24136 11756 24164 11784
rect 24673 11781 24685 11784
rect 24719 11781 24731 11815
rect 24673 11775 24731 11781
rect 21453 11747 21511 11753
rect 21453 11713 21465 11747
rect 21499 11713 21511 11747
rect 24029 11747 24087 11753
rect 24029 11744 24041 11747
rect 21453 11707 21511 11713
rect 23676 11716 24041 11744
rect 23676 11688 23704 11716
rect 24029 11713 24041 11716
rect 24075 11713 24087 11747
rect 24029 11707 24087 11713
rect 21269 11679 21327 11685
rect 21269 11676 21281 11679
rect 20640 11648 21281 11676
rect 21269 11645 21281 11648
rect 21315 11645 21327 11679
rect 21269 11639 21327 11645
rect 23658 11636 23664 11688
rect 23716 11636 23722 11688
rect 24044 11676 24072 11707
rect 24118 11704 24124 11756
rect 24176 11704 24182 11756
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24394 11744 24400 11756
rect 24351 11716 24400 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24394 11704 24400 11716
rect 24452 11744 24458 11756
rect 24581 11747 24639 11753
rect 24581 11744 24593 11747
rect 24452 11716 24593 11744
rect 24452 11704 24458 11716
rect 24581 11713 24593 11716
rect 24627 11713 24639 11747
rect 24581 11707 24639 11713
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11713 24915 11747
rect 24857 11707 24915 11713
rect 24872 11676 24900 11707
rect 25130 11704 25136 11756
rect 25188 11744 25194 11756
rect 25317 11747 25375 11753
rect 25317 11744 25329 11747
rect 25188 11716 25329 11744
rect 25188 11704 25194 11716
rect 25317 11713 25329 11716
rect 25363 11713 25375 11747
rect 25317 11707 25375 11713
rect 25501 11747 25559 11753
rect 25501 11713 25513 11747
rect 25547 11744 25559 11747
rect 25608 11744 25636 11840
rect 26329 11815 26387 11821
rect 26329 11812 26341 11815
rect 25792 11784 26341 11812
rect 25792 11753 25820 11784
rect 26329 11781 26341 11784
rect 26375 11781 26387 11815
rect 26329 11775 26387 11781
rect 28721 11815 28779 11821
rect 28721 11781 28733 11815
rect 28767 11812 28779 11815
rect 29012 11812 29040 11840
rect 28767 11784 29040 11812
rect 28767 11781 28779 11784
rect 28721 11775 28779 11781
rect 30098 11772 30104 11824
rect 30156 11772 30162 11824
rect 30650 11772 30656 11824
rect 30708 11812 30714 11824
rect 31202 11812 31208 11824
rect 30708 11784 31208 11812
rect 30708 11772 30714 11784
rect 31202 11772 31208 11784
rect 31260 11812 31266 11824
rect 31260 11784 31616 11812
rect 31260 11772 31266 11784
rect 25547 11716 25636 11744
rect 25777 11747 25835 11753
rect 25547 11713 25559 11716
rect 25501 11707 25559 11713
rect 25777 11713 25789 11747
rect 25823 11713 25835 11747
rect 25777 11707 25835 11713
rect 26237 11747 26295 11753
rect 26237 11713 26249 11747
rect 26283 11713 26295 11747
rect 26237 11707 26295 11713
rect 26421 11747 26479 11753
rect 26421 11713 26433 11747
rect 26467 11744 26479 11747
rect 26510 11744 26516 11756
rect 26467 11716 26516 11744
rect 26467 11713 26479 11716
rect 26421 11707 26479 11713
rect 24044 11648 24900 11676
rect 21177 11611 21235 11617
rect 21177 11608 21189 11611
rect 20456 11580 21189 11608
rect 21177 11577 21189 11580
rect 21223 11608 21235 11611
rect 23014 11608 23020 11620
rect 21223 11580 23020 11608
rect 21223 11577 21235 11580
rect 21177 11571 21235 11577
rect 23014 11568 23020 11580
rect 23072 11568 23078 11620
rect 25148 11617 25176 11704
rect 25409 11679 25467 11685
rect 25409 11645 25421 11679
rect 25455 11676 25467 11679
rect 25685 11679 25743 11685
rect 25685 11676 25697 11679
rect 25455 11648 25697 11676
rect 25455 11645 25467 11648
rect 25409 11639 25467 11645
rect 25685 11645 25697 11648
rect 25731 11645 25743 11679
rect 25685 11639 25743 11645
rect 26050 11636 26056 11688
rect 26108 11676 26114 11688
rect 26252 11676 26280 11707
rect 26510 11704 26516 11716
rect 26568 11744 26574 11756
rect 26697 11747 26755 11753
rect 26697 11744 26709 11747
rect 26568 11716 26709 11744
rect 26568 11704 26574 11716
rect 26697 11713 26709 11716
rect 26743 11713 26755 11747
rect 26697 11707 26755 11713
rect 26973 11747 27031 11753
rect 26973 11713 26985 11747
rect 27019 11744 27031 11747
rect 28074 11744 28080 11756
rect 27019 11716 28080 11744
rect 27019 11713 27031 11716
rect 26973 11707 27031 11713
rect 28074 11704 28080 11716
rect 28132 11704 28138 11756
rect 30837 11747 30895 11753
rect 30837 11744 30849 11747
rect 30576 11716 30849 11744
rect 30576 11688 30604 11716
rect 30837 11713 30849 11716
rect 30883 11713 30895 11747
rect 30837 11707 30895 11713
rect 31110 11704 31116 11756
rect 31168 11744 31174 11756
rect 31588 11753 31616 11784
rect 32508 11756 32536 11852
rect 33042 11840 33048 11852
rect 33100 11840 33106 11892
rect 34425 11815 34483 11821
rect 34425 11812 34437 11815
rect 33994 11784 34437 11812
rect 34425 11781 34437 11784
rect 34471 11781 34483 11815
rect 34425 11775 34483 11781
rect 31481 11747 31539 11753
rect 31481 11744 31493 11747
rect 31168 11716 31493 11744
rect 31168 11704 31174 11716
rect 31481 11713 31493 11716
rect 31527 11713 31539 11747
rect 31481 11707 31539 11713
rect 31573 11747 31631 11753
rect 31573 11713 31585 11747
rect 31619 11713 31631 11747
rect 31573 11707 31631 11713
rect 31754 11704 31760 11756
rect 31812 11704 31818 11756
rect 32490 11704 32496 11756
rect 32548 11704 32554 11756
rect 34514 11704 34520 11756
rect 34572 11744 34578 11756
rect 34885 11747 34943 11753
rect 34885 11744 34897 11747
rect 34572 11716 34897 11744
rect 34572 11704 34578 11716
rect 34885 11713 34897 11716
rect 34931 11713 34943 11747
rect 34885 11707 34943 11713
rect 26108 11648 26280 11676
rect 26108 11636 26114 11648
rect 26786 11636 26792 11688
rect 26844 11676 26850 11688
rect 28626 11676 28632 11688
rect 26844 11648 28632 11676
rect 26844 11636 26850 11648
rect 28626 11636 28632 11648
rect 28684 11676 28690 11688
rect 28813 11679 28871 11685
rect 28813 11676 28825 11679
rect 28684 11648 28825 11676
rect 28684 11636 28690 11648
rect 28813 11645 28825 11648
rect 28859 11645 28871 11679
rect 29089 11679 29147 11685
rect 29089 11676 29101 11679
rect 28813 11639 28871 11645
rect 28920 11648 29101 11676
rect 25133 11611 25191 11617
rect 25133 11608 25145 11611
rect 23584 11580 25145 11608
rect 18782 11540 18788 11552
rect 18156 11512 18788 11540
rect 18782 11500 18788 11512
rect 18840 11540 18846 11552
rect 20070 11540 20076 11552
rect 18840 11512 20076 11540
rect 18840 11500 18846 11512
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20180 11540 20208 11568
rect 20898 11540 20904 11552
rect 20180 11512 20904 11540
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 21266 11500 21272 11552
rect 21324 11540 21330 11552
rect 21637 11543 21695 11549
rect 21637 11540 21649 11543
rect 21324 11512 21649 11540
rect 21324 11500 21330 11512
rect 21637 11509 21649 11512
rect 21683 11509 21695 11543
rect 21637 11503 21695 11509
rect 21818 11500 21824 11552
rect 21876 11540 21882 11552
rect 23584 11540 23612 11580
rect 25133 11577 25145 11580
rect 25179 11577 25191 11611
rect 28920 11608 28948 11648
rect 29089 11645 29101 11648
rect 29135 11645 29147 11679
rect 29089 11639 29147 11645
rect 30558 11636 30564 11688
rect 30616 11636 30622 11688
rect 30929 11679 30987 11685
rect 30929 11645 30941 11679
rect 30975 11676 30987 11679
rect 31297 11679 31355 11685
rect 31297 11676 31309 11679
rect 30975 11648 31309 11676
rect 30975 11645 30987 11648
rect 30929 11639 30987 11645
rect 31297 11645 31309 11648
rect 31343 11645 31355 11679
rect 31297 11639 31355 11645
rect 32766 11636 32772 11688
rect 32824 11636 32830 11688
rect 25133 11571 25191 11577
rect 26068 11580 28948 11608
rect 31220 11580 31524 11608
rect 21876 11512 23612 11540
rect 23661 11543 23719 11549
rect 21876 11500 21882 11512
rect 23661 11509 23673 11543
rect 23707 11540 23719 11543
rect 24210 11540 24216 11552
rect 23707 11512 24216 11540
rect 23707 11509 23719 11512
rect 23661 11503 23719 11509
rect 24210 11500 24216 11512
rect 24268 11500 24274 11552
rect 25038 11500 25044 11552
rect 25096 11540 25102 11552
rect 26068 11540 26096 11580
rect 25096 11512 26096 11540
rect 25096 11500 25102 11512
rect 26142 11500 26148 11552
rect 26200 11500 26206 11552
rect 31220 11549 31248 11580
rect 31205 11543 31263 11549
rect 31205 11509 31217 11543
rect 31251 11509 31263 11543
rect 31496 11540 31524 11580
rect 31662 11568 31668 11620
rect 31720 11568 31726 11620
rect 32858 11540 32864 11552
rect 31496 11512 32864 11540
rect 31205 11503 31263 11509
rect 32858 11500 32864 11512
rect 32916 11500 32922 11552
rect 34238 11500 34244 11552
rect 34296 11500 34302 11552
rect 1104 11450 35248 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 35248 11450
rect 1104 11376 35248 11398
rect 2774 11296 2780 11348
rect 2832 11296 2838 11348
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 5442 11336 5448 11348
rect 3191 11308 5448 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6178 11296 6184 11348
rect 6236 11296 6242 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 15381 11339 15439 11345
rect 15381 11336 15393 11339
rect 13044 11308 15393 11336
rect 13044 11296 13050 11308
rect 15381 11305 15393 11308
rect 15427 11305 15439 11339
rect 15381 11299 15439 11305
rect 2792 11268 2820 11296
rect 3510 11268 3516 11280
rect 2792 11240 3516 11268
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 4525 11271 4583 11277
rect 4525 11237 4537 11271
rect 4571 11268 4583 11271
rect 4982 11268 4988 11280
rect 4571 11240 4988 11268
rect 4571 11237 4583 11240
rect 4525 11231 4583 11237
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4540 11132 4568 11231
rect 4982 11228 4988 11240
rect 5040 11228 5046 11280
rect 5350 11160 5356 11212
rect 5408 11160 5414 11212
rect 6196 11200 6224 11296
rect 15396 11268 15424 11299
rect 15746 11296 15752 11348
rect 15804 11296 15810 11348
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16117 11339 16175 11345
rect 16117 11336 16129 11339
rect 15988 11308 16129 11336
rect 15988 11296 15994 11308
rect 16117 11305 16129 11308
rect 16163 11305 16175 11339
rect 16117 11299 16175 11305
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 17129 11339 17187 11345
rect 17129 11336 17141 11339
rect 16540 11308 17141 11336
rect 16540 11296 16546 11308
rect 17129 11305 17141 11308
rect 17175 11305 17187 11339
rect 17129 11299 17187 11305
rect 15838 11268 15844 11280
rect 15396 11240 15844 11268
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 17144 11268 17172 11299
rect 17678 11296 17684 11348
rect 17736 11296 17742 11348
rect 17773 11339 17831 11345
rect 17773 11305 17785 11339
rect 17819 11336 17831 11339
rect 17862 11336 17868 11348
rect 17819 11308 17868 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18141 11339 18199 11345
rect 18141 11336 18153 11339
rect 18104 11308 18153 11336
rect 18104 11296 18110 11308
rect 18141 11305 18153 11308
rect 18187 11305 18199 11339
rect 18141 11299 18199 11305
rect 18601 11339 18659 11345
rect 18601 11305 18613 11339
rect 18647 11336 18659 11339
rect 18874 11336 18880 11348
rect 18647 11308 18880 11336
rect 18647 11305 18659 11308
rect 18601 11299 18659 11305
rect 18874 11296 18880 11308
rect 18932 11296 18938 11348
rect 19306 11308 19472 11336
rect 17543 11271 17601 11277
rect 17543 11268 17555 11271
rect 17144 11240 17555 11268
rect 17543 11237 17555 11240
rect 17589 11237 17601 11271
rect 17696 11268 17724 11296
rect 18506 11268 18512 11280
rect 17696 11240 18512 11268
rect 17543 11231 17601 11237
rect 18506 11228 18512 11240
rect 18564 11228 18570 11280
rect 19306 11268 19334 11308
rect 18800 11240 19334 11268
rect 6825 11203 6883 11209
rect 6825 11200 6837 11203
rect 6196 11172 6837 11200
rect 6825 11169 6837 11172
rect 6871 11169 6883 11203
rect 6825 11163 6883 11169
rect 8297 11203 8355 11209
rect 8297 11169 8309 11203
rect 8343 11200 8355 11203
rect 11057 11203 11115 11209
rect 8343 11172 8984 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 4203 11104 4568 11132
rect 5368 11132 5396 11160
rect 8956 11141 8984 11172
rect 11057 11169 11069 11203
rect 11103 11200 11115 11203
rect 11146 11200 11152 11212
rect 11103 11172 11152 11200
rect 11103 11169 11115 11172
rect 11057 11163 11115 11169
rect 11146 11160 11152 11172
rect 11204 11200 11210 11212
rect 18800 11200 18828 11240
rect 11204 11172 18828 11200
rect 19444 11200 19472 11308
rect 20438 11296 20444 11348
rect 20496 11336 20502 11348
rect 20901 11339 20959 11345
rect 20901 11336 20913 11339
rect 20496 11308 20913 11336
rect 20496 11296 20502 11308
rect 20901 11305 20913 11308
rect 20947 11305 20959 11339
rect 20901 11299 20959 11305
rect 21174 11296 21180 11348
rect 21232 11336 21238 11348
rect 21269 11339 21327 11345
rect 21269 11336 21281 11339
rect 21232 11308 21281 11336
rect 21232 11296 21238 11308
rect 21269 11305 21281 11308
rect 21315 11305 21327 11339
rect 21269 11299 21327 11305
rect 21542 11296 21548 11348
rect 21600 11336 21606 11348
rect 25225 11339 25283 11345
rect 21600 11308 25084 11336
rect 21600 11296 21606 11308
rect 22066 11240 23796 11268
rect 22066 11200 22094 11240
rect 19444 11172 22094 11200
rect 22204 11172 23336 11200
rect 11204 11160 11210 11172
rect 6549 11135 6607 11141
rect 6549 11132 6561 11135
rect 5368 11104 6561 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 6549 11101 6561 11104
rect 6595 11101 6607 11135
rect 6549 11095 6607 11101
rect 8573 11135 8631 11141
rect 8573 11101 8585 11135
rect 8619 11132 8631 11135
rect 8941 11135 8999 11141
rect 8619 11104 8708 11132
rect 8619 11101 8631 11104
rect 8573 11095 8631 11101
rect 8680 11076 8708 11104
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 12618 11132 12624 11144
rect 9815 11104 12624 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 17405 11135 17463 11141
rect 17405 11132 17417 11135
rect 17236 11104 17417 11132
rect 1578 11024 1584 11076
rect 1636 11064 1642 11076
rect 1673 11067 1731 11073
rect 1673 11064 1685 11067
rect 1636 11036 1685 11064
rect 1636 11024 1642 11036
rect 1673 11033 1685 11036
rect 1719 11033 1731 11067
rect 1673 11027 1731 11033
rect 2222 11024 2228 11076
rect 2280 11024 2286 11076
rect 4065 11067 4123 11073
rect 4065 11033 4077 11067
rect 4111 11064 4123 11067
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 4111 11036 4200 11064
rect 8050 11036 8493 11064
rect 4111 11033 4123 11036
rect 4065 11027 4123 11033
rect 4172 11008 4200 11036
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 8481 11027 8539 11033
rect 8662 11024 8668 11076
rect 8720 11024 8726 11076
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 15712 11036 16957 11064
rect 15712 11024 15718 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 16945 11027 17003 11033
rect 4154 10956 4160 11008
rect 4212 10956 4218 11008
rect 10686 10956 10692 11008
rect 10744 10956 10750 11008
rect 16960 10996 16988 11027
rect 17126 11024 17132 11076
rect 17184 11073 17190 11076
rect 17184 11067 17203 11073
rect 17191 11033 17203 11067
rect 17184 11027 17203 11033
rect 17184 11024 17190 11027
rect 17236 10996 17264 11104
rect 17405 11101 17417 11104
rect 17451 11101 17463 11135
rect 17405 11095 17463 11101
rect 17494 11092 17500 11144
rect 17552 11092 17558 11144
rect 17586 11092 17592 11144
rect 17644 11132 17650 11144
rect 17681 11135 17739 11141
rect 17681 11132 17693 11135
rect 17644 11104 17693 11132
rect 17644 11092 17650 11104
rect 17681 11101 17693 11104
rect 17727 11101 17739 11135
rect 17681 11095 17739 11101
rect 17957 11135 18015 11141
rect 17957 11101 17969 11135
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 18049 11135 18107 11141
rect 18049 11101 18061 11135
rect 18095 11132 18107 11135
rect 18138 11132 18144 11144
rect 18095 11104 18144 11132
rect 18095 11101 18107 11104
rect 18049 11095 18107 11101
rect 17512 11064 17540 11092
rect 17972 11064 18000 11095
rect 18138 11092 18144 11104
rect 18196 11092 18202 11144
rect 18230 11092 18236 11144
rect 18288 11092 18294 11144
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 18414 11092 18420 11144
rect 18472 11092 18478 11144
rect 18506 11092 18512 11144
rect 18564 11132 18570 11144
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 18564 11104 18889 11132
rect 18564 11092 18570 11104
rect 18877 11101 18889 11104
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 18966 11092 18972 11144
rect 19024 11132 19030 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 19024 11104 19257 11132
rect 19024 11092 19030 11104
rect 19245 11101 19257 11104
rect 19291 11132 19303 11135
rect 19334 11132 19340 11144
rect 19291 11104 19340 11132
rect 19291 11101 19303 11104
rect 19245 11095 19303 11101
rect 19334 11092 19340 11104
rect 19392 11092 19398 11144
rect 19794 11092 19800 11144
rect 19852 11092 19858 11144
rect 19886 11092 19892 11144
rect 19944 11132 19950 11144
rect 19981 11135 20039 11141
rect 19981 11132 19993 11135
rect 19944 11104 19993 11132
rect 19944 11092 19950 11104
rect 19981 11101 19993 11104
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 20349 11135 20407 11141
rect 20349 11132 20361 11135
rect 20128 11104 20361 11132
rect 20128 11092 20134 11104
rect 20349 11101 20361 11104
rect 20395 11101 20407 11135
rect 20349 11095 20407 11101
rect 20806 11092 20812 11144
rect 20864 11092 20870 11144
rect 20898 11092 20904 11144
rect 20956 11132 20962 11144
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 20956 11104 21097 11132
rect 20956 11092 20962 11104
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 21358 11092 21364 11144
rect 21416 11132 21422 11144
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21416 11104 21649 11132
rect 21416 11092 21422 11104
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 18248 11064 18276 11092
rect 17512 11036 18000 11064
rect 18064 11036 18276 11064
rect 18340 11064 18368 11092
rect 19812 11064 19840 11092
rect 20625 11067 20683 11073
rect 18340 11036 20392 11064
rect 16960 10968 17264 10996
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 17770 10996 17776 11008
rect 17359 10968 17776 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 17770 10956 17776 10968
rect 17828 10956 17834 11008
rect 17957 10999 18015 11005
rect 17957 10965 17969 10999
rect 18003 10996 18015 10999
rect 18064 10996 18092 11036
rect 20364 11008 20392 11036
rect 20625 11033 20637 11067
rect 20671 11064 20683 11067
rect 22204 11064 22232 11172
rect 22554 11092 22560 11144
rect 22612 11132 22618 11144
rect 22741 11135 22799 11141
rect 22741 11132 22753 11135
rect 22612 11104 22753 11132
rect 22612 11092 22618 11104
rect 22741 11101 22753 11104
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 23106 11092 23112 11144
rect 23164 11132 23170 11144
rect 23201 11135 23259 11141
rect 23201 11132 23213 11135
rect 23164 11104 23213 11132
rect 23164 11092 23170 11104
rect 23201 11101 23213 11104
rect 23247 11101 23259 11135
rect 23308 11132 23336 11172
rect 23308 11126 23520 11132
rect 23658 11126 23664 11144
rect 23308 11104 23664 11126
rect 23201 11095 23259 11101
rect 23492 11098 23664 11104
rect 23658 11092 23664 11098
rect 23716 11092 23722 11144
rect 23768 11132 23796 11240
rect 23842 11228 23848 11280
rect 23900 11228 23906 11280
rect 24118 11228 24124 11280
rect 24176 11268 24182 11280
rect 24213 11271 24271 11277
rect 24213 11268 24225 11271
rect 24176 11240 24225 11268
rect 24176 11228 24182 11240
rect 24213 11237 24225 11240
rect 24259 11237 24271 11271
rect 25056 11268 25084 11308
rect 25225 11305 25237 11339
rect 25271 11336 25283 11339
rect 25590 11336 25596 11348
rect 25271 11308 25596 11336
rect 25271 11305 25283 11308
rect 25225 11299 25283 11305
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 26142 11296 26148 11348
rect 26200 11296 26206 11348
rect 29822 11296 29828 11348
rect 29880 11296 29886 11348
rect 30098 11296 30104 11348
rect 30156 11296 30162 11348
rect 30558 11296 30564 11348
rect 30616 11296 30622 11348
rect 30650 11296 30656 11348
rect 30708 11336 30714 11348
rect 30745 11339 30803 11345
rect 30745 11336 30757 11339
rect 30708 11308 30757 11336
rect 30708 11296 30714 11308
rect 30745 11305 30757 11308
rect 30791 11305 30803 11339
rect 30745 11299 30803 11305
rect 31205 11339 31263 11345
rect 31205 11305 31217 11339
rect 31251 11336 31263 11339
rect 31294 11336 31300 11348
rect 31251 11308 31300 11336
rect 31251 11305 31263 11308
rect 31205 11299 31263 11305
rect 31294 11296 31300 11308
rect 31352 11296 31358 11348
rect 31386 11296 31392 11348
rect 31444 11296 31450 11348
rect 31849 11339 31907 11345
rect 31849 11305 31861 11339
rect 31895 11336 31907 11339
rect 32766 11336 32772 11348
rect 31895 11308 32772 11336
rect 31895 11305 31907 11308
rect 31849 11299 31907 11305
rect 32766 11296 32772 11308
rect 32824 11296 32830 11348
rect 32858 11296 32864 11348
rect 32916 11296 32922 11348
rect 34514 11296 34520 11348
rect 34572 11296 34578 11348
rect 26050 11268 26056 11280
rect 25056 11240 26056 11268
rect 24213 11231 24271 11237
rect 26050 11228 26056 11240
rect 26108 11228 26114 11280
rect 26160 11200 26188 11296
rect 27065 11203 27123 11209
rect 27065 11200 27077 11203
rect 26160 11172 27077 11200
rect 27065 11169 27077 11172
rect 27111 11169 27123 11203
rect 27065 11163 27123 11169
rect 28537 11203 28595 11209
rect 28537 11169 28549 11203
rect 28583 11169 28595 11203
rect 28537 11163 28595 11169
rect 26605 11135 26663 11141
rect 26605 11132 26617 11135
rect 23768 11104 26617 11132
rect 26605 11101 26617 11104
rect 26651 11132 26663 11135
rect 26786 11132 26792 11144
rect 26651 11104 26792 11132
rect 26651 11101 26663 11104
rect 26605 11095 26663 11101
rect 26786 11092 26792 11104
rect 26844 11092 26850 11144
rect 20671 11036 22232 11064
rect 20671 11033 20683 11036
rect 20625 11027 20683 11033
rect 22278 11024 22284 11076
rect 22336 11064 22342 11076
rect 24210 11064 24216 11076
rect 22336 11036 24216 11064
rect 22336 11024 22342 11036
rect 24210 11024 24216 11036
rect 24268 11024 24274 11076
rect 27798 11024 27804 11076
rect 27856 11024 27862 11076
rect 28552 11064 28580 11163
rect 29840 11132 29868 11296
rect 30193 11135 30251 11141
rect 30193 11132 30205 11135
rect 29840 11104 30205 11132
rect 30193 11101 30205 11104
rect 30239 11101 30251 11135
rect 30576 11132 30604 11296
rect 30834 11160 30840 11212
rect 30892 11200 30898 11212
rect 31404 11200 31432 11296
rect 32490 11228 32496 11280
rect 32548 11268 32554 11280
rect 32585 11271 32643 11277
rect 32585 11268 32597 11271
rect 32548 11240 32597 11268
rect 32548 11228 32554 11240
rect 32585 11237 32597 11240
rect 32631 11237 32643 11271
rect 32585 11231 32643 11237
rect 31481 11203 31539 11209
rect 31481 11200 31493 11203
rect 30892 11172 31248 11200
rect 31404 11172 31493 11200
rect 30892 11160 30898 11172
rect 30745 11135 30803 11141
rect 30745 11132 30757 11135
rect 30576 11104 30757 11132
rect 30193 11095 30251 11101
rect 30745 11101 30757 11104
rect 30791 11101 30803 11135
rect 30745 11095 30803 11101
rect 31021 11135 31079 11141
rect 31021 11101 31033 11135
rect 31067 11132 31079 11135
rect 31110 11132 31116 11144
rect 31067 11104 31116 11132
rect 31067 11101 31079 11104
rect 31021 11095 31079 11101
rect 31110 11092 31116 11104
rect 31168 11092 31174 11144
rect 31220 11132 31248 11172
rect 31481 11169 31493 11172
rect 31527 11169 31539 11203
rect 31481 11163 31539 11169
rect 31573 11135 31631 11141
rect 31573 11132 31585 11135
rect 31220 11104 31585 11132
rect 31573 11101 31585 11104
rect 31619 11132 31631 11135
rect 31662 11132 31668 11144
rect 31619 11104 31668 11132
rect 31619 11101 31631 11104
rect 31573 11095 31631 11101
rect 31662 11092 31668 11104
rect 31720 11092 31726 11144
rect 32600 11132 32628 11231
rect 32876 11200 32904 11296
rect 34532 11268 34560 11296
rect 34532 11240 34744 11268
rect 33045 11203 33103 11209
rect 33045 11200 33057 11203
rect 32876 11172 33057 11200
rect 33045 11169 33057 11172
rect 33091 11169 33103 11203
rect 33045 11163 33103 11169
rect 34422 11160 34428 11212
rect 34480 11200 34486 11212
rect 34517 11203 34575 11209
rect 34517 11200 34529 11203
rect 34480 11172 34529 11200
rect 34480 11160 34486 11172
rect 34517 11169 34529 11172
rect 34563 11169 34575 11203
rect 34517 11163 34575 11169
rect 34716 11141 34744 11240
rect 32769 11135 32827 11141
rect 32769 11132 32781 11135
rect 32600 11104 32781 11132
rect 32769 11101 32781 11104
rect 32815 11101 32827 11135
rect 32769 11095 32827 11101
rect 34701 11135 34759 11141
rect 34701 11101 34713 11135
rect 34747 11101 34759 11135
rect 34701 11095 34759 11101
rect 30650 11064 30656 11076
rect 28552 11036 30656 11064
rect 30650 11024 30656 11036
rect 30708 11024 30714 11076
rect 34793 11067 34851 11073
rect 34793 11064 34805 11067
rect 34270 11036 34805 11064
rect 34793 11033 34805 11036
rect 34839 11033 34851 11067
rect 34793 11027 34851 11033
rect 18003 10968 18092 10996
rect 18693 10999 18751 11005
rect 18003 10965 18015 10968
rect 17957 10959 18015 10965
rect 18693 10965 18705 10999
rect 18739 10996 18751 10999
rect 18782 10996 18788 11008
rect 18739 10968 18788 10996
rect 18739 10965 18751 10968
rect 18693 10959 18751 10965
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 20346 10956 20352 11008
rect 20404 10956 20410 11008
rect 21726 10956 21732 11008
rect 21784 10956 21790 11008
rect 28074 10956 28080 11008
rect 28132 10996 28138 11008
rect 28813 10999 28871 11005
rect 28813 10996 28825 10999
rect 28132 10968 28825 10996
rect 28132 10956 28138 10968
rect 28813 10965 28825 10968
rect 28859 10965 28871 10999
rect 28813 10959 28871 10965
rect 1104 10906 35236 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 35236 10906
rect 1104 10832 35236 10854
rect 1581 10795 1639 10801
rect 1581 10761 1593 10795
rect 1627 10792 1639 10795
rect 1670 10792 1676 10804
rect 1627 10764 1676 10792
rect 1627 10761 1639 10764
rect 1581 10755 1639 10761
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 4617 10795 4675 10801
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 5534 10792 5540 10804
rect 4663 10764 5540 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5721 10795 5779 10801
rect 5721 10761 5733 10795
rect 5767 10792 5779 10795
rect 5994 10792 6000 10804
rect 5767 10764 6000 10792
rect 5767 10761 5779 10764
rect 5721 10755 5779 10761
rect 5994 10752 6000 10764
rect 6052 10752 6058 10804
rect 6454 10752 6460 10804
rect 6512 10792 6518 10804
rect 8297 10795 8355 10801
rect 8297 10792 8309 10795
rect 6512 10764 8309 10792
rect 6512 10752 6518 10764
rect 8297 10761 8309 10764
rect 8343 10792 8355 10795
rect 8343 10764 20852 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 4154 10684 4160 10736
rect 4212 10684 4218 10736
rect 8662 10684 8668 10736
rect 8720 10684 8726 10736
rect 9030 10684 9036 10736
rect 9088 10724 9094 10736
rect 9125 10727 9183 10733
rect 9125 10724 9137 10727
rect 9088 10696 9137 10724
rect 9088 10684 9094 10696
rect 9125 10693 9137 10696
rect 9171 10693 9183 10727
rect 9125 10687 9183 10693
rect 16666 10684 16672 10736
rect 16724 10724 16730 10736
rect 17310 10724 17316 10736
rect 16724 10696 17316 10724
rect 16724 10684 16730 10696
rect 17310 10684 17316 10696
rect 17368 10724 17374 10736
rect 17586 10724 17592 10736
rect 17368 10696 17592 10724
rect 17368 10684 17374 10696
rect 17586 10684 17592 10696
rect 17644 10724 17650 10736
rect 18506 10724 18512 10736
rect 17644 10696 18512 10724
rect 17644 10684 17650 10696
rect 18506 10684 18512 10696
rect 18564 10684 18570 10736
rect 934 10616 940 10668
rect 992 10656 998 10668
rect 1397 10659 1455 10665
rect 1397 10656 1409 10659
rect 992 10628 1409 10656
rect 992 10616 998 10628
rect 1397 10625 1409 10628
rect 1443 10625 1455 10659
rect 1397 10619 1455 10625
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10625 5595 10659
rect 5537 10619 5595 10625
rect 2869 10591 2927 10597
rect 2869 10557 2881 10591
rect 2915 10557 2927 10591
rect 2869 10551 2927 10557
rect 1394 10480 1400 10532
rect 1452 10520 1458 10532
rect 2774 10520 2780 10532
rect 1452 10492 2780 10520
rect 1452 10480 1458 10492
rect 2774 10480 2780 10492
rect 2832 10520 2838 10532
rect 2884 10520 2912 10551
rect 3142 10548 3148 10600
rect 3200 10548 3206 10600
rect 3878 10548 3884 10600
rect 3936 10588 3942 10600
rect 5552 10588 5580 10619
rect 17126 10616 17132 10668
rect 17184 10656 17190 10668
rect 17494 10656 17500 10668
rect 17184 10628 17500 10656
rect 17184 10616 17190 10628
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17770 10616 17776 10668
rect 17828 10616 17834 10668
rect 17954 10616 17960 10668
rect 18012 10616 18018 10668
rect 3936 10560 5580 10588
rect 3936 10548 3942 10560
rect 2832 10492 2912 10520
rect 2832 10480 2838 10492
rect 2884 10452 2912 10492
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 12710 10520 12716 10532
rect 10744 10492 12716 10520
rect 10744 10480 10750 10492
rect 12710 10480 12716 10492
rect 12768 10520 12774 10532
rect 17770 10520 17776 10532
rect 12768 10492 17776 10520
rect 12768 10480 12774 10492
rect 17770 10480 17776 10492
rect 17828 10480 17834 10532
rect 17957 10523 18015 10529
rect 17957 10489 17969 10523
rect 18003 10520 18015 10523
rect 19242 10520 19248 10532
rect 18003 10492 19248 10520
rect 18003 10489 18015 10492
rect 17957 10483 18015 10489
rect 19242 10480 19248 10492
rect 19300 10480 19306 10532
rect 20824 10464 20852 10764
rect 20898 10752 20904 10804
rect 20956 10752 20962 10804
rect 21085 10795 21143 10801
rect 21085 10761 21097 10795
rect 21131 10792 21143 10795
rect 21919 10795 21977 10801
rect 21919 10792 21931 10795
rect 21131 10764 21931 10792
rect 21131 10761 21143 10764
rect 21085 10755 21143 10761
rect 21919 10761 21931 10764
rect 21965 10761 21977 10795
rect 21919 10755 21977 10761
rect 23477 10795 23535 10801
rect 23477 10761 23489 10795
rect 23523 10792 23535 10795
rect 24302 10792 24308 10804
rect 23523 10764 24308 10792
rect 23523 10761 23535 10764
rect 23477 10755 23535 10761
rect 24302 10752 24308 10764
rect 24360 10752 24366 10804
rect 31110 10752 31116 10804
rect 31168 10752 31174 10804
rect 31754 10792 31760 10804
rect 31496 10764 31760 10792
rect 20916 10656 20944 10752
rect 20990 10684 20996 10736
rect 21048 10684 21054 10736
rect 21266 10684 21272 10736
rect 21324 10684 21330 10736
rect 21358 10684 21364 10736
rect 21416 10724 21422 10736
rect 21821 10727 21879 10733
rect 21821 10724 21833 10727
rect 21416 10696 21833 10724
rect 21416 10684 21422 10696
rect 21821 10693 21833 10696
rect 21867 10693 21879 10727
rect 21821 10687 21879 10693
rect 22922 10684 22928 10736
rect 22980 10684 22986 10736
rect 23124 10696 23980 10724
rect 23124 10668 23152 10696
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 20916 10628 22017 10656
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 22278 10616 22284 10668
rect 22336 10616 22342 10668
rect 22554 10616 22560 10668
rect 22612 10616 22618 10668
rect 22646 10616 22652 10668
rect 22704 10656 22710 10668
rect 23106 10656 23112 10668
rect 22704 10628 23112 10656
rect 22704 10616 22710 10628
rect 23106 10616 23112 10628
rect 23164 10616 23170 10668
rect 23474 10616 23480 10668
rect 23532 10616 23538 10668
rect 23952 10665 23980 10696
rect 23937 10659 23995 10665
rect 23937 10625 23949 10659
rect 23983 10625 23995 10659
rect 23937 10619 23995 10625
rect 24210 10616 24216 10668
rect 24268 10616 24274 10668
rect 24394 10616 24400 10668
rect 24452 10616 24458 10668
rect 30650 10616 30656 10668
rect 30708 10656 30714 10668
rect 30837 10659 30895 10665
rect 30837 10656 30849 10659
rect 30708 10628 30849 10656
rect 30708 10616 30714 10628
rect 30837 10625 30849 10628
rect 30883 10625 30895 10659
rect 31128 10656 31156 10752
rect 31496 10665 31524 10764
rect 31754 10752 31760 10764
rect 31812 10752 31818 10804
rect 34514 10752 34520 10804
rect 34572 10752 34578 10804
rect 31297 10659 31355 10665
rect 31297 10656 31309 10659
rect 31128 10628 31309 10656
rect 30837 10619 30895 10625
rect 31297 10625 31309 10628
rect 31343 10625 31355 10659
rect 31297 10619 31355 10625
rect 31481 10659 31539 10665
rect 31481 10625 31493 10659
rect 31527 10625 31539 10659
rect 31481 10619 31539 10625
rect 22572 10520 22600 10616
rect 23201 10591 23259 10597
rect 23201 10557 23213 10591
rect 23247 10588 23259 10591
rect 24412 10588 24440 10616
rect 23247 10560 24440 10588
rect 30929 10591 30987 10597
rect 23247 10557 23259 10560
rect 23201 10551 23259 10557
rect 30929 10557 30941 10591
rect 30975 10588 30987 10591
rect 31389 10591 31447 10597
rect 31389 10588 31401 10591
rect 30975 10560 31401 10588
rect 30975 10557 30987 10560
rect 30929 10551 30987 10557
rect 31389 10557 31401 10560
rect 31435 10557 31447 10591
rect 31389 10551 31447 10557
rect 21560 10492 22600 10520
rect 31205 10523 31263 10529
rect 4893 10455 4951 10461
rect 4893 10452 4905 10455
rect 2884 10424 4905 10452
rect 4893 10421 4905 10424
rect 4939 10421 4951 10455
rect 4893 10415 4951 10421
rect 20806 10412 20812 10464
rect 20864 10412 20870 10464
rect 21560 10461 21588 10492
rect 31205 10489 31217 10523
rect 31251 10520 31263 10523
rect 32398 10520 32404 10532
rect 31251 10492 32404 10520
rect 31251 10489 31263 10492
rect 31205 10483 31263 10489
rect 32398 10480 32404 10492
rect 32456 10480 32462 10532
rect 21545 10455 21603 10461
rect 21545 10421 21557 10455
rect 21591 10421 21603 10455
rect 21545 10415 21603 10421
rect 1104 10362 35248 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 35248 10362
rect 1104 10288 35248 10310
rect 2774 10208 2780 10260
rect 2832 10208 2838 10260
rect 3145 10251 3203 10257
rect 3145 10217 3157 10251
rect 3191 10248 3203 10251
rect 3878 10248 3884 10260
rect 3191 10220 3884 10248
rect 3191 10217 3203 10220
rect 3145 10211 3203 10217
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 16025 10251 16083 10257
rect 16025 10217 16037 10251
rect 16071 10248 16083 10251
rect 16071 10220 17172 10248
rect 16071 10217 16083 10220
rect 16025 10211 16083 10217
rect 2792 10180 2820 10208
rect 3513 10183 3571 10189
rect 3513 10180 3525 10183
rect 2792 10152 3525 10180
rect 3513 10149 3525 10152
rect 3559 10149 3571 10183
rect 17037 10183 17095 10189
rect 17037 10180 17049 10183
rect 3513 10143 3571 10149
rect 16408 10152 17049 10180
rect 1394 10072 1400 10124
rect 1452 10072 1458 10124
rect 16117 10115 16175 10121
rect 16117 10081 16129 10115
rect 16163 10112 16175 10115
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 16163 10084 16313 10112
rect 16163 10081 16175 10084
rect 16117 10075 16175 10081
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 16301 10075 16359 10081
rect 2774 10004 2780 10056
rect 2832 10004 2838 10056
rect 15654 10004 15660 10056
rect 15712 10004 15718 10056
rect 16209 10047 16267 10053
rect 16209 10013 16221 10047
rect 16255 10044 16267 10047
rect 16408 10044 16436 10152
rect 17037 10149 17049 10152
rect 17083 10149 17095 10183
rect 17144 10180 17172 10220
rect 17218 10208 17224 10260
rect 17276 10208 17282 10260
rect 17494 10208 17500 10260
rect 17552 10248 17558 10260
rect 18322 10248 18328 10260
rect 17552 10220 18328 10248
rect 17552 10208 17558 10220
rect 18322 10208 18328 10220
rect 18380 10208 18386 10260
rect 22094 10248 22100 10260
rect 20732 10220 22100 10248
rect 20732 10189 20760 10220
rect 22094 10208 22100 10220
rect 22152 10208 22158 10260
rect 22281 10251 22339 10257
rect 22281 10217 22293 10251
rect 22327 10248 22339 10251
rect 23474 10248 23480 10260
rect 22327 10220 23480 10248
rect 22327 10217 22339 10220
rect 22281 10211 22339 10217
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 20717 10183 20775 10189
rect 17144 10152 18184 10180
rect 17037 10143 17095 10149
rect 17218 10112 17224 10124
rect 16776 10084 17224 10112
rect 16255 10016 16436 10044
rect 16255 10013 16267 10016
rect 16209 10007 16267 10013
rect 16482 10004 16488 10056
rect 16540 10004 16546 10056
rect 16574 10004 16580 10056
rect 16632 10004 16638 10056
rect 16666 10004 16672 10056
rect 16724 10004 16730 10056
rect 16776 10053 16804 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10013 16819 10047
rect 16761 10007 16819 10013
rect 16945 10047 17003 10053
rect 16945 10013 16957 10047
rect 16991 10013 17003 10047
rect 16945 10007 17003 10013
rect 1670 9936 1676 9988
rect 1728 9936 1734 9988
rect 15749 9911 15807 9917
rect 15749 9877 15761 9911
rect 15795 9908 15807 9911
rect 16500 9908 16528 10004
rect 15795 9880 16528 9908
rect 16960 9908 16988 10007
rect 17034 10004 17040 10056
rect 17092 10004 17098 10056
rect 17494 10044 17500 10056
rect 17420 10016 17500 10044
rect 17052 9976 17080 10004
rect 17420 9985 17448 10016
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 17678 10044 17684 10056
rect 17635 10016 17684 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17205 9979 17263 9985
rect 17205 9976 17217 9979
rect 17052 9948 17217 9976
rect 17205 9945 17217 9948
rect 17251 9945 17263 9979
rect 17205 9939 17263 9945
rect 17405 9979 17463 9985
rect 17405 9945 17417 9979
rect 17451 9945 17463 9979
rect 17405 9939 17463 9945
rect 17604 9908 17632 10007
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10044 17831 10047
rect 17862 10044 17868 10056
rect 17819 10016 17868 10044
rect 17819 10013 17831 10016
rect 17773 10007 17831 10013
rect 17862 10004 17868 10016
rect 17920 10004 17926 10056
rect 18156 10053 18184 10152
rect 20717 10149 20729 10183
rect 20763 10149 20775 10183
rect 20717 10143 20775 10149
rect 20806 10140 20812 10192
rect 20864 10180 20870 10192
rect 31481 10183 31539 10189
rect 20864 10152 22094 10180
rect 20864 10140 20870 10152
rect 20438 10072 20444 10124
rect 20496 10072 20502 10124
rect 20990 10072 20996 10124
rect 21048 10112 21054 10124
rect 21637 10115 21695 10121
rect 21637 10112 21649 10115
rect 21048 10084 21649 10112
rect 21048 10072 21054 10084
rect 21637 10081 21649 10084
rect 21683 10081 21695 10115
rect 21637 10075 21695 10081
rect 21726 10072 21732 10124
rect 21784 10112 21790 10124
rect 21821 10115 21879 10121
rect 21821 10112 21833 10115
rect 21784 10084 21833 10112
rect 21784 10072 21790 10084
rect 21821 10081 21833 10084
rect 21867 10081 21879 10115
rect 22066 10112 22094 10152
rect 31481 10149 31493 10183
rect 31527 10180 31539 10183
rect 31527 10152 31754 10180
rect 31527 10149 31539 10152
rect 31481 10143 31539 10149
rect 22066 10084 26096 10112
rect 21821 10075 21879 10081
rect 18141 10047 18199 10053
rect 18141 10013 18153 10047
rect 18187 10013 18199 10047
rect 18141 10007 18199 10013
rect 18322 10004 18328 10056
rect 18380 10004 18386 10056
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 18543 10047 18601 10053
rect 18543 10013 18555 10047
rect 18589 10044 18601 10047
rect 19978 10044 19984 10056
rect 18589 10016 19984 10044
rect 18589 10013 18601 10016
rect 18543 10007 18601 10013
rect 19978 10004 19984 10016
rect 20036 10004 20042 10056
rect 20346 10004 20352 10056
rect 20404 10004 20410 10056
rect 21266 10004 21272 10056
rect 21324 10044 21330 10056
rect 21913 10047 21971 10053
rect 21913 10044 21925 10047
rect 21324 10016 21925 10044
rect 21324 10004 21330 10016
rect 21913 10013 21925 10016
rect 21959 10013 21971 10047
rect 22646 10044 22652 10056
rect 21913 10007 21971 10013
rect 22066 10016 22652 10044
rect 18785 9979 18843 9985
rect 18785 9945 18797 9979
rect 18831 9976 18843 9979
rect 22066 9976 22094 10016
rect 22646 10004 22652 10016
rect 22704 10004 22710 10056
rect 26068 10053 26096 10084
rect 26053 10047 26111 10053
rect 26053 10013 26065 10047
rect 26099 10044 26111 10047
rect 27522 10044 27528 10056
rect 26099 10016 27528 10044
rect 26099 10013 26111 10016
rect 26053 10007 26111 10013
rect 27522 10004 27528 10016
rect 27580 10044 27586 10056
rect 28074 10044 28080 10056
rect 27580 10016 28080 10044
rect 27580 10004 27586 10016
rect 28074 10004 28080 10016
rect 28132 10004 28138 10056
rect 31110 10004 31116 10056
rect 31168 10044 31174 10056
rect 31297 10047 31355 10053
rect 31297 10044 31309 10047
rect 31168 10016 31309 10044
rect 31168 10004 31174 10016
rect 31297 10013 31309 10016
rect 31343 10013 31355 10047
rect 31726 10044 31754 10152
rect 34057 10115 34115 10121
rect 34057 10081 34069 10115
rect 34103 10081 34115 10115
rect 34057 10075 34115 10081
rect 32033 10047 32091 10053
rect 32033 10044 32045 10047
rect 31726 10016 32045 10044
rect 31297 10007 31355 10013
rect 32033 10013 32045 10016
rect 32079 10013 32091 10047
rect 32033 10007 32091 10013
rect 32677 10047 32735 10053
rect 32677 10013 32689 10047
rect 32723 10044 32735 10047
rect 32723 10016 32757 10044
rect 32723 10013 32735 10016
rect 32677 10007 32735 10013
rect 32585 9979 32643 9985
rect 32585 9976 32597 9979
rect 18831 9948 22094 9976
rect 22204 9948 26004 9976
rect 18831 9945 18843 9948
rect 18785 9939 18843 9945
rect 16960 9880 17632 9908
rect 15795 9877 15807 9880
rect 15749 9871 15807 9877
rect 17678 9868 17684 9920
rect 17736 9868 17742 9920
rect 17770 9868 17776 9920
rect 17828 9908 17834 9920
rect 22204 9908 22232 9948
rect 17828 9880 22232 9908
rect 25976 9908 26004 9948
rect 27356 9948 32597 9976
rect 27356 9917 27384 9948
rect 32585 9945 32597 9948
rect 32631 9976 32643 9979
rect 32692 9976 32720 10007
rect 34072 9988 34100 10075
rect 34422 10004 34428 10056
rect 34480 10004 34486 10056
rect 32631 9948 33272 9976
rect 32631 9945 32643 9948
rect 32585 9939 32643 9945
rect 27341 9911 27399 9917
rect 27341 9908 27353 9911
rect 25976 9880 27353 9908
rect 17828 9868 17834 9880
rect 27341 9877 27353 9880
rect 27387 9877 27399 9911
rect 27341 9871 27399 9877
rect 32217 9911 32275 9917
rect 32217 9877 32229 9911
rect 32263 9908 32275 9911
rect 32306 9908 32312 9920
rect 32263 9880 32312 9908
rect 32263 9877 32275 9880
rect 32217 9871 32275 9877
rect 32306 9868 32312 9880
rect 32364 9868 32370 9920
rect 32769 9911 32827 9917
rect 32769 9877 32781 9911
rect 32815 9908 32827 9911
rect 33134 9908 33140 9920
rect 32815 9880 33140 9908
rect 32815 9877 32827 9880
rect 32769 9871 32827 9877
rect 33134 9868 33140 9880
rect 33192 9868 33198 9920
rect 33244 9908 33272 9948
rect 34054 9936 34060 9988
rect 34112 9936 34118 9988
rect 34146 9908 34152 9920
rect 33244 9880 34152 9908
rect 34146 9868 34152 9880
rect 34204 9868 34210 9920
rect 1104 9818 35236 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 35236 9818
rect 1104 9744 35236 9766
rect 2774 9664 2780 9716
rect 2832 9664 2838 9716
rect 17497 9707 17555 9713
rect 17497 9673 17509 9707
rect 17543 9673 17555 9707
rect 17497 9667 17555 9673
rect 18141 9707 18199 9713
rect 18141 9673 18153 9707
rect 18187 9704 18199 9707
rect 18414 9704 18420 9716
rect 18187 9676 18420 9704
rect 18187 9673 18199 9676
rect 18141 9667 18199 9673
rect 2409 9639 2467 9645
rect 2409 9605 2421 9639
rect 2455 9636 2467 9639
rect 2792 9636 2820 9664
rect 2455 9608 2820 9636
rect 2455 9605 2467 9608
rect 2409 9599 2467 9605
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 16853 9639 16911 9645
rect 16853 9636 16865 9639
rect 16724 9608 16865 9636
rect 16724 9596 16730 9608
rect 16853 9605 16865 9608
rect 16899 9605 16911 9639
rect 17512 9636 17540 9667
rect 18414 9664 18420 9676
rect 18472 9664 18478 9716
rect 18322 9636 18328 9648
rect 17512 9608 18328 9636
rect 16853 9599 16911 9605
rect 18322 9596 18328 9608
rect 18380 9596 18386 9648
rect 20990 9636 20996 9648
rect 18524 9608 19472 9636
rect 20378 9608 20996 9636
rect 2317 9571 2375 9577
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2682 9568 2688 9580
rect 2363 9540 2688 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2682 9528 2688 9540
rect 2740 9568 2746 9580
rect 2777 9571 2835 9577
rect 2777 9568 2789 9571
rect 2740 9540 2789 9568
rect 2740 9528 2746 9540
rect 2777 9537 2789 9540
rect 2823 9537 2835 9571
rect 2777 9531 2835 9537
rect 16482 9528 16488 9580
rect 16540 9528 16546 9580
rect 17218 9528 17224 9580
rect 17276 9528 17282 9580
rect 17862 9577 17868 9580
rect 17313 9571 17371 9577
rect 17313 9537 17325 9571
rect 17359 9568 17371 9571
rect 17851 9571 17868 9577
rect 17359 9540 17816 9568
rect 17359 9537 17371 9540
rect 17313 9531 17371 9537
rect 15654 9460 15660 9512
rect 15712 9460 15718 9512
rect 16500 9500 16528 9528
rect 17328 9500 17356 9531
rect 16500 9472 17356 9500
rect 17678 9460 17684 9512
rect 17736 9460 17742 9512
rect 17788 9500 17816 9540
rect 17851 9537 17863 9571
rect 17920 9568 17926 9580
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 17920 9540 18429 9568
rect 17851 9531 17868 9537
rect 17862 9528 17868 9531
rect 17920 9528 17926 9540
rect 18417 9537 18429 9540
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 17788 9472 17908 9500
rect 15672 9432 15700 9460
rect 17880 9432 17908 9472
rect 18138 9460 18144 9512
rect 18196 9500 18202 9512
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 18196 9472 18245 9500
rect 18196 9460 18202 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 18524 9432 18552 9608
rect 18708 9577 18736 9608
rect 19444 9580 19472 9608
rect 20990 9596 20996 9608
rect 21048 9596 21054 9648
rect 32398 9596 32404 9648
rect 32456 9596 32462 9648
rect 33134 9596 33140 9648
rect 33192 9596 33198 9648
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18693 9571 18751 9577
rect 18693 9537 18705 9571
rect 18739 9537 18751 9571
rect 18877 9571 18935 9577
rect 18877 9568 18889 9571
rect 18693 9531 18751 9537
rect 18800 9540 18889 9568
rect 15672 9404 17816 9432
rect 17880 9404 18552 9432
rect 18616 9500 18644 9531
rect 18800 9500 18828 9540
rect 18877 9537 18889 9540
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 19426 9528 19432 9580
rect 19484 9528 19490 9580
rect 27157 9571 27215 9577
rect 27157 9537 27169 9571
rect 27203 9568 27215 9571
rect 27338 9568 27344 9580
rect 27203 9540 27344 9568
rect 27203 9537 27215 9540
rect 27157 9531 27215 9537
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 27522 9528 27528 9580
rect 27580 9528 27586 9580
rect 34146 9528 34152 9580
rect 34204 9568 34210 9580
rect 34425 9571 34483 9577
rect 34425 9568 34437 9571
rect 34204 9540 34437 9568
rect 34204 9528 34210 9540
rect 34425 9537 34437 9540
rect 34471 9537 34483 9571
rect 34425 9531 34483 9537
rect 18616 9472 18828 9500
rect 27433 9503 27491 9509
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 16945 9367 17003 9373
rect 16945 9364 16957 9367
rect 16632 9336 16957 9364
rect 16632 9324 16638 9336
rect 16945 9333 16957 9336
rect 16991 9333 17003 9367
rect 17788 9364 17816 9404
rect 18616 9376 18644 9472
rect 27433 9469 27445 9503
rect 27479 9500 27491 9503
rect 27540 9500 27568 9528
rect 27479 9472 27568 9500
rect 31941 9503 31999 9509
rect 27479 9469 27491 9472
rect 27433 9463 27491 9469
rect 31941 9469 31953 9503
rect 31987 9500 31999 9503
rect 32030 9500 32036 9512
rect 31987 9472 32036 9500
rect 31987 9469 31999 9472
rect 31941 9463 31999 9469
rect 32030 9460 32036 9472
rect 32088 9500 32094 9512
rect 32125 9503 32183 9509
rect 32125 9500 32137 9503
rect 32088 9472 32137 9500
rect 32088 9460 32094 9472
rect 32125 9469 32137 9472
rect 32171 9500 32183 9503
rect 32490 9500 32496 9512
rect 32171 9472 32496 9500
rect 32171 9469 32183 9472
rect 32125 9463 32183 9469
rect 32490 9460 32496 9472
rect 32548 9460 32554 9512
rect 18598 9364 18604 9376
rect 17788 9336 18604 9364
rect 16945 9327 17003 9333
rect 18598 9324 18604 9336
rect 18656 9324 18662 9376
rect 33870 9324 33876 9376
rect 33928 9324 33934 9376
rect 34054 9324 34060 9376
rect 34112 9324 34118 9376
rect 1104 9274 35248 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 35248 9274
rect 1104 9200 35248 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 2866 9160 2872 9172
rect 1627 9132 2872 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 16666 9120 16672 9172
rect 16724 9120 16730 9172
rect 17681 9163 17739 9169
rect 17681 9129 17693 9163
rect 17727 9160 17739 9163
rect 17862 9160 17868 9172
rect 17727 9132 17868 9160
rect 17727 9129 17739 9132
rect 17681 9123 17739 9129
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18598 9120 18604 9172
rect 18656 9120 18662 9172
rect 19521 9163 19579 9169
rect 19521 9129 19533 9163
rect 19567 9160 19579 9163
rect 19978 9160 19984 9172
rect 19567 9132 19984 9160
rect 19567 9129 19579 9132
rect 19521 9123 19579 9129
rect 19978 9120 19984 9132
rect 20036 9120 20042 9172
rect 32030 9120 32036 9172
rect 32088 9120 32094 9172
rect 16684 9024 16712 9120
rect 16684 8996 17724 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 17696 8965 17724 8996
rect 17497 8959 17555 8965
rect 17497 8956 17509 8959
rect 16632 8928 17509 8956
rect 16632 8916 16638 8928
rect 17497 8925 17509 8928
rect 17543 8925 17555 8959
rect 17497 8919 17555 8925
rect 17681 8959 17739 8965
rect 17681 8925 17693 8959
rect 17727 8925 17739 8959
rect 18616 8956 18644 9120
rect 19426 9052 19432 9104
rect 19484 9052 19490 9104
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 18616 8928 19349 8956
rect 17681 8919 17739 8925
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19444 8956 19472 9052
rect 32048 9024 32076 9120
rect 32125 9027 32183 9033
rect 32125 9024 32137 9027
rect 32048 8996 32137 9024
rect 32125 8993 32137 8996
rect 32171 8993 32183 9027
rect 32125 8987 32183 8993
rect 19521 8959 19579 8965
rect 19521 8956 19533 8959
rect 19444 8928 19533 8956
rect 19337 8919 19395 8925
rect 19521 8925 19533 8928
rect 19567 8925 19579 8959
rect 34054 8956 34060 8968
rect 33534 8928 34060 8956
rect 19521 8919 19579 8925
rect 34054 8916 34060 8928
rect 34112 8916 34118 8968
rect 32306 8848 32312 8900
rect 32364 8888 32370 8900
rect 32401 8891 32459 8897
rect 32401 8888 32413 8891
rect 32364 8860 32413 8888
rect 32364 8848 32370 8860
rect 32401 8857 32413 8860
rect 32447 8857 32459 8891
rect 32401 8851 32459 8857
rect 33318 8780 33324 8832
rect 33376 8820 33382 8832
rect 33873 8823 33931 8829
rect 33873 8820 33885 8823
rect 33376 8792 33885 8820
rect 33376 8780 33382 8792
rect 33873 8789 33885 8792
rect 33919 8789 33931 8823
rect 33873 8783 33931 8789
rect 1104 8730 35236 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 35236 8730
rect 1104 8656 35236 8678
rect 1104 8186 35248 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 35248 8186
rect 1104 8112 35248 8134
rect 34057 7939 34115 7945
rect 34057 7905 34069 7939
rect 34103 7936 34115 7939
rect 34103 7908 34652 7936
rect 34103 7905 34115 7908
rect 34057 7899 34115 7905
rect 34238 7828 34244 7880
rect 34296 7868 34302 7880
rect 34333 7871 34391 7877
rect 34333 7868 34345 7871
rect 34296 7840 34345 7868
rect 34296 7828 34302 7840
rect 34333 7837 34345 7840
rect 34379 7837 34391 7871
rect 34333 7831 34391 7837
rect 34624 7812 34652 7908
rect 34606 7760 34612 7812
rect 34664 7760 34670 7812
rect 1104 7642 35236 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 35236 7642
rect 1104 7568 35236 7590
rect 1104 7098 35248 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 35248 7098
rect 1104 7024 35248 7046
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 992 6752 1409 6780
rect 992 6740 998 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1578 6604 1584 6656
rect 1636 6604 1642 6656
rect 1104 6554 35236 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 35236 6554
rect 1104 6480 35236 6502
rect 1104 6010 35248 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 35248 6010
rect 1104 5936 35248 5958
rect 33321 5695 33379 5701
rect 33321 5661 33333 5695
rect 33367 5692 33379 5695
rect 33870 5692 33876 5704
rect 33367 5664 33876 5692
rect 33367 5661 33379 5664
rect 33321 5655 33379 5661
rect 33870 5652 33876 5664
rect 33928 5652 33934 5704
rect 34330 5584 34336 5636
rect 34388 5584 34394 5636
rect 1104 5466 35236 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 35236 5466
rect 1104 5392 35236 5414
rect 1104 4922 35248 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 35248 4922
rect 1104 4848 35248 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 2958 4808 2964 4820
rect 1627 4780 2964 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1104 4378 35236 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 35236 4378
rect 1104 4304 35236 4326
rect 1104 3834 35248 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 35248 3834
rect 1104 3760 35248 3782
rect 33318 3476 33324 3528
rect 33376 3476 33382 3528
rect 34333 3451 34391 3457
rect 34333 3417 34345 3451
rect 34379 3448 34391 3451
rect 34882 3448 34888 3460
rect 34379 3420 34888 3448
rect 34379 3417 34391 3420
rect 34333 3411 34391 3417
rect 34882 3408 34888 3420
rect 34940 3408 34946 3460
rect 1104 3290 35236 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 35236 3290
rect 1104 3216 35236 3238
rect 1104 2746 35248 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 35248 2746
rect 1104 2672 35248 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 1581 2635 1639 2641
rect 1581 2632 1593 2635
rect 1544 2604 1593 2632
rect 1544 2592 1550 2604
rect 1581 2601 1593 2604
rect 1627 2601 1639 2635
rect 1581 2595 1639 2601
rect 27338 2592 27344 2644
rect 27396 2592 27402 2644
rect 9030 2456 9036 2508
rect 9088 2496 9094 2508
rect 9585 2499 9643 2505
rect 9585 2496 9597 2499
rect 9088 2468 9597 2496
rect 9088 2456 9094 2468
rect 9585 2465 9597 2468
rect 9631 2465 9643 2499
rect 9585 2459 9643 2465
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 27246 2388 27252 2440
rect 27304 2428 27310 2440
rect 27525 2431 27583 2437
rect 27525 2428 27537 2431
rect 27304 2400 27537 2428
rect 27304 2388 27310 2400
rect 27525 2397 27537 2400
rect 27571 2397 27583 2431
rect 27525 2391 27583 2397
rect 1104 2202 35236 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 35236 2202
rect 1104 2128 35236 2150
<< via1 >>
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 940 36116 992 36168
rect 33876 36116 33928 36168
rect 34336 36091 34388 36100
rect 34336 36057 34345 36091
rect 34345 36057 34379 36091
rect 34379 36057 34388 36091
rect 34336 36048 34388 36057
rect 1584 36023 1636 36032
rect 1584 35989 1593 36023
rect 1593 35989 1627 36023
rect 1627 35989 1636 36023
rect 1584 35980 1636 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 940 35028 992 35080
rect 2872 34892 2924 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 34612 33872 34664 33924
rect 34704 33804 34756 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 940 32852 992 32904
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 34520 31807 34572 31816
rect 34520 31773 34529 31807
rect 34529 31773 34563 31807
rect 34563 31773 34572 31807
rect 34520 31764 34572 31773
rect 34060 31628 34112 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 3700 30540 3752 30592
rect 33140 30540 33192 30592
rect 34428 30540 34480 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 29276 30268 29328 30320
rect 33140 30268 33192 30320
rect 28816 30175 28868 30184
rect 28816 30141 28825 30175
rect 28825 30141 28859 30175
rect 28859 30141 28868 30175
rect 28816 30132 28868 30141
rect 31852 30200 31904 30252
rect 31024 30175 31076 30184
rect 31024 30141 31033 30175
rect 31033 30141 31067 30175
rect 31067 30141 31076 30175
rect 31024 30132 31076 30141
rect 33876 30107 33928 30116
rect 33876 30073 33885 30107
rect 33885 30073 33919 30107
rect 33919 30073 33928 30107
rect 33876 30064 33928 30073
rect 29828 29996 29880 30048
rect 31852 30039 31904 30048
rect 31852 30005 31861 30039
rect 31861 30005 31895 30039
rect 31895 30005 31904 30039
rect 31852 29996 31904 30005
rect 34244 30039 34296 30048
rect 34244 30005 34253 30039
rect 34253 30005 34287 30039
rect 34287 30005 34296 30039
rect 34244 29996 34296 30005
rect 34428 29996 34480 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 28816 29792 28868 29844
rect 29276 29835 29328 29844
rect 29276 29801 29285 29835
rect 29285 29801 29319 29835
rect 29319 29801 29328 29835
rect 29276 29792 29328 29801
rect 34520 29835 34572 29844
rect 34520 29801 34529 29835
rect 34529 29801 34563 29835
rect 34563 29801 34572 29835
rect 34520 29792 34572 29801
rect 25136 29699 25188 29708
rect 25136 29665 25145 29699
rect 25145 29665 25179 29699
rect 25179 29665 25188 29699
rect 25136 29656 25188 29665
rect 29828 29656 29880 29708
rect 32220 29699 32272 29708
rect 32220 29665 32229 29699
rect 32229 29665 32263 29699
rect 32263 29665 32272 29699
rect 32220 29656 32272 29665
rect 24860 29588 24912 29640
rect 24676 29520 24728 29572
rect 26976 29588 27028 29640
rect 28356 29588 28408 29640
rect 29184 29631 29236 29640
rect 29184 29597 29193 29631
rect 29193 29597 29227 29631
rect 29227 29597 29236 29631
rect 29184 29588 29236 29597
rect 31668 29588 31720 29640
rect 27068 29520 27120 29572
rect 23388 29452 23440 29504
rect 24308 29452 24360 29504
rect 24400 29452 24452 29504
rect 30380 29520 30432 29572
rect 31852 29520 31904 29572
rect 32588 29588 32640 29640
rect 34244 29724 34296 29776
rect 29184 29452 29236 29504
rect 30196 29452 30248 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 23664 29248 23716 29300
rect 23940 29223 23992 29232
rect 23940 29189 23949 29223
rect 23949 29189 23983 29223
rect 23983 29189 23992 29223
rect 23940 29180 23992 29189
rect 23572 29155 23624 29164
rect 23572 29121 23581 29155
rect 23581 29121 23615 29155
rect 23615 29121 23624 29155
rect 23572 29112 23624 29121
rect 24860 29248 24912 29300
rect 25136 29291 25188 29300
rect 25136 29257 25145 29291
rect 25145 29257 25179 29291
rect 25179 29257 25188 29291
rect 25136 29248 25188 29257
rect 29828 29248 29880 29300
rect 30380 29291 30432 29300
rect 30380 29257 30389 29291
rect 30389 29257 30423 29291
rect 30423 29257 30432 29291
rect 30380 29248 30432 29257
rect 32588 29291 32640 29300
rect 32588 29257 32597 29291
rect 32597 29257 32631 29291
rect 32631 29257 32640 29291
rect 32588 29248 32640 29257
rect 24308 29180 24360 29232
rect 24400 29155 24452 29164
rect 24400 29121 24409 29155
rect 24409 29121 24443 29155
rect 24443 29121 24452 29155
rect 24400 29112 24452 29121
rect 24860 29155 24912 29164
rect 24860 29121 24869 29155
rect 24869 29121 24903 29155
rect 24903 29121 24912 29155
rect 24860 29112 24912 29121
rect 25044 29112 25096 29164
rect 25136 29155 25188 29164
rect 25136 29121 25145 29155
rect 25145 29121 25179 29155
rect 25179 29121 25188 29155
rect 25136 29112 25188 29121
rect 26976 28976 27028 29028
rect 34704 29248 34756 29300
rect 34796 29180 34848 29232
rect 23480 28951 23532 28960
rect 23480 28917 23489 28951
rect 23489 28917 23523 28951
rect 23523 28917 23532 28951
rect 23480 28908 23532 28917
rect 26240 28908 26292 28960
rect 27988 28908 28040 28960
rect 28540 28908 28592 28960
rect 30196 28951 30248 28960
rect 30196 28917 30205 28951
rect 30205 28917 30239 28951
rect 30239 28917 30248 28951
rect 30196 28908 30248 28917
rect 33048 28908 33100 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 23940 28704 23992 28756
rect 28356 28747 28408 28756
rect 24768 28679 24820 28688
rect 24768 28645 24777 28679
rect 24777 28645 24811 28679
rect 24811 28645 24820 28679
rect 24768 28636 24820 28645
rect 26516 28636 26568 28688
rect 940 28500 992 28552
rect 23480 28500 23532 28552
rect 24492 28568 24544 28620
rect 25136 28568 25188 28620
rect 28356 28713 28365 28747
rect 28365 28713 28399 28747
rect 28399 28713 28408 28747
rect 28356 28704 28408 28713
rect 31024 28704 31076 28756
rect 33048 28704 33100 28756
rect 34796 28747 34848 28756
rect 34796 28713 34805 28747
rect 34805 28713 34839 28747
rect 34839 28713 34848 28747
rect 34796 28704 34848 28713
rect 28264 28636 28316 28688
rect 26976 28611 27028 28620
rect 26976 28577 26985 28611
rect 26985 28577 27019 28611
rect 27019 28577 27028 28611
rect 26976 28568 27028 28577
rect 28080 28568 28132 28620
rect 23664 28432 23716 28484
rect 26240 28500 26292 28552
rect 26332 28500 26384 28552
rect 27068 28500 27120 28552
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 23572 28407 23624 28416
rect 23572 28373 23581 28407
rect 23581 28373 23615 28407
rect 23615 28373 23624 28407
rect 23572 28364 23624 28373
rect 25044 28432 25096 28484
rect 25412 28432 25464 28484
rect 27988 28543 28040 28552
rect 27988 28509 27997 28543
rect 27997 28509 28031 28543
rect 28031 28509 28040 28543
rect 27988 28500 28040 28509
rect 28172 28543 28224 28552
rect 28172 28509 28181 28543
rect 28181 28509 28215 28543
rect 28215 28509 28224 28543
rect 28172 28500 28224 28509
rect 28080 28432 28132 28484
rect 24860 28364 24912 28416
rect 26240 28364 26292 28416
rect 27712 28364 27764 28416
rect 28540 28475 28592 28484
rect 28540 28441 28549 28475
rect 28549 28441 28583 28475
rect 28583 28441 28592 28475
rect 28540 28432 28592 28441
rect 31668 28679 31720 28688
rect 31668 28645 31677 28679
rect 31677 28645 31711 28679
rect 31711 28645 31720 28679
rect 31668 28636 31720 28645
rect 32220 28636 32272 28688
rect 29828 28568 29880 28620
rect 32312 28611 32364 28620
rect 32312 28577 32321 28611
rect 32321 28577 32355 28611
rect 32355 28577 32364 28611
rect 32312 28568 32364 28577
rect 34060 28611 34112 28620
rect 34060 28577 34069 28611
rect 34069 28577 34103 28611
rect 34103 28577 34112 28611
rect 34060 28568 34112 28577
rect 30288 28432 30340 28484
rect 31760 28543 31812 28552
rect 31760 28509 31769 28543
rect 31769 28509 31803 28543
rect 31803 28509 31812 28543
rect 31760 28500 31812 28509
rect 32036 28500 32088 28552
rect 31760 28364 31812 28416
rect 34520 28543 34572 28552
rect 34520 28509 34529 28543
rect 34529 28509 34563 28543
rect 34563 28509 34572 28543
rect 34520 28500 34572 28509
rect 32772 28364 32824 28416
rect 34428 28364 34480 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 27712 28203 27764 28212
rect 27712 28169 27721 28203
rect 27721 28169 27755 28203
rect 27755 28169 27764 28203
rect 27712 28160 27764 28169
rect 28080 28160 28132 28212
rect 30288 28203 30340 28212
rect 30288 28169 30297 28203
rect 30297 28169 30331 28203
rect 30331 28169 30340 28203
rect 30288 28160 30340 28169
rect 32312 28160 32364 28212
rect 27528 28067 27580 28076
rect 27528 28033 27537 28067
rect 27537 28033 27571 28067
rect 27571 28033 27580 28067
rect 27528 28024 27580 28033
rect 27712 28067 27764 28076
rect 27712 28033 27721 28067
rect 27721 28033 27755 28067
rect 27755 28033 27764 28067
rect 27712 28024 27764 28033
rect 30196 28067 30248 28076
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 31668 28024 31720 28076
rect 23572 27956 23624 28008
rect 28172 27956 28224 28008
rect 32036 27956 32088 28008
rect 32772 27956 32824 28008
rect 31300 27820 31352 27872
rect 31760 27820 31812 27872
rect 32312 27820 32364 27872
rect 34428 27820 34480 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 21364 27616 21416 27668
rect 24400 27616 24452 27668
rect 24768 27659 24820 27668
rect 24768 27625 24777 27659
rect 24777 27625 24811 27659
rect 24811 27625 24820 27659
rect 24768 27616 24820 27625
rect 26240 27659 26292 27668
rect 26240 27625 26249 27659
rect 26249 27625 26283 27659
rect 26283 27625 26292 27659
rect 26240 27616 26292 27625
rect 26332 27659 26384 27668
rect 26332 27625 26341 27659
rect 26341 27625 26375 27659
rect 26375 27625 26384 27659
rect 26332 27616 26384 27625
rect 31760 27659 31812 27668
rect 31760 27625 31769 27659
rect 31769 27625 31803 27659
rect 31803 27625 31812 27659
rect 31760 27616 31812 27625
rect 34520 27659 34572 27668
rect 34520 27625 34529 27659
rect 34529 27625 34563 27659
rect 34563 27625 34572 27659
rect 34520 27616 34572 27625
rect 23388 27548 23440 27600
rect 22468 27480 22520 27532
rect 19248 27455 19300 27464
rect 19248 27421 19257 27455
rect 19257 27421 19291 27455
rect 19291 27421 19300 27455
rect 19248 27412 19300 27421
rect 19340 27455 19392 27464
rect 19340 27421 19349 27455
rect 19349 27421 19383 27455
rect 19383 27421 19392 27455
rect 19340 27412 19392 27421
rect 19432 27412 19484 27464
rect 18972 27344 19024 27396
rect 19984 27455 20036 27464
rect 19984 27421 19993 27455
rect 19993 27421 20027 27455
rect 20027 27421 20036 27455
rect 19984 27412 20036 27421
rect 20076 27455 20128 27464
rect 20076 27421 20085 27455
rect 20085 27421 20119 27455
rect 20119 27421 20128 27455
rect 20076 27412 20128 27421
rect 17592 27276 17644 27328
rect 20260 27276 20312 27328
rect 20444 27319 20496 27328
rect 20444 27285 20453 27319
rect 20453 27285 20487 27319
rect 20487 27285 20496 27319
rect 20444 27276 20496 27285
rect 22192 27276 22244 27328
rect 23204 27276 23256 27328
rect 24492 27412 24544 27464
rect 27712 27480 27764 27532
rect 25412 27412 25464 27464
rect 25964 27455 26016 27464
rect 25964 27421 25973 27455
rect 25973 27421 26007 27455
rect 26007 27421 26016 27455
rect 25964 27412 26016 27421
rect 26148 27412 26200 27464
rect 26332 27387 26384 27396
rect 26332 27353 26341 27387
rect 26341 27353 26375 27387
rect 26375 27353 26384 27387
rect 26332 27344 26384 27353
rect 26424 27344 26476 27396
rect 27528 27344 27580 27396
rect 28540 27412 28592 27464
rect 31668 27480 31720 27532
rect 32128 27523 32180 27532
rect 32128 27489 32137 27523
rect 32137 27489 32171 27523
rect 32171 27489 32180 27523
rect 32128 27480 32180 27489
rect 32588 27480 32640 27532
rect 34520 27412 34572 27464
rect 25044 27276 25096 27328
rect 25872 27276 25924 27328
rect 29092 27319 29144 27328
rect 29092 27285 29101 27319
rect 29101 27285 29135 27319
rect 29135 27285 29144 27319
rect 29092 27276 29144 27285
rect 31484 27276 31536 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 17592 27115 17644 27124
rect 17592 27081 17601 27115
rect 17601 27081 17635 27115
rect 17635 27081 17644 27115
rect 17592 27072 17644 27081
rect 18972 27072 19024 27124
rect 19248 27072 19300 27124
rect 19984 27072 20036 27124
rect 20444 27072 20496 27124
rect 24400 27072 24452 27124
rect 24492 27115 24544 27124
rect 24492 27081 24501 27115
rect 24501 27081 24535 27115
rect 24535 27081 24544 27115
rect 24492 27072 24544 27081
rect 13360 26979 13412 26988
rect 13360 26945 13369 26979
rect 13369 26945 13403 26979
rect 13403 26945 13412 26979
rect 13360 26936 13412 26945
rect 13176 26911 13228 26920
rect 13176 26877 13185 26911
rect 13185 26877 13219 26911
rect 13219 26877 13228 26911
rect 13176 26868 13228 26877
rect 17500 26936 17552 26988
rect 18788 26979 18840 26988
rect 18788 26945 18797 26979
rect 18797 26945 18831 26979
rect 18831 26945 18840 26979
rect 18788 26936 18840 26945
rect 19064 26979 19116 26988
rect 19064 26945 19073 26979
rect 19073 26945 19107 26979
rect 19107 26945 19116 26979
rect 19064 26936 19116 26945
rect 20260 27004 20312 27056
rect 18880 26868 18932 26920
rect 19340 26800 19392 26852
rect 13544 26775 13596 26784
rect 13544 26741 13553 26775
rect 13553 26741 13587 26775
rect 13587 26741 13596 26775
rect 13544 26732 13596 26741
rect 15936 26732 15988 26784
rect 16120 26732 16172 26784
rect 17224 26732 17276 26784
rect 18512 26732 18564 26784
rect 18788 26732 18840 26784
rect 19248 26732 19300 26784
rect 20076 26936 20128 26988
rect 20996 27004 21048 27056
rect 22100 27004 22152 27056
rect 25136 27072 25188 27124
rect 26148 27072 26200 27124
rect 26240 27072 26292 27124
rect 26332 27072 26384 27124
rect 28540 27072 28592 27124
rect 29092 27072 29144 27124
rect 29644 27072 29696 27124
rect 29828 27072 29880 27124
rect 31484 27072 31536 27124
rect 32128 27072 32180 27124
rect 32588 27115 32640 27124
rect 32588 27081 32597 27115
rect 32597 27081 32631 27115
rect 32631 27081 32640 27115
rect 32588 27072 32640 27081
rect 25228 27004 25280 27056
rect 25412 27004 25464 27056
rect 25872 27004 25924 27056
rect 21272 26979 21324 26988
rect 21272 26945 21281 26979
rect 21281 26945 21315 26979
rect 21315 26945 21324 26979
rect 21272 26936 21324 26945
rect 21364 26979 21416 26988
rect 21364 26945 21373 26979
rect 21373 26945 21407 26979
rect 21407 26945 21416 26979
rect 21364 26936 21416 26945
rect 22468 26936 22520 26988
rect 23204 26979 23256 26988
rect 23204 26945 23213 26979
rect 23213 26945 23247 26979
rect 23247 26945 23256 26979
rect 23204 26936 23256 26945
rect 24308 26936 24360 26988
rect 24768 26936 24820 26988
rect 25136 26936 25188 26988
rect 26056 26979 26108 26988
rect 26056 26945 26065 26979
rect 26065 26945 26099 26979
rect 26099 26945 26108 26979
rect 26056 26936 26108 26945
rect 26332 26979 26384 26988
rect 26332 26945 26341 26979
rect 26341 26945 26375 26979
rect 26375 26945 26384 26979
rect 26332 26936 26384 26945
rect 22192 26800 22244 26852
rect 25688 26911 25740 26920
rect 25688 26877 25697 26911
rect 25697 26877 25731 26911
rect 25731 26877 25740 26911
rect 25688 26868 25740 26877
rect 26792 26979 26844 26988
rect 26792 26945 26801 26979
rect 26801 26945 26835 26979
rect 26835 26945 26844 26979
rect 26792 26936 26844 26945
rect 27068 26936 27120 26988
rect 27252 26936 27304 26988
rect 31300 26936 31352 26988
rect 31668 26936 31720 26988
rect 32312 26979 32364 26988
rect 32312 26945 32321 26979
rect 32321 26945 32355 26979
rect 32355 26945 32364 26979
rect 32312 26936 32364 26945
rect 34704 26979 34756 26988
rect 34704 26945 34713 26979
rect 34713 26945 34747 26979
rect 34747 26945 34756 26979
rect 34704 26936 34756 26945
rect 34796 26936 34848 26988
rect 29644 26911 29696 26920
rect 29644 26877 29653 26911
rect 29653 26877 29687 26911
rect 29687 26877 29696 26911
rect 29644 26868 29696 26877
rect 22928 26732 22980 26784
rect 23572 26732 23624 26784
rect 25044 26775 25096 26784
rect 25044 26741 25053 26775
rect 25053 26741 25087 26775
rect 25087 26741 25096 26775
rect 25044 26732 25096 26741
rect 25872 26732 25924 26784
rect 26516 26843 26568 26852
rect 26516 26809 26525 26843
rect 26525 26809 26559 26843
rect 26559 26809 26568 26843
rect 26516 26800 26568 26809
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 13176 26528 13228 26580
rect 13544 26528 13596 26580
rect 16396 26528 16448 26580
rect 20996 26528 21048 26580
rect 22192 26571 22244 26580
rect 22192 26537 22201 26571
rect 22201 26537 22235 26571
rect 22235 26537 22244 26571
rect 22192 26528 22244 26537
rect 22468 26571 22520 26580
rect 22468 26537 22477 26571
rect 22477 26537 22511 26571
rect 22511 26537 22520 26571
rect 22468 26528 22520 26537
rect 24676 26528 24728 26580
rect 25964 26528 26016 26580
rect 32588 26571 32640 26580
rect 32588 26537 32597 26571
rect 32597 26537 32631 26571
rect 32631 26537 32640 26571
rect 32588 26528 32640 26537
rect 34704 26528 34756 26580
rect 13268 26460 13320 26512
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 11980 26324 12032 26376
rect 12992 26367 13044 26376
rect 12992 26333 13001 26367
rect 13001 26333 13035 26367
rect 13035 26333 13044 26367
rect 12992 26324 13044 26333
rect 13084 26324 13136 26376
rect 17040 26460 17092 26512
rect 18144 26392 18196 26444
rect 11060 26256 11112 26308
rect 12532 26256 12584 26308
rect 1860 26188 1912 26240
rect 9496 26231 9548 26240
rect 9496 26197 9505 26231
rect 9505 26197 9539 26231
rect 9539 26197 9548 26231
rect 9496 26188 9548 26197
rect 12716 26231 12768 26240
rect 12716 26197 12725 26231
rect 12725 26197 12759 26231
rect 12759 26197 12768 26231
rect 12716 26188 12768 26197
rect 13636 26188 13688 26240
rect 13912 26188 13964 26240
rect 15936 26256 15988 26308
rect 16488 26367 16540 26376
rect 16488 26333 16497 26367
rect 16497 26333 16531 26367
rect 16531 26333 16540 26367
rect 16488 26324 16540 26333
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 17408 26367 17460 26376
rect 17408 26333 17417 26367
rect 17417 26333 17451 26367
rect 17451 26333 17460 26367
rect 17408 26324 17460 26333
rect 18512 26324 18564 26376
rect 19340 26392 19392 26444
rect 16580 26256 16632 26308
rect 18788 26367 18840 26376
rect 18788 26333 18797 26367
rect 18797 26333 18831 26367
rect 18831 26333 18840 26367
rect 18788 26324 18840 26333
rect 19064 26324 19116 26376
rect 19156 26324 19208 26376
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 16304 26188 16356 26240
rect 17132 26188 17184 26240
rect 18236 26188 18288 26240
rect 21088 26435 21140 26444
rect 21088 26401 21097 26435
rect 21097 26401 21131 26435
rect 21131 26401 21140 26435
rect 21088 26392 21140 26401
rect 22928 26392 22980 26444
rect 23756 26392 23808 26444
rect 21456 26299 21508 26308
rect 21456 26265 21465 26299
rect 21465 26265 21499 26299
rect 21499 26265 21508 26299
rect 21456 26256 21508 26265
rect 23296 26324 23348 26376
rect 23572 26367 23624 26376
rect 23572 26333 23581 26367
rect 23581 26333 23615 26367
rect 23615 26333 23624 26367
rect 23572 26324 23624 26333
rect 24308 26460 24360 26512
rect 25688 26367 25740 26376
rect 25688 26333 25717 26367
rect 25717 26333 25740 26367
rect 25688 26324 25740 26333
rect 25872 26367 25924 26376
rect 25872 26333 25881 26367
rect 25881 26333 25915 26367
rect 25915 26333 25924 26367
rect 25872 26324 25924 26333
rect 26056 26367 26108 26376
rect 26056 26333 26065 26367
rect 26065 26333 26099 26367
rect 26099 26333 26108 26367
rect 26056 26324 26108 26333
rect 27252 26324 27304 26376
rect 34520 26324 34572 26376
rect 20720 26231 20772 26240
rect 20720 26197 20729 26231
rect 20729 26197 20763 26231
rect 20763 26197 20772 26231
rect 20720 26188 20772 26197
rect 21364 26188 21416 26240
rect 22192 26188 22244 26240
rect 26240 26256 26292 26308
rect 27068 26256 27120 26308
rect 33048 26299 33100 26308
rect 33048 26265 33057 26299
rect 33057 26265 33091 26299
rect 33091 26265 33100 26299
rect 33048 26256 33100 26265
rect 26332 26188 26384 26240
rect 30656 26188 30708 26240
rect 31300 26231 31352 26240
rect 31300 26197 31309 26231
rect 31309 26197 31343 26231
rect 31343 26197 31352 26231
rect 31300 26188 31352 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 13360 25984 13412 26036
rect 9404 25848 9456 25900
rect 10232 25848 10284 25900
rect 11336 25848 11388 25900
rect 11980 25916 12032 25968
rect 13728 25984 13780 26036
rect 16488 25984 16540 26036
rect 16580 25984 16632 26036
rect 18236 25984 18288 26036
rect 19432 26027 19484 26036
rect 19432 25993 19441 26027
rect 19441 25993 19475 26027
rect 19475 25993 19484 26027
rect 19432 25984 19484 25993
rect 21272 25984 21324 26036
rect 27252 26027 27304 26036
rect 27252 25993 27261 26027
rect 27261 25993 27295 26027
rect 27295 25993 27304 26027
rect 27252 25984 27304 25993
rect 8852 25644 8904 25696
rect 9496 25644 9548 25696
rect 9864 25644 9916 25696
rect 11704 25780 11756 25832
rect 11888 25780 11940 25832
rect 12532 25891 12584 25900
rect 12532 25857 12541 25891
rect 12541 25857 12575 25891
rect 12575 25857 12584 25891
rect 12532 25848 12584 25857
rect 12808 25891 12860 25900
rect 12808 25857 12817 25891
rect 12817 25857 12851 25891
rect 12851 25857 12860 25891
rect 12808 25848 12860 25857
rect 12992 25891 13044 25900
rect 12992 25857 13001 25891
rect 13001 25857 13035 25891
rect 13035 25857 13044 25891
rect 12992 25848 13044 25857
rect 13452 25891 13504 25900
rect 13452 25857 13461 25891
rect 13461 25857 13495 25891
rect 13495 25857 13504 25891
rect 13452 25848 13504 25857
rect 13636 25891 13688 25900
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 12716 25780 12768 25832
rect 13820 25891 13872 25900
rect 13820 25857 13829 25891
rect 13829 25857 13863 25891
rect 13863 25857 13872 25891
rect 13820 25848 13872 25857
rect 14096 25891 14148 25900
rect 14096 25857 14105 25891
rect 14105 25857 14139 25891
rect 14139 25857 14148 25891
rect 14096 25848 14148 25857
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 12900 25712 12952 25764
rect 14464 25755 14516 25764
rect 14464 25721 14473 25755
rect 14473 25721 14507 25755
rect 14507 25721 14516 25755
rect 14464 25712 14516 25721
rect 16028 25916 16080 25968
rect 15752 25848 15804 25900
rect 16120 25891 16172 25900
rect 16120 25857 16129 25891
rect 16129 25857 16163 25891
rect 16163 25857 16172 25891
rect 16120 25848 16172 25857
rect 16396 25848 16448 25900
rect 17592 25916 17644 25968
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 18144 25916 18196 25968
rect 19064 25916 19116 25968
rect 16212 25780 16264 25832
rect 18328 25823 18380 25832
rect 18328 25789 18337 25823
rect 18337 25789 18371 25823
rect 18371 25789 18380 25823
rect 18328 25780 18380 25789
rect 18788 25780 18840 25832
rect 19156 25891 19208 25900
rect 19156 25857 19165 25891
rect 19165 25857 19199 25891
rect 19199 25857 19208 25891
rect 19156 25848 19208 25857
rect 19340 25959 19392 25968
rect 19340 25925 19349 25959
rect 19349 25925 19383 25959
rect 19383 25925 19392 25959
rect 19340 25916 19392 25925
rect 26332 25916 26384 25968
rect 29552 25916 29604 25968
rect 31668 25984 31720 26036
rect 33048 25984 33100 26036
rect 30564 25916 30616 25968
rect 20996 25848 21048 25900
rect 26148 25848 26200 25900
rect 16672 25712 16724 25764
rect 19248 25823 19300 25832
rect 19248 25789 19257 25823
rect 19257 25789 19291 25823
rect 19291 25789 19300 25823
rect 19248 25780 19300 25789
rect 27160 25848 27212 25900
rect 27344 25780 27396 25832
rect 13176 25687 13228 25696
rect 13176 25653 13185 25687
rect 13185 25653 13219 25687
rect 13219 25653 13228 25687
rect 13176 25644 13228 25653
rect 13268 25644 13320 25696
rect 13820 25644 13872 25696
rect 14924 25687 14976 25696
rect 14924 25653 14933 25687
rect 14933 25653 14967 25687
rect 14967 25653 14976 25687
rect 14924 25644 14976 25653
rect 15660 25644 15712 25696
rect 15936 25644 15988 25696
rect 16028 25687 16080 25696
rect 16028 25653 16037 25687
rect 16037 25653 16071 25687
rect 16071 25653 16080 25687
rect 16028 25644 16080 25653
rect 16488 25644 16540 25696
rect 16580 25644 16632 25696
rect 20904 25644 20956 25696
rect 21272 25644 21324 25696
rect 22376 25687 22428 25696
rect 22376 25653 22385 25687
rect 22385 25653 22419 25687
rect 22419 25653 22428 25687
rect 22376 25644 22428 25653
rect 22652 25687 22704 25696
rect 22652 25653 22661 25687
rect 22661 25653 22695 25687
rect 22695 25653 22704 25687
rect 22652 25644 22704 25653
rect 22928 25644 22980 25696
rect 23296 25712 23348 25764
rect 28080 25712 28132 25764
rect 23388 25687 23440 25696
rect 23388 25653 23397 25687
rect 23397 25653 23431 25687
rect 23431 25653 23440 25687
rect 23388 25644 23440 25653
rect 31852 25823 31904 25832
rect 31852 25789 31861 25823
rect 31861 25789 31895 25823
rect 31895 25789 31904 25823
rect 31852 25780 31904 25789
rect 32220 25823 32272 25832
rect 32220 25789 32229 25823
rect 32229 25789 32263 25823
rect 32263 25789 32272 25823
rect 32220 25780 32272 25789
rect 31760 25712 31812 25764
rect 34520 25687 34572 25696
rect 34520 25653 34529 25687
rect 34529 25653 34563 25687
rect 34563 25653 34572 25687
rect 34520 25644 34572 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 9680 25372 9732 25424
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 9404 25236 9456 25288
rect 9496 25279 9548 25288
rect 9496 25245 9505 25279
rect 9505 25245 9539 25279
rect 9539 25245 9548 25279
rect 9496 25236 9548 25245
rect 10232 25279 10284 25288
rect 10232 25245 10241 25279
rect 10241 25245 10275 25279
rect 10275 25245 10284 25279
rect 10232 25236 10284 25245
rect 11060 25236 11112 25288
rect 13176 25440 13228 25492
rect 13360 25440 13412 25492
rect 13728 25440 13780 25492
rect 14096 25440 14148 25492
rect 14924 25440 14976 25492
rect 15844 25440 15896 25492
rect 11704 25372 11756 25424
rect 11888 25304 11940 25356
rect 12808 25372 12860 25424
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 9036 25168 9088 25220
rect 10416 25211 10468 25220
rect 10416 25177 10425 25211
rect 10425 25177 10459 25211
rect 10459 25177 10468 25211
rect 10416 25168 10468 25177
rect 10876 25168 10928 25220
rect 11336 25168 11388 25220
rect 12992 25236 13044 25288
rect 13268 25236 13320 25288
rect 13452 25372 13504 25424
rect 13912 25372 13964 25424
rect 8852 25100 8904 25152
rect 10508 25100 10560 25152
rect 11244 25100 11296 25152
rect 12072 25143 12124 25152
rect 12072 25109 12081 25143
rect 12081 25109 12115 25143
rect 12115 25109 12124 25143
rect 12072 25100 12124 25109
rect 12256 25100 12308 25152
rect 12348 25100 12400 25152
rect 12808 25100 12860 25152
rect 12992 25100 13044 25152
rect 13636 25168 13688 25220
rect 16580 25440 16632 25492
rect 17040 25440 17092 25492
rect 23664 25440 23716 25492
rect 23756 25483 23808 25492
rect 23756 25449 23765 25483
rect 23765 25449 23799 25483
rect 23799 25449 23808 25483
rect 23756 25440 23808 25449
rect 24860 25483 24912 25492
rect 24860 25449 24869 25483
rect 24869 25449 24903 25483
rect 24903 25449 24912 25483
rect 24860 25440 24912 25449
rect 30564 25483 30616 25492
rect 30564 25449 30573 25483
rect 30573 25449 30607 25483
rect 30607 25449 30616 25483
rect 30564 25440 30616 25449
rect 32220 25440 32272 25492
rect 14096 25236 14148 25288
rect 15292 25279 15344 25288
rect 15292 25245 15301 25279
rect 15301 25245 15335 25279
rect 15335 25245 15344 25279
rect 15292 25236 15344 25245
rect 16120 25372 16172 25424
rect 15568 25347 15620 25356
rect 15568 25313 15577 25347
rect 15577 25313 15611 25347
rect 15611 25313 15620 25347
rect 15568 25304 15620 25313
rect 16212 25304 16264 25356
rect 16304 25347 16356 25356
rect 16304 25313 16313 25347
rect 16313 25313 16347 25347
rect 16347 25313 16356 25347
rect 16304 25304 16356 25313
rect 16672 25304 16724 25356
rect 15752 25236 15804 25288
rect 20720 25372 20772 25424
rect 20904 25236 20956 25288
rect 22652 25372 22704 25424
rect 21824 25347 21876 25356
rect 21824 25313 21833 25347
rect 21833 25313 21867 25347
rect 21867 25313 21876 25347
rect 21824 25304 21876 25313
rect 23296 25372 23348 25424
rect 22928 25236 22980 25288
rect 23204 25279 23256 25288
rect 23204 25245 23213 25279
rect 23213 25245 23247 25279
rect 23247 25245 23256 25279
rect 23204 25236 23256 25245
rect 24768 25304 24820 25356
rect 26148 25304 26200 25356
rect 27344 25304 27396 25356
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 13728 25100 13780 25152
rect 13820 25100 13872 25152
rect 16212 25143 16264 25152
rect 16212 25109 16221 25143
rect 16221 25109 16255 25143
rect 16255 25109 16264 25143
rect 16212 25100 16264 25109
rect 20076 25143 20128 25152
rect 20076 25109 20085 25143
rect 20085 25109 20119 25143
rect 20119 25109 20128 25143
rect 20076 25100 20128 25109
rect 20444 25143 20496 25152
rect 20444 25109 20453 25143
rect 20453 25109 20487 25143
rect 20487 25109 20496 25143
rect 20444 25100 20496 25109
rect 20812 25143 20864 25152
rect 20812 25109 20821 25143
rect 20821 25109 20855 25143
rect 20855 25109 20864 25143
rect 20812 25100 20864 25109
rect 21272 25143 21324 25152
rect 21272 25109 21281 25143
rect 21281 25109 21315 25143
rect 21315 25109 21324 25143
rect 21272 25100 21324 25109
rect 21732 25100 21784 25152
rect 23296 25211 23348 25220
rect 23296 25177 23305 25211
rect 23305 25177 23339 25211
rect 23339 25177 23348 25211
rect 23296 25168 23348 25177
rect 24032 25279 24084 25288
rect 24032 25245 24041 25279
rect 24041 25245 24075 25279
rect 24075 25245 24084 25279
rect 24032 25236 24084 25245
rect 24400 25279 24452 25288
rect 24400 25245 24409 25279
rect 24409 25245 24443 25279
rect 24443 25245 24452 25279
rect 24400 25236 24452 25245
rect 24860 25236 24912 25288
rect 25780 25236 25832 25288
rect 25964 25279 26016 25288
rect 25964 25245 25973 25279
rect 25973 25245 26007 25279
rect 26007 25245 26016 25279
rect 25964 25236 26016 25245
rect 32312 25304 32364 25356
rect 27620 25279 27672 25288
rect 27620 25245 27629 25279
rect 27629 25245 27663 25279
rect 27663 25245 27672 25279
rect 27620 25236 27672 25245
rect 27804 25236 27856 25288
rect 24308 25100 24360 25152
rect 27344 25143 27396 25152
rect 27344 25109 27353 25143
rect 27353 25109 27387 25143
rect 27387 25109 27396 25143
rect 27344 25100 27396 25109
rect 31760 25236 31812 25288
rect 31852 25279 31904 25288
rect 31852 25245 31861 25279
rect 31861 25245 31895 25279
rect 31895 25245 31904 25279
rect 31852 25236 31904 25245
rect 32956 25236 33008 25288
rect 34888 25236 34940 25288
rect 34060 25168 34112 25220
rect 30656 25100 30708 25152
rect 31944 25100 31996 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9404 24896 9456 24948
rect 11336 24939 11388 24948
rect 11336 24905 11345 24939
rect 11345 24905 11379 24939
rect 11379 24905 11388 24939
rect 11336 24896 11388 24905
rect 11704 24896 11756 24948
rect 12348 24896 12400 24948
rect 15660 24896 15712 24948
rect 16212 24896 16264 24948
rect 20812 24896 20864 24948
rect 8576 24760 8628 24812
rect 8852 24828 8904 24880
rect 9036 24803 9088 24812
rect 9036 24769 9045 24803
rect 9045 24769 9079 24803
rect 9079 24769 9088 24803
rect 9036 24760 9088 24769
rect 9220 24760 9272 24812
rect 12440 24828 12492 24880
rect 13728 24760 13780 24812
rect 15660 24803 15712 24812
rect 15660 24769 15669 24803
rect 15669 24769 15703 24803
rect 15703 24769 15712 24803
rect 15660 24760 15712 24769
rect 8852 24624 8904 24676
rect 10784 24556 10836 24608
rect 13820 24692 13872 24744
rect 15200 24692 15252 24744
rect 15936 24760 15988 24812
rect 20996 24828 21048 24880
rect 21088 24828 21140 24880
rect 21824 24896 21876 24948
rect 22376 24896 22428 24948
rect 23204 24896 23256 24948
rect 23756 24896 23808 24948
rect 24860 24939 24912 24948
rect 24860 24905 24869 24939
rect 24869 24905 24903 24939
rect 24903 24905 24912 24939
rect 24860 24896 24912 24905
rect 22468 24828 22520 24880
rect 22652 24871 22704 24880
rect 22652 24837 22661 24871
rect 22661 24837 22695 24871
rect 22695 24837 22704 24871
rect 22652 24828 22704 24837
rect 18328 24760 18380 24812
rect 19340 24760 19392 24812
rect 19984 24803 20036 24812
rect 19984 24769 19993 24803
rect 19993 24769 20027 24803
rect 20027 24769 20036 24803
rect 19984 24760 20036 24769
rect 20444 24760 20496 24812
rect 15844 24735 15896 24744
rect 15844 24701 15853 24735
rect 15853 24701 15887 24735
rect 15887 24701 15896 24735
rect 15844 24692 15896 24701
rect 19064 24735 19116 24744
rect 19064 24701 19073 24735
rect 19073 24701 19107 24735
rect 19107 24701 19116 24735
rect 19064 24692 19116 24701
rect 11060 24624 11112 24676
rect 13084 24624 13136 24676
rect 12440 24556 12492 24608
rect 12716 24556 12768 24608
rect 15384 24624 15436 24676
rect 15752 24624 15804 24676
rect 16396 24624 16448 24676
rect 16488 24624 16540 24676
rect 17960 24624 18012 24676
rect 21364 24624 21416 24676
rect 22100 24667 22152 24676
rect 22100 24633 22109 24667
rect 22109 24633 22143 24667
rect 22143 24633 22152 24667
rect 22100 24624 22152 24633
rect 13728 24556 13780 24608
rect 22468 24599 22520 24608
rect 22468 24565 22477 24599
rect 22477 24565 22511 24599
rect 22511 24565 22520 24599
rect 29644 24939 29696 24948
rect 29644 24905 29653 24939
rect 29653 24905 29687 24939
rect 29687 24905 29696 24939
rect 29644 24896 29696 24905
rect 34888 24939 34940 24948
rect 34888 24905 34897 24939
rect 34897 24905 34931 24939
rect 34931 24905 34940 24939
rect 34888 24896 34940 24905
rect 23756 24803 23808 24812
rect 23756 24769 23765 24803
rect 23765 24769 23799 24803
rect 23799 24769 23808 24803
rect 23756 24760 23808 24769
rect 24032 24803 24084 24812
rect 24032 24769 24041 24803
rect 24041 24769 24075 24803
rect 24075 24769 24084 24803
rect 24032 24760 24084 24769
rect 23664 24624 23716 24676
rect 24308 24803 24360 24812
rect 24308 24769 24317 24803
rect 24317 24769 24351 24803
rect 24351 24769 24360 24803
rect 24308 24760 24360 24769
rect 24952 24760 25004 24812
rect 25780 24828 25832 24880
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 22468 24556 22520 24565
rect 23204 24556 23256 24608
rect 25964 24692 26016 24744
rect 31760 24760 31812 24812
rect 31944 24760 31996 24812
rect 34152 24828 34204 24880
rect 32956 24803 33008 24812
rect 32956 24769 32973 24803
rect 32973 24769 33007 24803
rect 33007 24769 33008 24803
rect 32956 24760 33008 24769
rect 33048 24692 33100 24744
rect 25596 24624 25648 24676
rect 27160 24556 27212 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 9220 24352 9272 24404
rect 11152 24352 11204 24404
rect 12716 24352 12768 24404
rect 10416 24259 10468 24268
rect 10416 24225 10425 24259
rect 10425 24225 10459 24259
rect 10459 24225 10468 24259
rect 10416 24216 10468 24225
rect 940 24148 992 24200
rect 4068 24148 4120 24200
rect 9036 24148 9088 24200
rect 11888 24284 11940 24336
rect 12072 24284 12124 24336
rect 15200 24352 15252 24404
rect 15292 24395 15344 24404
rect 15292 24361 15301 24395
rect 15301 24361 15335 24395
rect 15335 24361 15344 24395
rect 15292 24352 15344 24361
rect 15844 24352 15896 24404
rect 17132 24352 17184 24404
rect 10692 24216 10744 24268
rect 11060 24148 11112 24200
rect 11244 24191 11296 24200
rect 11244 24157 11253 24191
rect 11253 24157 11287 24191
rect 11287 24157 11296 24191
rect 11244 24148 11296 24157
rect 2044 24012 2096 24064
rect 2964 24055 3016 24064
rect 2964 24021 2973 24055
rect 2973 24021 3007 24055
rect 3007 24021 3016 24055
rect 2964 24012 3016 24021
rect 3424 24055 3476 24064
rect 3424 24021 3433 24055
rect 3433 24021 3467 24055
rect 3467 24021 3476 24055
rect 3424 24012 3476 24021
rect 6644 24012 6696 24064
rect 10692 24080 10744 24132
rect 11888 24191 11940 24200
rect 11888 24157 11897 24191
rect 11897 24157 11931 24191
rect 11931 24157 11940 24191
rect 11888 24148 11940 24157
rect 12808 24216 12860 24268
rect 13084 24284 13136 24336
rect 15752 24284 15804 24336
rect 16304 24284 16356 24336
rect 14004 24216 14056 24268
rect 12532 24148 12584 24200
rect 13084 24148 13136 24200
rect 13176 24148 13228 24200
rect 15292 24216 15344 24268
rect 16396 24259 16448 24268
rect 16396 24225 16405 24259
rect 16405 24225 16439 24259
rect 16439 24225 16448 24259
rect 16396 24216 16448 24225
rect 14556 24148 14608 24200
rect 15476 24191 15528 24200
rect 15476 24157 15485 24191
rect 15485 24157 15519 24191
rect 15519 24157 15528 24191
rect 15476 24148 15528 24157
rect 15752 24191 15804 24200
rect 15752 24157 15761 24191
rect 15761 24157 15795 24191
rect 15795 24157 15804 24191
rect 15752 24148 15804 24157
rect 22192 24352 22244 24404
rect 22376 24352 22428 24404
rect 22836 24352 22888 24404
rect 25872 24352 25924 24404
rect 28080 24352 28132 24404
rect 18236 24259 18288 24268
rect 18236 24225 18245 24259
rect 18245 24225 18279 24259
rect 18279 24225 18288 24259
rect 18236 24216 18288 24225
rect 12164 24080 12216 24132
rect 12348 24080 12400 24132
rect 20260 24284 20312 24336
rect 21088 24284 21140 24336
rect 20996 24148 21048 24200
rect 21732 24148 21784 24200
rect 22192 24148 22244 24200
rect 25596 24191 25648 24200
rect 25596 24157 25605 24191
rect 25605 24157 25639 24191
rect 25639 24157 25648 24191
rect 25596 24148 25648 24157
rect 11980 24055 12032 24064
rect 11980 24021 11989 24055
rect 11989 24021 12023 24055
rect 12023 24021 12032 24055
rect 11980 24012 12032 24021
rect 12808 24012 12860 24064
rect 21364 24123 21416 24132
rect 21364 24089 21373 24123
rect 21373 24089 21407 24123
rect 21407 24089 21416 24123
rect 27068 24327 27120 24336
rect 27068 24293 27077 24327
rect 27077 24293 27111 24327
rect 27111 24293 27120 24327
rect 27068 24284 27120 24293
rect 27344 24216 27396 24268
rect 27620 24216 27672 24268
rect 26976 24191 27028 24200
rect 26976 24157 26985 24191
rect 26985 24157 27019 24191
rect 27019 24157 27028 24191
rect 26976 24148 27028 24157
rect 27436 24191 27488 24200
rect 27436 24157 27445 24191
rect 27445 24157 27479 24191
rect 27479 24157 27488 24191
rect 27436 24148 27488 24157
rect 21364 24080 21416 24089
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 14372 24012 14424 24064
rect 20076 24012 20128 24064
rect 20444 24012 20496 24064
rect 22192 24055 22244 24064
rect 22192 24021 22201 24055
rect 22201 24021 22235 24055
rect 22235 24021 22244 24055
rect 22192 24012 22244 24021
rect 22928 24012 22980 24064
rect 23388 24055 23440 24064
rect 23388 24021 23397 24055
rect 23397 24021 23431 24055
rect 23431 24021 23440 24055
rect 23388 24012 23440 24021
rect 27804 24080 27856 24132
rect 27988 24080 28040 24132
rect 28724 24284 28776 24336
rect 27528 24012 27580 24064
rect 29092 24259 29144 24268
rect 29092 24225 29101 24259
rect 29101 24225 29135 24259
rect 29135 24225 29144 24259
rect 29092 24216 29144 24225
rect 31944 24352 31996 24404
rect 34152 24352 34204 24404
rect 29644 24216 29696 24268
rect 28632 24191 28684 24200
rect 28632 24157 28641 24191
rect 28641 24157 28675 24191
rect 28675 24157 28684 24191
rect 28632 24148 28684 24157
rect 29000 24191 29052 24200
rect 29000 24157 29009 24191
rect 29009 24157 29043 24191
rect 29043 24157 29052 24191
rect 29000 24148 29052 24157
rect 29368 24148 29420 24200
rect 28908 24012 28960 24064
rect 30840 24080 30892 24132
rect 34520 24148 34572 24200
rect 32680 24012 32732 24064
rect 33048 24012 33100 24064
rect 34060 24055 34112 24064
rect 34060 24021 34069 24055
rect 34069 24021 34103 24055
rect 34103 24021 34112 24055
rect 34060 24012 34112 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 11704 23851 11756 23860
rect 11704 23817 11713 23851
rect 11713 23817 11747 23851
rect 11747 23817 11756 23851
rect 11704 23808 11756 23817
rect 11980 23808 12032 23860
rect 12348 23808 12400 23860
rect 13176 23808 13228 23860
rect 15476 23808 15528 23860
rect 15752 23808 15804 23860
rect 15844 23808 15896 23860
rect 18236 23808 18288 23860
rect 20536 23808 20588 23860
rect 21732 23808 21784 23860
rect 1860 23783 1912 23792
rect 1860 23749 1869 23783
rect 1869 23749 1903 23783
rect 1903 23749 1912 23783
rect 1860 23740 1912 23749
rect 3700 23783 3752 23792
rect 3700 23749 3709 23783
rect 3709 23749 3743 23783
rect 3743 23749 3752 23783
rect 3700 23740 3752 23749
rect 4712 23740 4764 23792
rect 2964 23672 3016 23724
rect 3424 23715 3476 23724
rect 3424 23681 3433 23715
rect 3433 23681 3467 23715
rect 3467 23681 3476 23715
rect 3424 23672 3476 23681
rect 6644 23740 6696 23792
rect 8300 23740 8352 23792
rect 10968 23740 11020 23792
rect 1400 23604 1452 23656
rect 5356 23647 5408 23656
rect 5356 23613 5365 23647
rect 5365 23613 5399 23647
rect 5399 23613 5408 23647
rect 5356 23604 5408 23613
rect 10600 23672 10652 23724
rect 4804 23468 4856 23520
rect 5172 23511 5224 23520
rect 5172 23477 5181 23511
rect 5181 23477 5215 23511
rect 5215 23477 5224 23511
rect 5172 23468 5224 23477
rect 10232 23468 10284 23520
rect 10600 23468 10652 23520
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 12532 23672 12584 23724
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 14556 23740 14608 23792
rect 14280 23672 14332 23724
rect 15292 23672 15344 23724
rect 15384 23672 15436 23724
rect 15752 23715 15804 23724
rect 15752 23681 15761 23715
rect 15761 23681 15795 23715
rect 15795 23681 15804 23715
rect 15752 23672 15804 23681
rect 12164 23536 12216 23588
rect 14004 23647 14056 23656
rect 14004 23613 14013 23647
rect 14013 23613 14047 23647
rect 14047 23613 14056 23647
rect 14004 23604 14056 23613
rect 16488 23672 16540 23724
rect 17960 23740 18012 23792
rect 21088 23740 21140 23792
rect 23664 23808 23716 23860
rect 17592 23672 17644 23724
rect 16304 23604 16356 23656
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20536 23715 20588 23724
rect 20536 23681 20545 23715
rect 20545 23681 20579 23715
rect 20579 23681 20588 23715
rect 20536 23672 20588 23681
rect 22100 23672 22152 23724
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22468 23715 22520 23724
rect 22468 23681 22477 23715
rect 22477 23681 22511 23715
rect 22511 23681 22520 23715
rect 22468 23672 22520 23681
rect 10784 23468 10836 23477
rect 12440 23468 12492 23520
rect 15200 23468 15252 23520
rect 17132 23511 17184 23520
rect 17132 23477 17141 23511
rect 17141 23477 17175 23511
rect 17175 23477 17184 23511
rect 17132 23468 17184 23477
rect 19248 23468 19300 23520
rect 21824 23647 21876 23656
rect 21824 23613 21833 23647
rect 21833 23613 21867 23647
rect 21867 23613 21876 23647
rect 21824 23604 21876 23613
rect 23388 23740 23440 23792
rect 22652 23715 22704 23724
rect 22652 23681 22661 23715
rect 22661 23681 22695 23715
rect 22695 23681 22704 23715
rect 22652 23672 22704 23681
rect 22744 23715 22796 23724
rect 22744 23681 22753 23715
rect 22753 23681 22787 23715
rect 22787 23681 22796 23715
rect 22744 23672 22796 23681
rect 22836 23672 22888 23724
rect 24492 23672 24544 23724
rect 25044 23740 25096 23792
rect 26976 23851 27028 23860
rect 26976 23817 26985 23851
rect 26985 23817 27019 23851
rect 27019 23817 27028 23851
rect 26976 23808 27028 23817
rect 27160 23851 27212 23860
rect 27160 23817 27187 23851
rect 27187 23817 27212 23851
rect 27160 23808 27212 23817
rect 28632 23808 28684 23860
rect 28724 23808 28776 23860
rect 28908 23808 28960 23860
rect 29000 23851 29052 23860
rect 29000 23817 29009 23851
rect 29009 23817 29043 23851
rect 29043 23817 29052 23851
rect 29000 23808 29052 23817
rect 29092 23808 29144 23860
rect 30840 23851 30892 23860
rect 30840 23817 30849 23851
rect 30849 23817 30883 23851
rect 30883 23817 30892 23851
rect 30840 23808 30892 23817
rect 25596 23740 25648 23792
rect 27436 23740 27488 23792
rect 27804 23740 27856 23792
rect 28356 23783 28408 23792
rect 28356 23749 28365 23783
rect 28365 23749 28399 23783
rect 28399 23749 28408 23783
rect 28356 23740 28408 23749
rect 27988 23604 28040 23656
rect 21272 23468 21324 23520
rect 22744 23468 22796 23520
rect 23020 23468 23072 23520
rect 23204 23468 23256 23520
rect 24308 23468 24360 23520
rect 24860 23468 24912 23520
rect 27252 23468 27304 23520
rect 27528 23468 27580 23520
rect 29092 23715 29144 23724
rect 29092 23681 29101 23715
rect 29101 23681 29135 23715
rect 29135 23681 29144 23715
rect 29092 23672 29144 23681
rect 29368 23715 29420 23724
rect 29368 23681 29377 23715
rect 29377 23681 29411 23715
rect 29411 23681 29420 23715
rect 29368 23672 29420 23681
rect 30656 23511 30708 23520
rect 30656 23477 30665 23511
rect 30665 23477 30699 23511
rect 30699 23477 30708 23511
rect 30656 23468 30708 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 3424 23307 3476 23316
rect 3424 23273 3433 23307
rect 3433 23273 3467 23307
rect 3467 23273 3476 23307
rect 3424 23264 3476 23273
rect 4712 23264 4764 23316
rect 8300 23307 8352 23316
rect 8300 23273 8309 23307
rect 8309 23273 8343 23307
rect 8343 23273 8352 23307
rect 8300 23264 8352 23273
rect 8852 23264 8904 23316
rect 1676 23171 1728 23180
rect 1676 23137 1685 23171
rect 1685 23137 1719 23171
rect 1719 23137 1728 23171
rect 1676 23128 1728 23137
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 2228 22992 2280 23044
rect 4160 23196 4212 23248
rect 5264 23171 5316 23180
rect 5264 23137 5273 23171
rect 5273 23137 5307 23171
rect 5307 23137 5316 23171
rect 5264 23128 5316 23137
rect 6644 23128 6696 23180
rect 13912 23264 13964 23316
rect 14372 23264 14424 23316
rect 15292 23264 15344 23316
rect 15752 23264 15804 23316
rect 19432 23264 19484 23316
rect 19984 23264 20036 23316
rect 20260 23264 20312 23316
rect 21824 23264 21876 23316
rect 22100 23264 22152 23316
rect 4804 23060 4856 23112
rect 5448 23060 5500 23112
rect 8208 23060 8260 23112
rect 15384 23128 15436 23180
rect 17132 23171 17184 23180
rect 17132 23137 17141 23171
rect 17141 23137 17175 23171
rect 17175 23137 17184 23171
rect 17132 23128 17184 23137
rect 10048 23103 10100 23112
rect 10048 23069 10057 23103
rect 10057 23069 10091 23103
rect 10091 23069 10100 23103
rect 10048 23060 10100 23069
rect 10232 23103 10284 23112
rect 10232 23069 10241 23103
rect 10241 23069 10275 23103
rect 10275 23069 10284 23103
rect 10232 23060 10284 23069
rect 15568 23103 15620 23112
rect 15568 23069 15578 23103
rect 15578 23069 15620 23103
rect 22468 23264 22520 23316
rect 22652 23264 22704 23316
rect 23204 23264 23256 23316
rect 24400 23264 24452 23316
rect 24860 23264 24912 23316
rect 15568 23060 15620 23069
rect 2596 22924 2648 22976
rect 4712 22992 4764 23044
rect 7656 22992 7708 23044
rect 11152 22992 11204 23044
rect 15200 22992 15252 23044
rect 12716 22924 12768 22976
rect 14372 22967 14424 22976
rect 14372 22933 14381 22967
rect 14381 22933 14415 22967
rect 14415 22933 14424 22967
rect 14372 22924 14424 22933
rect 18420 23103 18472 23112
rect 18420 23069 18429 23103
rect 18429 23069 18463 23103
rect 18463 23069 18472 23103
rect 18420 23060 18472 23069
rect 18604 22924 18656 22976
rect 19340 22967 19392 22976
rect 19340 22933 19349 22967
rect 19349 22933 19383 22967
rect 19383 22933 19392 22967
rect 19340 22924 19392 22933
rect 20996 23103 21048 23112
rect 20996 23069 21005 23103
rect 21005 23069 21039 23103
rect 21039 23069 21048 23103
rect 20996 23060 21048 23069
rect 21088 23060 21140 23112
rect 23020 23171 23072 23180
rect 23020 23137 23029 23171
rect 23029 23137 23063 23171
rect 23063 23137 23072 23171
rect 23020 23128 23072 23137
rect 21456 22924 21508 22976
rect 21548 22967 21600 22976
rect 21548 22933 21557 22967
rect 21557 22933 21591 22967
rect 21591 22933 21600 22967
rect 21548 22924 21600 22933
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22879 23103
rect 22879 23069 22888 23103
rect 22836 23060 22888 23069
rect 23112 23103 23164 23112
rect 23112 23069 23121 23103
rect 23121 23069 23155 23103
rect 23155 23069 23164 23103
rect 23112 23060 23164 23069
rect 24032 23060 24084 23112
rect 24308 23060 24360 23112
rect 24492 23060 24544 23112
rect 24768 23060 24820 23112
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 25780 23171 25832 23180
rect 25780 23137 25789 23171
rect 25789 23137 25823 23171
rect 25823 23137 25832 23171
rect 25780 23128 25832 23137
rect 22928 22992 22980 23044
rect 22468 22924 22520 22976
rect 22744 22924 22796 22976
rect 22836 22924 22888 22976
rect 24492 22924 24544 22976
rect 34612 22992 34664 23044
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2228 22763 2280 22772
rect 2228 22729 2237 22763
rect 2237 22729 2271 22763
rect 2271 22729 2280 22763
rect 2228 22720 2280 22729
rect 7656 22720 7708 22772
rect 2872 22695 2924 22704
rect 2872 22661 2881 22695
rect 2881 22661 2915 22695
rect 2915 22661 2924 22695
rect 2872 22652 2924 22661
rect 3884 22652 3936 22704
rect 8208 22720 8260 22772
rect 12440 22763 12492 22772
rect 9680 22584 9732 22636
rect 2596 22559 2648 22568
rect 2596 22525 2605 22559
rect 2605 22525 2639 22559
rect 2639 22525 2648 22559
rect 2596 22516 2648 22525
rect 2688 22380 2740 22432
rect 4804 22516 4856 22568
rect 10324 22584 10376 22636
rect 12440 22729 12449 22763
rect 12449 22729 12483 22763
rect 12483 22729 12492 22763
rect 12440 22720 12492 22729
rect 12716 22627 12768 22636
rect 11888 22516 11940 22568
rect 10048 22448 10100 22500
rect 4896 22380 4948 22432
rect 6644 22380 6696 22432
rect 9312 22380 9364 22432
rect 9496 22380 9548 22432
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 10784 22448 10836 22500
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 14096 22720 14148 22772
rect 14280 22720 14332 22772
rect 14464 22720 14516 22772
rect 13452 22627 13504 22636
rect 13452 22593 13461 22627
rect 13461 22593 13495 22627
rect 13495 22593 13504 22627
rect 13452 22584 13504 22593
rect 12992 22448 13044 22500
rect 13912 22627 13964 22636
rect 13912 22593 13921 22627
rect 13921 22593 13955 22627
rect 13955 22593 13964 22627
rect 13912 22584 13964 22593
rect 15568 22720 15620 22772
rect 17592 22720 17644 22772
rect 18604 22720 18656 22772
rect 20904 22720 20956 22772
rect 21180 22720 21232 22772
rect 21548 22720 21600 22772
rect 22836 22720 22888 22772
rect 23020 22720 23072 22772
rect 24492 22720 24544 22772
rect 24860 22720 24912 22772
rect 29644 22720 29696 22772
rect 14188 22516 14240 22568
rect 14372 22516 14424 22568
rect 20996 22584 21048 22636
rect 18052 22516 18104 22568
rect 18420 22516 18472 22568
rect 21732 22516 21784 22568
rect 9772 22380 9824 22389
rect 10600 22423 10652 22432
rect 10600 22389 10609 22423
rect 10609 22389 10643 22423
rect 10643 22389 10652 22423
rect 10600 22380 10652 22389
rect 11060 22380 11112 22432
rect 13268 22423 13320 22432
rect 13268 22389 13277 22423
rect 13277 22389 13311 22423
rect 13311 22389 13320 22423
rect 13268 22380 13320 22389
rect 13452 22380 13504 22432
rect 19524 22448 19576 22500
rect 21456 22448 21508 22500
rect 22192 22584 22244 22636
rect 23296 22695 23348 22704
rect 23296 22661 23305 22695
rect 23305 22661 23339 22695
rect 23339 22661 23348 22695
rect 23296 22652 23348 22661
rect 22560 22627 22612 22636
rect 22560 22593 22569 22627
rect 22569 22593 22603 22627
rect 22603 22593 22612 22627
rect 22560 22584 22612 22593
rect 22376 22559 22428 22568
rect 22376 22525 22385 22559
rect 22385 22525 22419 22559
rect 22419 22525 22428 22559
rect 22376 22516 22428 22525
rect 22836 22516 22888 22568
rect 26240 22584 26292 22636
rect 28448 22584 28500 22636
rect 30932 22652 30984 22704
rect 34152 22652 34204 22704
rect 25044 22516 25096 22568
rect 27620 22516 27672 22568
rect 30380 22559 30432 22568
rect 30380 22525 30389 22559
rect 30389 22525 30423 22559
rect 30423 22525 30432 22559
rect 30380 22516 30432 22525
rect 32036 22584 32088 22636
rect 32496 22584 32548 22636
rect 32956 22627 33008 22636
rect 32956 22593 32965 22627
rect 32965 22593 32999 22627
rect 32999 22593 33008 22627
rect 32956 22584 33008 22593
rect 32588 22448 32640 22500
rect 14280 22423 14332 22432
rect 14280 22389 14289 22423
rect 14289 22389 14323 22423
rect 14323 22389 14332 22423
rect 14280 22380 14332 22389
rect 23112 22423 23164 22432
rect 23112 22389 23121 22423
rect 23121 22389 23155 22423
rect 23155 22389 23164 22423
rect 23112 22380 23164 22389
rect 23388 22380 23440 22432
rect 27528 22423 27580 22432
rect 27528 22389 27537 22423
rect 27537 22389 27571 22423
rect 27571 22389 27580 22423
rect 27528 22380 27580 22389
rect 27896 22423 27948 22432
rect 27896 22389 27905 22423
rect 27905 22389 27939 22423
rect 27939 22389 27948 22423
rect 27896 22380 27948 22389
rect 32680 22380 32732 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3884 22219 3936 22228
rect 3884 22185 3893 22219
rect 3893 22185 3927 22219
rect 3927 22185 3936 22219
rect 3884 22176 3936 22185
rect 4896 22176 4948 22228
rect 5264 22176 5316 22228
rect 5448 22176 5500 22228
rect 14004 22176 14056 22228
rect 5448 22040 5500 22092
rect 940 21972 992 22024
rect 4068 21972 4120 22024
rect 5356 22015 5408 22024
rect 5356 21981 5365 22015
rect 5365 21981 5399 22015
rect 5399 21981 5408 22015
rect 5356 21972 5408 21981
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 2688 21836 2740 21888
rect 4620 21836 4672 21888
rect 5172 21836 5224 21888
rect 5724 21972 5776 22024
rect 5908 22015 5960 22024
rect 5908 21981 5917 22015
rect 5917 21981 5951 22015
rect 5951 21981 5960 22015
rect 5908 21972 5960 21981
rect 8024 22015 8076 22024
rect 8024 21981 8033 22015
rect 8033 21981 8067 22015
rect 8067 21981 8076 22015
rect 8024 21972 8076 21981
rect 9772 22040 9824 22092
rect 9680 22015 9732 22024
rect 9680 21981 9689 22015
rect 9689 21981 9723 22015
rect 9723 21981 9732 22015
rect 9680 21972 9732 21981
rect 9312 21904 9364 21956
rect 7656 21879 7708 21888
rect 7656 21845 7665 21879
rect 7665 21845 7699 21879
rect 7699 21845 7708 21879
rect 7656 21836 7708 21845
rect 7748 21836 7800 21888
rect 8024 21836 8076 21888
rect 9496 21836 9548 21888
rect 9588 21879 9640 21888
rect 9588 21845 9597 21879
rect 9597 21845 9631 21879
rect 9631 21845 9640 21879
rect 9588 21836 9640 21845
rect 10968 22108 11020 22160
rect 14648 22108 14700 22160
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 10876 22015 10928 22024
rect 10876 21981 10885 22015
rect 10885 21981 10919 22015
rect 10919 21981 10928 22015
rect 10876 21972 10928 21981
rect 11796 22040 11848 22092
rect 11888 22015 11940 22024
rect 11888 21981 11897 22015
rect 11897 21981 11931 22015
rect 11931 21981 11940 22015
rect 11888 21972 11940 21981
rect 12532 22040 12584 22092
rect 13268 22040 13320 22092
rect 15292 22176 15344 22228
rect 20904 22176 20956 22228
rect 23388 22176 23440 22228
rect 30380 22219 30432 22228
rect 30380 22185 30389 22219
rect 30389 22185 30423 22219
rect 30423 22185 30432 22219
rect 30380 22176 30432 22185
rect 30932 22219 30984 22228
rect 30932 22185 30941 22219
rect 30941 22185 30975 22219
rect 30975 22185 30984 22219
rect 30932 22176 30984 22185
rect 34152 22176 34204 22228
rect 18052 22151 18104 22160
rect 18052 22117 18061 22151
rect 18061 22117 18095 22151
rect 18095 22117 18104 22151
rect 18052 22108 18104 22117
rect 26240 22151 26292 22160
rect 12716 21972 12768 22024
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 10140 21836 10192 21888
rect 11060 21879 11112 21888
rect 11060 21845 11069 21879
rect 11069 21845 11103 21879
rect 11103 21845 11112 21879
rect 11060 21836 11112 21845
rect 11704 21836 11756 21888
rect 11796 21836 11848 21888
rect 12624 21836 12676 21888
rect 14280 21972 14332 22024
rect 15016 21972 15068 22024
rect 17592 22083 17644 22092
rect 17592 22049 17601 22083
rect 17601 22049 17635 22083
rect 17635 22049 17644 22083
rect 17592 22040 17644 22049
rect 19340 22040 19392 22092
rect 26240 22117 26249 22151
rect 26249 22117 26283 22151
rect 26283 22117 26292 22151
rect 26240 22108 26292 22117
rect 26332 22151 26384 22160
rect 26332 22117 26341 22151
rect 26341 22117 26375 22151
rect 26375 22117 26384 22151
rect 26332 22108 26384 22117
rect 15660 21972 15712 22024
rect 17684 22015 17736 22024
rect 17684 21981 17693 22015
rect 17693 21981 17727 22015
rect 17727 21981 17736 22015
rect 17684 21972 17736 21981
rect 19524 22015 19576 22024
rect 19524 21981 19533 22015
rect 19533 21981 19567 22015
rect 19567 21981 19576 22015
rect 19524 21972 19576 21981
rect 21732 22083 21784 22092
rect 21732 22049 21741 22083
rect 21741 22049 21775 22083
rect 21775 22049 21784 22083
rect 21732 22040 21784 22049
rect 22560 22040 22612 22092
rect 26056 22040 26108 22092
rect 20076 21972 20128 22024
rect 26608 22040 26660 22092
rect 13820 21904 13872 21956
rect 14372 21947 14424 21956
rect 14372 21913 14381 21947
rect 14381 21913 14415 21947
rect 14415 21913 14424 21947
rect 14372 21904 14424 21913
rect 22192 21904 22244 21956
rect 22468 21904 22520 21956
rect 27252 22040 27304 22092
rect 27896 22108 27948 22160
rect 26884 22015 26936 22024
rect 26884 21981 26893 22015
rect 26893 21981 26927 22015
rect 26927 21981 26936 22015
rect 26884 21972 26936 21981
rect 27344 22015 27396 22024
rect 27344 21981 27353 22015
rect 27353 21981 27387 22015
rect 27387 21981 27396 22015
rect 27344 21972 27396 21981
rect 27712 21972 27764 22024
rect 27804 22015 27856 22024
rect 27804 21981 27813 22015
rect 27813 21981 27847 22015
rect 27847 21981 27856 22015
rect 27804 21972 27856 21981
rect 26792 21904 26844 21956
rect 27160 21947 27212 21956
rect 27160 21913 27169 21947
rect 27169 21913 27203 21947
rect 27203 21913 27212 21947
rect 27160 21904 27212 21913
rect 27988 21904 28040 21956
rect 14096 21836 14148 21888
rect 15292 21879 15344 21888
rect 15292 21845 15301 21879
rect 15301 21845 15335 21879
rect 15335 21845 15344 21879
rect 15292 21836 15344 21845
rect 26516 21836 26568 21888
rect 26608 21879 26660 21888
rect 26608 21845 26617 21879
rect 26617 21845 26651 21879
rect 26651 21845 26660 21879
rect 26608 21836 26660 21845
rect 26884 21836 26936 21888
rect 27528 21836 27580 21888
rect 28448 22015 28500 22024
rect 28448 21981 28457 22015
rect 28457 21981 28491 22015
rect 28491 21981 28500 22015
rect 28448 21972 28500 21981
rect 31760 22040 31812 22092
rect 29092 21904 29144 21956
rect 29920 21947 29972 21956
rect 29920 21913 29929 21947
rect 29929 21913 29963 21947
rect 29963 21913 29972 21947
rect 29920 21904 29972 21913
rect 32036 22015 32088 22024
rect 32036 21981 32045 22015
rect 32045 21981 32079 22015
rect 32079 21981 32088 22015
rect 32036 21972 32088 21981
rect 34060 21972 34112 22024
rect 32496 21904 32548 21956
rect 28816 21836 28868 21888
rect 30656 21879 30708 21888
rect 30656 21845 30665 21879
rect 30665 21845 30699 21879
rect 30699 21845 30708 21879
rect 30656 21836 30708 21845
rect 32680 21836 32732 21888
rect 34428 21836 34480 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1584 21632 1636 21684
rect 4620 21675 4672 21684
rect 4620 21641 4629 21675
rect 4629 21641 4663 21675
rect 4663 21641 4672 21675
rect 4620 21632 4672 21641
rect 4988 21607 5040 21616
rect 4988 21573 4997 21607
rect 4997 21573 5031 21607
rect 5031 21573 5040 21607
rect 4988 21564 5040 21573
rect 2688 21496 2740 21548
rect 4896 21539 4948 21548
rect 4896 21505 4905 21539
rect 4905 21505 4939 21539
rect 4939 21505 4948 21539
rect 4896 21496 4948 21505
rect 5172 21539 5224 21548
rect 5172 21505 5181 21539
rect 5181 21505 5215 21539
rect 5215 21505 5224 21539
rect 5172 21496 5224 21505
rect 5264 21539 5316 21548
rect 5264 21505 5273 21539
rect 5273 21505 5307 21539
rect 5307 21505 5316 21539
rect 5264 21496 5316 21505
rect 5356 21496 5408 21548
rect 5908 21632 5960 21684
rect 9312 21632 9364 21684
rect 10508 21632 10560 21684
rect 11796 21632 11848 21684
rect 11888 21632 11940 21684
rect 12072 21632 12124 21684
rect 12164 21675 12216 21684
rect 12164 21641 12173 21675
rect 12173 21641 12207 21675
rect 12207 21641 12216 21675
rect 12164 21632 12216 21641
rect 12716 21632 12768 21684
rect 13820 21632 13872 21684
rect 14464 21632 14516 21684
rect 14648 21675 14700 21684
rect 14648 21641 14657 21675
rect 14657 21641 14691 21675
rect 14691 21641 14700 21675
rect 14648 21632 14700 21641
rect 17592 21632 17644 21684
rect 19248 21632 19300 21684
rect 21732 21632 21784 21684
rect 5816 21564 5868 21616
rect 5724 21496 5776 21548
rect 8024 21564 8076 21616
rect 1400 21428 1452 21480
rect 2596 21428 2648 21480
rect 3148 21428 3200 21480
rect 5080 21360 5132 21412
rect 8852 21539 8904 21548
rect 8852 21505 8861 21539
rect 8861 21505 8895 21539
rect 8895 21505 8904 21539
rect 8852 21496 8904 21505
rect 6460 21428 6512 21480
rect 6828 21428 6880 21480
rect 6368 21360 6420 21412
rect 6644 21360 6696 21412
rect 10232 21496 10284 21548
rect 9496 21471 9548 21480
rect 9496 21437 9505 21471
rect 9505 21437 9539 21471
rect 9539 21437 9548 21471
rect 9496 21428 9548 21437
rect 10324 21428 10376 21480
rect 11060 21496 11112 21548
rect 13636 21564 13688 21616
rect 14004 21564 14056 21616
rect 11980 21539 12032 21548
rect 11980 21505 11989 21539
rect 11989 21505 12023 21539
rect 12023 21505 12032 21539
rect 11980 21496 12032 21505
rect 13084 21496 13136 21548
rect 15016 21496 15068 21548
rect 15292 21496 15344 21548
rect 12532 21428 12584 21480
rect 14648 21428 14700 21480
rect 12808 21360 12860 21412
rect 2228 21335 2280 21344
rect 2228 21301 2237 21335
rect 2237 21301 2271 21335
rect 2271 21301 2280 21335
rect 2228 21292 2280 21301
rect 2688 21335 2740 21344
rect 2688 21301 2697 21335
rect 2697 21301 2731 21335
rect 2731 21301 2740 21335
rect 2688 21292 2740 21301
rect 2872 21292 2924 21344
rect 4988 21292 5040 21344
rect 6552 21292 6604 21344
rect 6736 21335 6788 21344
rect 6736 21301 6745 21335
rect 6745 21301 6779 21335
rect 6779 21301 6788 21335
rect 6736 21292 6788 21301
rect 10968 21292 11020 21344
rect 11980 21292 12032 21344
rect 12900 21292 12952 21344
rect 15660 21539 15712 21548
rect 15660 21505 15669 21539
rect 15669 21505 15703 21539
rect 15703 21505 15712 21539
rect 15660 21496 15712 21505
rect 16672 21496 16724 21548
rect 16948 21471 17000 21480
rect 16948 21437 16957 21471
rect 16957 21437 16991 21471
rect 16991 21437 17000 21471
rect 16948 21428 17000 21437
rect 20628 21496 20680 21548
rect 19432 21471 19484 21480
rect 19432 21437 19441 21471
rect 19441 21437 19475 21471
rect 19475 21437 19484 21471
rect 19432 21428 19484 21437
rect 22560 21632 22612 21684
rect 23572 21632 23624 21684
rect 26792 21675 26844 21684
rect 26792 21641 26801 21675
rect 26801 21641 26835 21675
rect 26835 21641 26844 21675
rect 26792 21632 26844 21641
rect 27160 21675 27212 21684
rect 27160 21641 27169 21675
rect 27169 21641 27203 21675
rect 27203 21641 27212 21675
rect 27160 21632 27212 21641
rect 22836 21564 22888 21616
rect 19708 21403 19760 21412
rect 19708 21369 19717 21403
rect 19717 21369 19751 21403
rect 19751 21369 19760 21403
rect 19708 21360 19760 21369
rect 26332 21471 26384 21480
rect 26332 21437 26341 21471
rect 26341 21437 26375 21471
rect 26375 21437 26384 21471
rect 26332 21428 26384 21437
rect 26608 21564 26660 21616
rect 27712 21632 27764 21684
rect 27896 21632 27948 21684
rect 29092 21675 29144 21684
rect 29092 21641 29101 21675
rect 29101 21641 29135 21675
rect 29135 21641 29144 21675
rect 29092 21632 29144 21641
rect 29920 21632 29972 21684
rect 28724 21607 28776 21616
rect 28724 21573 28733 21607
rect 28733 21573 28767 21607
rect 28767 21573 28776 21607
rect 28724 21564 28776 21573
rect 28816 21564 28868 21616
rect 26516 21539 26568 21548
rect 26516 21505 26525 21539
rect 26525 21505 26559 21539
rect 26559 21505 26568 21539
rect 26516 21496 26568 21505
rect 26792 21496 26844 21548
rect 27528 21496 27580 21548
rect 27804 21496 27856 21548
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 26700 21360 26752 21412
rect 29000 21428 29052 21480
rect 20720 21292 20772 21344
rect 21824 21292 21876 21344
rect 23112 21292 23164 21344
rect 23296 21292 23348 21344
rect 26424 21292 26476 21344
rect 27528 21335 27580 21344
rect 27528 21301 27537 21335
rect 27537 21301 27571 21335
rect 27571 21301 27580 21335
rect 27528 21292 27580 21301
rect 27620 21335 27672 21344
rect 27620 21301 27629 21335
rect 27629 21301 27663 21335
rect 27663 21301 27672 21335
rect 27620 21292 27672 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3148 21088 3200 21140
rect 4896 21088 4948 21140
rect 5356 21088 5408 21140
rect 6644 21131 6696 21140
rect 6644 21097 6653 21131
rect 6653 21097 6687 21131
rect 6687 21097 6696 21131
rect 6644 21088 6696 21097
rect 6736 21088 6788 21140
rect 8852 21088 8904 21140
rect 10324 21088 10376 21140
rect 1676 20995 1728 21004
rect 1676 20961 1685 20995
rect 1685 20961 1719 20995
rect 1719 20961 1728 20995
rect 1676 20952 1728 20961
rect 4804 20952 4856 21004
rect 6368 20952 6420 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 6552 20884 6604 20936
rect 6736 20927 6788 20936
rect 6736 20893 6745 20927
rect 6745 20893 6779 20927
rect 6779 20893 6788 20927
rect 6736 20884 6788 20893
rect 10876 21088 10928 21140
rect 11888 21088 11940 21140
rect 11980 21131 12032 21140
rect 11980 21097 11989 21131
rect 11989 21097 12023 21131
rect 12023 21097 12032 21131
rect 11980 21088 12032 21097
rect 12440 21088 12492 21140
rect 12624 21088 12676 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 10968 20952 11020 21004
rect 11336 20884 11388 20936
rect 12716 20952 12768 21004
rect 12900 20995 12952 21004
rect 12900 20961 12909 20995
rect 12909 20961 12943 20995
rect 12943 20961 12952 20995
rect 13912 21088 13964 21140
rect 12900 20952 12952 20961
rect 2228 20816 2280 20868
rect 7748 20816 7800 20868
rect 11888 20927 11940 20936
rect 11888 20893 11897 20927
rect 11897 20893 11931 20927
rect 11931 20893 11940 20927
rect 11888 20884 11940 20893
rect 13268 20927 13320 20936
rect 13268 20893 13277 20927
rect 13277 20893 13311 20927
rect 13311 20893 13320 20927
rect 13268 20884 13320 20893
rect 13636 20995 13688 21004
rect 13636 20961 13645 20995
rect 13645 20961 13679 20995
rect 13679 20961 13688 20995
rect 13636 20952 13688 20961
rect 13820 20952 13872 21004
rect 5264 20748 5316 20800
rect 6736 20748 6788 20800
rect 8944 20748 8996 20800
rect 11980 20816 12032 20868
rect 12256 20816 12308 20868
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 14372 20816 14424 20868
rect 17132 20927 17184 20936
rect 17132 20893 17141 20927
rect 17141 20893 17175 20927
rect 17175 20893 17184 20927
rect 17132 20884 17184 20893
rect 17868 21020 17920 21072
rect 17592 20884 17644 20936
rect 11796 20748 11848 20800
rect 12532 20791 12584 20800
rect 12532 20757 12541 20791
rect 12541 20757 12575 20791
rect 12575 20757 12584 20791
rect 12532 20748 12584 20757
rect 13820 20748 13872 20800
rect 16948 20748 17000 20800
rect 17868 20748 17920 20800
rect 19708 20884 19760 20936
rect 20444 21088 20496 21140
rect 21824 21131 21876 21140
rect 21824 21097 21833 21131
rect 21833 21097 21867 21131
rect 21867 21097 21876 21131
rect 21824 21088 21876 21097
rect 20076 21063 20128 21072
rect 20076 21029 20085 21063
rect 20085 21029 20119 21063
rect 20119 21029 20128 21063
rect 20076 21020 20128 21029
rect 20260 20884 20312 20936
rect 22560 20929 22612 20936
rect 22560 20895 22577 20929
rect 22577 20895 22611 20929
rect 22611 20895 22612 20929
rect 23112 20952 23164 21004
rect 23572 21131 23624 21140
rect 23572 21097 23581 21131
rect 23581 21097 23615 21131
rect 23615 21097 23624 21131
rect 23572 21088 23624 21097
rect 24032 21088 24084 21140
rect 24952 21088 25004 21140
rect 26332 21088 26384 21140
rect 26700 21131 26752 21140
rect 26700 21097 26709 21131
rect 26709 21097 26743 21131
rect 26743 21097 26752 21131
rect 26700 21088 26752 21097
rect 27620 21088 27672 21140
rect 22560 20884 22612 20895
rect 22836 20927 22888 20936
rect 22836 20893 22845 20927
rect 22845 20893 22879 20927
rect 22879 20893 22888 20927
rect 22836 20884 22888 20893
rect 18328 20791 18380 20800
rect 18328 20757 18337 20791
rect 18337 20757 18371 20791
rect 18371 20757 18380 20791
rect 18328 20748 18380 20757
rect 20168 20748 20220 20800
rect 22928 20816 22980 20868
rect 23204 20884 23256 20936
rect 23480 20952 23532 21004
rect 25320 21020 25372 21072
rect 24492 20995 24544 21004
rect 24492 20961 24501 20995
rect 24501 20961 24535 20995
rect 24535 20961 24544 20995
rect 24492 20952 24544 20961
rect 23664 20927 23716 20936
rect 23664 20893 23673 20927
rect 23673 20893 23707 20927
rect 23707 20893 23716 20927
rect 23664 20884 23716 20893
rect 23848 20927 23900 20936
rect 23848 20893 23857 20927
rect 23857 20893 23891 20927
rect 23891 20893 23900 20927
rect 23848 20884 23900 20893
rect 23756 20816 23808 20868
rect 24124 20884 24176 20936
rect 24860 20884 24912 20936
rect 25780 20927 25832 20936
rect 25780 20893 25789 20927
rect 25789 20893 25823 20927
rect 25823 20893 25832 20927
rect 25780 20884 25832 20893
rect 25872 20927 25924 20936
rect 25872 20893 25881 20927
rect 25881 20893 25915 20927
rect 25915 20893 25924 20927
rect 25872 20884 25924 20893
rect 34520 20927 34572 20936
rect 34520 20893 34529 20927
rect 34529 20893 34563 20927
rect 34563 20893 34572 20927
rect 34520 20884 34572 20893
rect 34060 20816 34112 20868
rect 25504 20791 25556 20800
rect 25504 20757 25513 20791
rect 25513 20757 25547 20791
rect 25547 20757 25556 20791
rect 25504 20748 25556 20757
rect 25872 20748 25924 20800
rect 26424 20748 26476 20800
rect 27896 20748 27948 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 9496 20544 9548 20596
rect 11704 20544 11756 20596
rect 13912 20587 13964 20596
rect 13912 20553 13921 20587
rect 13921 20553 13955 20587
rect 13955 20553 13964 20587
rect 13912 20544 13964 20553
rect 14188 20544 14240 20596
rect 10692 20476 10744 20528
rect 11520 20476 11572 20528
rect 11796 20519 11848 20528
rect 11796 20485 11805 20519
rect 11805 20485 11839 20519
rect 11839 20485 11848 20519
rect 11796 20476 11848 20485
rect 13268 20476 13320 20528
rect 14372 20519 14424 20528
rect 14372 20485 14381 20519
rect 14381 20485 14415 20519
rect 14415 20485 14424 20519
rect 14372 20476 14424 20485
rect 15108 20476 15160 20528
rect 16856 20519 16908 20528
rect 16856 20485 16865 20519
rect 16865 20485 16899 20519
rect 16899 20485 16908 20519
rect 16856 20476 16908 20485
rect 17132 20544 17184 20596
rect 17684 20544 17736 20596
rect 22560 20544 22612 20596
rect 22744 20544 22796 20596
rect 22836 20544 22888 20596
rect 23480 20544 23532 20596
rect 11060 20408 11112 20460
rect 12072 20451 12124 20460
rect 12072 20417 12081 20451
rect 12081 20417 12115 20451
rect 12115 20417 12124 20451
rect 12072 20408 12124 20417
rect 12256 20451 12308 20460
rect 12256 20417 12265 20451
rect 12265 20417 12299 20451
rect 12299 20417 12308 20451
rect 12256 20408 12308 20417
rect 12532 20451 12584 20460
rect 12532 20417 12541 20451
rect 12541 20417 12575 20451
rect 12575 20417 12584 20451
rect 12532 20408 12584 20417
rect 13176 20451 13228 20460
rect 13176 20417 13185 20451
rect 13185 20417 13219 20451
rect 13219 20417 13228 20451
rect 13176 20408 13228 20417
rect 13912 20408 13964 20460
rect 14188 20408 14240 20460
rect 14280 20451 14332 20460
rect 14280 20417 14289 20451
rect 14289 20417 14323 20451
rect 14323 20417 14332 20451
rect 14280 20408 14332 20417
rect 14464 20451 14516 20460
rect 14464 20417 14473 20451
rect 14473 20417 14507 20451
rect 14507 20417 14516 20451
rect 14464 20408 14516 20417
rect 15476 20408 15528 20460
rect 16948 20408 17000 20460
rect 24492 20587 24544 20596
rect 24492 20553 24501 20587
rect 24501 20553 24535 20587
rect 24535 20553 24544 20587
rect 24492 20544 24544 20553
rect 25320 20587 25372 20596
rect 25320 20553 25329 20587
rect 25329 20553 25363 20587
rect 25363 20553 25372 20587
rect 25320 20544 25372 20553
rect 23848 20476 23900 20528
rect 12164 20340 12216 20392
rect 2320 20247 2372 20256
rect 2320 20213 2329 20247
rect 2329 20213 2363 20247
rect 2363 20213 2372 20247
rect 2320 20204 2372 20213
rect 2872 20204 2924 20256
rect 3056 20204 3108 20256
rect 8944 20204 8996 20256
rect 9496 20204 9548 20256
rect 10232 20247 10284 20256
rect 10232 20213 10241 20247
rect 10241 20213 10275 20247
rect 10275 20213 10284 20247
rect 10232 20204 10284 20213
rect 10508 20204 10560 20256
rect 11244 20204 11296 20256
rect 12716 20247 12768 20256
rect 12716 20213 12725 20247
rect 12725 20213 12759 20247
rect 12759 20213 12768 20247
rect 12716 20204 12768 20213
rect 15384 20383 15436 20392
rect 15384 20349 15393 20383
rect 15393 20349 15427 20383
rect 15427 20349 15436 20383
rect 15384 20340 15436 20349
rect 16672 20340 16724 20392
rect 23664 20408 23716 20460
rect 20444 20383 20496 20392
rect 20444 20349 20453 20383
rect 20453 20349 20487 20383
rect 20487 20349 20496 20383
rect 20444 20340 20496 20349
rect 23756 20340 23808 20392
rect 28724 20544 28776 20596
rect 13636 20272 13688 20324
rect 17408 20272 17460 20324
rect 20168 20272 20220 20324
rect 14188 20247 14240 20256
rect 14188 20213 14197 20247
rect 14197 20213 14231 20247
rect 14231 20213 14240 20247
rect 14188 20204 14240 20213
rect 14924 20204 14976 20256
rect 17776 20204 17828 20256
rect 20260 20247 20312 20256
rect 20260 20213 20269 20247
rect 20269 20213 20303 20247
rect 20303 20213 20312 20247
rect 20260 20204 20312 20213
rect 22836 20247 22888 20256
rect 22836 20213 22845 20247
rect 22845 20213 22879 20247
rect 22879 20213 22888 20247
rect 22836 20204 22888 20213
rect 23572 20272 23624 20324
rect 25780 20408 25832 20460
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 28172 20408 28224 20460
rect 24860 20204 24912 20256
rect 25596 20204 25648 20256
rect 27620 20340 27672 20392
rect 28172 20247 28224 20256
rect 28172 20213 28181 20247
rect 28181 20213 28215 20247
rect 28215 20213 28224 20247
rect 28172 20204 28224 20213
rect 28448 20204 28500 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4712 20000 4764 20052
rect 10692 20043 10744 20052
rect 10692 20009 10701 20043
rect 10701 20009 10735 20043
rect 10735 20009 10744 20043
rect 10692 20000 10744 20009
rect 11060 20043 11112 20052
rect 11060 20009 11069 20043
rect 11069 20009 11103 20043
rect 11103 20009 11112 20043
rect 11060 20000 11112 20009
rect 11336 20000 11388 20052
rect 2044 19907 2096 19916
rect 2044 19873 2053 19907
rect 2053 19873 2087 19907
rect 2087 19873 2096 19907
rect 2044 19864 2096 19873
rect 940 19796 992 19848
rect 3056 19796 3108 19848
rect 4436 19932 4488 19984
rect 4252 19907 4304 19916
rect 4252 19873 4261 19907
rect 4261 19873 4295 19907
rect 4295 19873 4304 19907
rect 4252 19864 4304 19873
rect 4988 19907 5040 19916
rect 4988 19873 4997 19907
rect 4997 19873 5031 19907
rect 5031 19873 5040 19907
rect 4988 19864 5040 19873
rect 5448 19864 5500 19916
rect 8944 19864 8996 19916
rect 11980 20000 12032 20052
rect 11980 19864 12032 19916
rect 12164 19907 12216 19916
rect 12164 19873 12173 19907
rect 12173 19873 12207 19907
rect 12207 19873 12216 19907
rect 12164 19864 12216 19873
rect 12256 19864 12308 19916
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 5264 19839 5316 19848
rect 5264 19805 5273 19839
rect 5273 19805 5307 19839
rect 5307 19805 5316 19839
rect 5264 19796 5316 19805
rect 7656 19796 7708 19848
rect 1400 19660 1452 19712
rect 1676 19660 1728 19712
rect 4160 19660 4212 19712
rect 4896 19660 4948 19712
rect 4988 19703 5040 19712
rect 4988 19669 4997 19703
rect 4997 19669 5031 19703
rect 5031 19669 5040 19703
rect 4988 19660 5040 19669
rect 7564 19660 7616 19712
rect 8576 19839 8628 19848
rect 8576 19805 8585 19839
rect 8585 19805 8619 19839
rect 8619 19805 8628 19839
rect 8576 19796 8628 19805
rect 9496 19796 9548 19848
rect 11244 19839 11296 19848
rect 11244 19805 11253 19839
rect 11253 19805 11287 19839
rect 11287 19805 11296 19839
rect 11244 19796 11296 19805
rect 11520 19796 11572 19848
rect 11796 19839 11848 19848
rect 11796 19805 11805 19839
rect 11805 19805 11839 19839
rect 11839 19805 11848 19839
rect 12716 20000 12768 20052
rect 13176 20043 13228 20052
rect 13176 20009 13185 20043
rect 13185 20009 13219 20043
rect 13219 20009 13228 20043
rect 13176 20000 13228 20009
rect 13360 20043 13412 20052
rect 13360 20009 13369 20043
rect 13369 20009 13403 20043
rect 13403 20009 13412 20043
rect 13360 20000 13412 20009
rect 14188 20000 14240 20052
rect 15384 20000 15436 20052
rect 15476 20000 15528 20052
rect 16856 20000 16908 20052
rect 16948 20000 17000 20052
rect 17684 20000 17736 20052
rect 17868 20043 17920 20052
rect 17868 20009 17877 20043
rect 17877 20009 17911 20043
rect 17911 20009 17920 20043
rect 17868 20000 17920 20009
rect 17960 20000 18012 20052
rect 20996 20000 21048 20052
rect 22468 20000 22520 20052
rect 11796 19796 11848 19805
rect 12440 19839 12492 19848
rect 12440 19805 12449 19839
rect 12449 19805 12483 19839
rect 12483 19805 12492 19839
rect 12440 19796 12492 19805
rect 14096 19864 14148 19916
rect 13820 19839 13872 19848
rect 13820 19805 13829 19839
rect 13829 19805 13863 19839
rect 13863 19805 13872 19839
rect 13820 19796 13872 19805
rect 15108 19907 15160 19916
rect 15108 19873 15117 19907
rect 15117 19873 15151 19907
rect 15151 19873 15160 19907
rect 15108 19864 15160 19873
rect 15384 19839 15436 19848
rect 15384 19805 15393 19839
rect 15393 19805 15427 19839
rect 15427 19805 15436 19839
rect 15384 19796 15436 19805
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 15660 19796 15712 19805
rect 16120 19796 16172 19848
rect 16856 19864 16908 19916
rect 18788 19932 18840 19984
rect 9036 19771 9088 19780
rect 9036 19737 9045 19771
rect 9045 19737 9079 19771
rect 9079 19737 9088 19771
rect 9036 19728 9088 19737
rect 12256 19728 12308 19780
rect 13452 19728 13504 19780
rect 14924 19728 14976 19780
rect 8484 19660 8536 19712
rect 8760 19703 8812 19712
rect 8760 19669 8769 19703
rect 8769 19669 8803 19703
rect 8803 19669 8812 19703
rect 8760 19660 8812 19669
rect 10140 19703 10192 19712
rect 10140 19669 10149 19703
rect 10149 19669 10183 19703
rect 10183 19669 10192 19703
rect 10140 19660 10192 19669
rect 12164 19660 12216 19712
rect 14464 19660 14516 19712
rect 15384 19660 15436 19712
rect 16212 19660 16264 19712
rect 19064 19864 19116 19916
rect 17684 19839 17736 19848
rect 17684 19805 17693 19839
rect 17693 19805 17727 19839
rect 17727 19805 17736 19839
rect 17684 19796 17736 19805
rect 17776 19839 17828 19848
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 19340 19796 19392 19848
rect 20260 19907 20312 19916
rect 20260 19873 20269 19907
rect 20269 19873 20303 19907
rect 20303 19873 20312 19907
rect 20260 19864 20312 19873
rect 20812 19864 20864 19916
rect 24124 20000 24176 20052
rect 22928 19864 22980 19916
rect 17960 19771 18012 19780
rect 17960 19737 17969 19771
rect 17969 19737 18003 19771
rect 18003 19737 18012 19771
rect 17960 19728 18012 19737
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 20904 19796 20956 19848
rect 21916 19796 21968 19848
rect 22744 19796 22796 19848
rect 21088 19728 21140 19780
rect 23664 19796 23716 19848
rect 25504 19864 25556 19916
rect 23296 19728 23348 19780
rect 19432 19660 19484 19712
rect 19984 19660 20036 19712
rect 22100 19660 22152 19712
rect 22836 19660 22888 19712
rect 25596 19839 25648 19848
rect 25596 19805 25605 19839
rect 25605 19805 25639 19839
rect 25639 19805 25648 19839
rect 25596 19796 25648 19805
rect 25780 19796 25832 19848
rect 26056 19932 26108 19984
rect 28172 20000 28224 20052
rect 34520 20043 34572 20052
rect 34520 20009 34529 20043
rect 34529 20009 34563 20043
rect 34563 20009 34572 20043
rect 34520 20000 34572 20009
rect 27528 19864 27580 19916
rect 27804 19796 27856 19848
rect 29644 19864 29696 19916
rect 32680 19932 32732 19984
rect 28448 19796 28500 19848
rect 31852 19907 31904 19916
rect 31852 19873 31861 19907
rect 31861 19873 31895 19907
rect 31895 19873 31904 19907
rect 31852 19864 31904 19873
rect 32128 19796 32180 19848
rect 34520 19796 34572 19848
rect 26608 19728 26660 19780
rect 27620 19728 27672 19780
rect 27896 19771 27948 19780
rect 27896 19737 27905 19771
rect 27905 19737 27939 19771
rect 27939 19737 27948 19771
rect 27896 19728 27948 19737
rect 27804 19660 27856 19712
rect 30748 19728 30800 19780
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4252 19499 4304 19508
rect 4252 19465 4261 19499
rect 4261 19465 4295 19499
rect 4295 19465 4304 19499
rect 4252 19456 4304 19465
rect 4712 19499 4764 19508
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 5172 19456 5224 19508
rect 8576 19456 8628 19508
rect 11796 19499 11848 19508
rect 11796 19465 11805 19499
rect 11805 19465 11839 19499
rect 11839 19465 11848 19499
rect 11796 19456 11848 19465
rect 12072 19456 12124 19508
rect 12808 19499 12860 19508
rect 12808 19465 12817 19499
rect 12817 19465 12851 19499
rect 12851 19465 12860 19499
rect 12808 19456 12860 19465
rect 13452 19456 13504 19508
rect 15660 19456 15712 19508
rect 16212 19456 16264 19508
rect 17960 19456 18012 19508
rect 2320 19388 2372 19440
rect 1400 19363 1452 19372
rect 1400 19329 1409 19363
rect 1409 19329 1443 19363
rect 1443 19329 1452 19363
rect 1400 19320 1452 19329
rect 4160 19388 4212 19440
rect 1768 19252 1820 19304
rect 4988 19388 5040 19440
rect 6736 19388 6788 19440
rect 8760 19388 8812 19440
rect 10140 19388 10192 19440
rect 11244 19431 11296 19440
rect 11244 19397 11253 19431
rect 11253 19397 11287 19431
rect 11287 19397 11296 19431
rect 11244 19388 11296 19397
rect 11980 19388 12032 19440
rect 12532 19388 12584 19440
rect 16396 19431 16448 19440
rect 16396 19397 16405 19431
rect 16405 19397 16439 19431
rect 16439 19397 16448 19431
rect 16396 19388 16448 19397
rect 17684 19388 17736 19440
rect 18788 19456 18840 19508
rect 19064 19388 19116 19440
rect 5264 19320 5316 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 11520 19320 11572 19372
rect 17868 19320 17920 19372
rect 20168 19499 20220 19508
rect 20168 19465 20177 19499
rect 20177 19465 20211 19499
rect 20211 19465 20220 19499
rect 20168 19456 20220 19465
rect 20628 19456 20680 19508
rect 21548 19456 21600 19508
rect 4804 19252 4856 19304
rect 5172 19252 5224 19304
rect 5632 19295 5684 19304
rect 5632 19261 5641 19295
rect 5641 19261 5675 19295
rect 5675 19261 5684 19295
rect 5632 19252 5684 19261
rect 8484 19252 8536 19304
rect 14648 19252 14700 19304
rect 15384 19252 15436 19304
rect 18052 19252 18104 19304
rect 18328 19252 18380 19304
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 17684 19227 17736 19236
rect 17684 19193 17693 19227
rect 17693 19193 17727 19227
rect 17727 19193 17736 19227
rect 17684 19184 17736 19193
rect 3056 19116 3108 19168
rect 3424 19116 3476 19168
rect 3976 19116 4028 19168
rect 4436 19159 4488 19168
rect 4436 19125 4445 19159
rect 4445 19125 4479 19159
rect 4479 19125 4488 19159
rect 4436 19116 4488 19125
rect 4988 19116 5040 19168
rect 5264 19116 5316 19168
rect 5448 19116 5500 19168
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 8944 19116 8996 19168
rect 18328 19116 18380 19168
rect 18696 19252 18748 19304
rect 19340 19320 19392 19372
rect 19616 19320 19668 19372
rect 20720 19388 20772 19440
rect 19984 19320 20036 19372
rect 20904 19320 20956 19372
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 21640 19363 21692 19372
rect 21640 19329 21649 19363
rect 21649 19329 21683 19363
rect 21683 19329 21692 19363
rect 21640 19320 21692 19329
rect 22744 19456 22796 19508
rect 23480 19456 23532 19508
rect 25964 19456 26016 19508
rect 29644 19499 29696 19508
rect 29644 19465 29653 19499
rect 29653 19465 29687 19499
rect 29687 19465 29696 19499
rect 29644 19456 29696 19465
rect 30748 19499 30800 19508
rect 30748 19465 30757 19499
rect 30757 19465 30791 19499
rect 30791 19465 30800 19499
rect 30748 19456 30800 19465
rect 31852 19456 31904 19508
rect 32496 19499 32548 19508
rect 32496 19465 32505 19499
rect 32505 19465 32539 19499
rect 32539 19465 32548 19499
rect 32496 19456 32548 19465
rect 26424 19388 26476 19440
rect 19064 19227 19116 19236
rect 19064 19193 19073 19227
rect 19073 19193 19107 19227
rect 19107 19193 19116 19227
rect 19064 19184 19116 19193
rect 22100 19252 22152 19304
rect 22928 19320 22980 19372
rect 26700 19320 26752 19372
rect 30656 19363 30708 19372
rect 25596 19295 25648 19304
rect 25596 19261 25605 19295
rect 25605 19261 25639 19295
rect 25639 19261 25648 19295
rect 25596 19252 25648 19261
rect 21732 19116 21784 19168
rect 24584 19184 24636 19236
rect 22192 19159 22244 19168
rect 22192 19125 22201 19159
rect 22201 19125 22235 19159
rect 22235 19125 22244 19159
rect 22192 19116 22244 19125
rect 22560 19159 22612 19168
rect 22560 19125 22569 19159
rect 22569 19125 22603 19159
rect 22603 19125 22612 19159
rect 22560 19116 22612 19125
rect 24676 19116 24728 19168
rect 25780 19159 25832 19168
rect 25780 19125 25789 19159
rect 25789 19125 25823 19159
rect 25823 19125 25832 19159
rect 25780 19116 25832 19125
rect 30196 19116 30248 19168
rect 30656 19329 30665 19363
rect 30665 19329 30699 19363
rect 30699 19329 30708 19363
rect 30656 19320 30708 19329
rect 31668 19363 31720 19372
rect 31668 19329 31677 19363
rect 31677 19329 31711 19363
rect 31711 19329 31720 19363
rect 31668 19320 31720 19329
rect 31944 19295 31996 19304
rect 31944 19261 31953 19295
rect 31953 19261 31987 19295
rect 31987 19261 31996 19295
rect 31944 19252 31996 19261
rect 32404 19320 32456 19372
rect 32128 19159 32180 19168
rect 32128 19125 32137 19159
rect 32137 19125 32171 19159
rect 32171 19125 32180 19159
rect 32128 19116 32180 19125
rect 34336 19116 34388 19168
rect 34520 19159 34572 19168
rect 34520 19125 34529 19159
rect 34529 19125 34563 19159
rect 34563 19125 34572 19159
rect 34520 19116 34572 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4712 18912 4764 18964
rect 4896 18912 4948 18964
rect 5632 18912 5684 18964
rect 9036 18912 9088 18964
rect 3976 18776 4028 18828
rect 10232 18912 10284 18964
rect 13452 18912 13504 18964
rect 14556 18912 14608 18964
rect 19616 18912 19668 18964
rect 22192 18912 22244 18964
rect 25780 18912 25832 18964
rect 26700 18955 26752 18964
rect 26700 18921 26709 18955
rect 26709 18921 26743 18955
rect 26743 18921 26752 18955
rect 26700 18912 26752 18921
rect 27896 18912 27948 18964
rect 9772 18844 9824 18896
rect 3056 18615 3108 18624
rect 3056 18581 3065 18615
rect 3065 18581 3099 18615
rect 3099 18581 3108 18615
rect 3056 18572 3108 18581
rect 3424 18751 3476 18760
rect 3424 18717 3433 18751
rect 3433 18717 3467 18751
rect 3467 18717 3476 18751
rect 10692 18776 10744 18828
rect 11244 18776 11296 18828
rect 3424 18708 3476 18717
rect 6552 18751 6604 18760
rect 6552 18717 6561 18751
rect 6561 18717 6595 18751
rect 6595 18717 6604 18751
rect 6552 18708 6604 18717
rect 8300 18708 8352 18760
rect 10416 18708 10468 18760
rect 7564 18640 7616 18692
rect 10876 18640 10928 18692
rect 4896 18572 4948 18624
rect 5172 18572 5224 18624
rect 5448 18572 5500 18624
rect 8484 18572 8536 18624
rect 9588 18572 9640 18624
rect 11060 18572 11112 18624
rect 11612 18751 11664 18760
rect 11612 18717 11621 18751
rect 11621 18717 11655 18751
rect 11655 18717 11664 18751
rect 11612 18708 11664 18717
rect 11796 18640 11848 18692
rect 15108 18708 15160 18760
rect 17224 18751 17276 18760
rect 17224 18717 17233 18751
rect 17233 18717 17267 18751
rect 17267 18717 17276 18751
rect 17224 18708 17276 18717
rect 17316 18751 17368 18760
rect 17316 18717 17325 18751
rect 17325 18717 17359 18751
rect 17359 18717 17368 18751
rect 17316 18708 17368 18717
rect 18604 18844 18656 18896
rect 18972 18844 19024 18896
rect 21916 18887 21968 18896
rect 21916 18853 21925 18887
rect 21925 18853 21959 18887
rect 21959 18853 21968 18887
rect 21916 18844 21968 18853
rect 19340 18776 19392 18828
rect 22560 18776 22612 18828
rect 27620 18844 27672 18896
rect 25688 18776 25740 18828
rect 18512 18751 18564 18760
rect 14004 18640 14056 18692
rect 16120 18640 16172 18692
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 19064 18708 19116 18760
rect 20904 18751 20956 18760
rect 20904 18717 20913 18751
rect 20913 18717 20947 18751
rect 20947 18717 20956 18751
rect 20904 18708 20956 18717
rect 13176 18572 13228 18624
rect 13268 18572 13320 18624
rect 16212 18572 16264 18624
rect 17224 18572 17276 18624
rect 20720 18640 20772 18692
rect 21088 18640 21140 18692
rect 21364 18708 21416 18760
rect 21824 18708 21876 18760
rect 22468 18708 22520 18760
rect 21548 18640 21600 18692
rect 23204 18708 23256 18760
rect 23848 18572 23900 18624
rect 24492 18751 24544 18760
rect 24492 18717 24501 18751
rect 24501 18717 24535 18751
rect 24535 18717 24544 18751
rect 24492 18708 24544 18717
rect 24676 18751 24728 18760
rect 24676 18717 24685 18751
rect 24685 18717 24719 18751
rect 24719 18717 24728 18751
rect 24676 18708 24728 18717
rect 26148 18776 26200 18828
rect 31944 18844 31996 18896
rect 25872 18640 25924 18692
rect 25412 18572 25464 18624
rect 25596 18615 25648 18624
rect 25596 18581 25605 18615
rect 25605 18581 25639 18615
rect 25639 18581 25648 18615
rect 25596 18572 25648 18581
rect 25688 18615 25740 18624
rect 25688 18581 25697 18615
rect 25697 18581 25731 18615
rect 25731 18581 25740 18615
rect 25688 18572 25740 18581
rect 26240 18751 26292 18760
rect 26240 18717 26249 18751
rect 26249 18717 26283 18751
rect 26283 18717 26292 18751
rect 26240 18708 26292 18717
rect 31668 18776 31720 18828
rect 26792 18708 26844 18760
rect 27804 18708 27856 18760
rect 29552 18751 29604 18760
rect 29552 18717 29561 18751
rect 29561 18717 29595 18751
rect 29595 18717 29604 18751
rect 29552 18708 29604 18717
rect 32680 18776 32732 18828
rect 33048 18776 33100 18828
rect 32404 18751 32456 18760
rect 32404 18717 32413 18751
rect 32413 18717 32447 18751
rect 32447 18717 32456 18751
rect 32404 18708 32456 18717
rect 32588 18751 32640 18760
rect 32588 18717 32597 18751
rect 32597 18717 32631 18751
rect 32631 18717 32640 18751
rect 32588 18708 32640 18717
rect 34336 18708 34388 18760
rect 30288 18640 30340 18692
rect 34520 18615 34572 18624
rect 34520 18581 34529 18615
rect 34529 18581 34563 18615
rect 34563 18581 34572 18615
rect 34520 18572 34572 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 12532 18300 12584 18352
rect 14004 18343 14056 18352
rect 14004 18309 14013 18343
rect 14013 18309 14047 18343
rect 14047 18309 14056 18343
rect 14004 18300 14056 18309
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 4988 18232 5040 18284
rect 5448 18275 5500 18284
rect 5448 18241 5457 18275
rect 5457 18241 5491 18275
rect 5491 18241 5500 18275
rect 5448 18232 5500 18241
rect 10692 18232 10744 18284
rect 8300 18096 8352 18148
rect 10876 18139 10928 18148
rect 10876 18105 10885 18139
rect 10885 18105 10919 18139
rect 10919 18105 10928 18139
rect 11336 18275 11388 18284
rect 11336 18241 11345 18275
rect 11345 18241 11379 18275
rect 11379 18241 11388 18275
rect 11336 18232 11388 18241
rect 12808 18275 12860 18284
rect 12808 18241 12817 18275
rect 12817 18241 12851 18275
rect 12851 18241 12860 18275
rect 12808 18232 12860 18241
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 13084 18275 13136 18284
rect 13084 18241 13093 18275
rect 13093 18241 13127 18275
rect 13127 18241 13136 18275
rect 13084 18232 13136 18241
rect 13268 18275 13320 18284
rect 13268 18241 13277 18275
rect 13277 18241 13311 18275
rect 13311 18241 13320 18275
rect 13268 18232 13320 18241
rect 13452 18232 13504 18284
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 11796 18207 11848 18216
rect 11796 18173 11805 18207
rect 11805 18173 11839 18207
rect 11839 18173 11848 18207
rect 11796 18164 11848 18173
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 17316 18300 17368 18352
rect 17592 18368 17644 18420
rect 21732 18368 21784 18420
rect 23388 18411 23440 18420
rect 23388 18377 23397 18411
rect 23397 18377 23431 18411
rect 23431 18377 23440 18411
rect 23388 18368 23440 18377
rect 23480 18300 23532 18352
rect 24492 18368 24544 18420
rect 24584 18368 24636 18420
rect 26240 18368 26292 18420
rect 30288 18411 30340 18420
rect 30288 18377 30297 18411
rect 30297 18377 30331 18411
rect 30331 18377 30340 18411
rect 30288 18368 30340 18377
rect 34520 18368 34572 18420
rect 14372 18207 14424 18216
rect 14372 18173 14381 18207
rect 14381 18173 14415 18207
rect 14415 18173 14424 18207
rect 14372 18164 14424 18173
rect 10876 18096 10928 18105
rect 13728 18096 13780 18148
rect 8484 18028 8536 18080
rect 8944 18028 8996 18080
rect 12440 18028 12492 18080
rect 13084 18028 13136 18080
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 15292 18275 15344 18284
rect 15292 18241 15301 18275
rect 15301 18241 15335 18275
rect 15335 18241 15344 18275
rect 15292 18232 15344 18241
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 15844 18275 15896 18284
rect 15844 18241 15853 18275
rect 15853 18241 15887 18275
rect 15887 18241 15896 18275
rect 15844 18232 15896 18241
rect 15936 18232 15988 18284
rect 16212 18275 16264 18284
rect 16212 18241 16221 18275
rect 16221 18241 16255 18275
rect 16255 18241 16264 18275
rect 16212 18232 16264 18241
rect 17040 18275 17092 18284
rect 17040 18241 17049 18275
rect 17049 18241 17083 18275
rect 17083 18241 17092 18275
rect 17040 18232 17092 18241
rect 17408 18232 17460 18284
rect 17500 18275 17552 18284
rect 17500 18241 17509 18275
rect 17509 18241 17543 18275
rect 17543 18241 17552 18275
rect 17500 18232 17552 18241
rect 17592 18275 17644 18284
rect 17592 18241 17601 18275
rect 17601 18241 17635 18275
rect 17635 18241 17644 18275
rect 17592 18232 17644 18241
rect 16672 18164 16724 18216
rect 17224 18096 17276 18148
rect 17408 18096 17460 18148
rect 15384 18028 15436 18080
rect 15936 18028 15988 18080
rect 16488 18028 16540 18080
rect 19708 18275 19760 18284
rect 19708 18241 19717 18275
rect 19717 18241 19751 18275
rect 19751 18241 19760 18275
rect 19708 18232 19760 18241
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 21364 18275 21416 18284
rect 21364 18241 21373 18275
rect 21373 18241 21407 18275
rect 21407 18241 21416 18275
rect 21364 18232 21416 18241
rect 21824 18232 21876 18284
rect 18512 18164 18564 18216
rect 24308 18275 24360 18284
rect 24308 18241 24317 18275
rect 24317 18241 24351 18275
rect 24351 18241 24360 18275
rect 24308 18232 24360 18241
rect 25596 18300 25648 18352
rect 25688 18232 25740 18284
rect 25964 18300 26016 18352
rect 25228 18164 25280 18216
rect 25412 18207 25464 18216
rect 25412 18173 25421 18207
rect 25421 18173 25455 18207
rect 25455 18173 25464 18207
rect 25412 18164 25464 18173
rect 20720 18139 20772 18148
rect 20720 18105 20729 18139
rect 20729 18105 20763 18139
rect 20763 18105 20772 18139
rect 20720 18096 20772 18105
rect 23756 18139 23808 18148
rect 23756 18105 23765 18139
rect 23765 18105 23799 18139
rect 23799 18105 23808 18139
rect 23756 18096 23808 18105
rect 25136 18096 25188 18148
rect 25872 18275 25924 18284
rect 25872 18241 25881 18275
rect 25881 18241 25915 18275
rect 25915 18241 25924 18275
rect 25872 18232 25924 18241
rect 30196 18275 30248 18284
rect 24400 18071 24452 18080
rect 24400 18037 24409 18071
rect 24409 18037 24443 18071
rect 24443 18037 24452 18071
rect 24400 18028 24452 18037
rect 25228 18071 25280 18080
rect 25228 18037 25237 18071
rect 25237 18037 25271 18071
rect 25271 18037 25280 18071
rect 30196 18241 30205 18275
rect 30205 18241 30239 18275
rect 30239 18241 30248 18275
rect 30196 18232 30248 18241
rect 34796 18232 34848 18284
rect 25228 18028 25280 18037
rect 26056 18028 26108 18080
rect 30012 18071 30064 18080
rect 30012 18037 30021 18071
rect 30021 18037 30055 18071
rect 30055 18037 30064 18071
rect 30012 18028 30064 18037
rect 33048 18028 33100 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 6552 17824 6604 17876
rect 8300 17824 8352 17876
rect 13820 17824 13872 17876
rect 1676 17731 1728 17740
rect 1676 17697 1685 17731
rect 1685 17697 1719 17731
rect 1719 17697 1728 17731
rect 1676 17688 1728 17697
rect 2320 17552 2372 17604
rect 3056 17552 3108 17604
rect 4896 17552 4948 17604
rect 5264 17688 5316 17740
rect 6368 17688 6420 17740
rect 13728 17756 13780 17808
rect 11336 17688 11388 17740
rect 14280 17824 14332 17876
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 15200 17867 15252 17876
rect 15200 17833 15209 17867
rect 15209 17833 15243 17867
rect 15243 17833 15252 17867
rect 15200 17824 15252 17833
rect 15292 17824 15344 17876
rect 15844 17824 15896 17876
rect 16488 17867 16540 17876
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 6736 17595 6788 17604
rect 6736 17561 6745 17595
rect 6745 17561 6779 17595
rect 6779 17561 6788 17595
rect 6736 17552 6788 17561
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 11796 17620 11848 17672
rect 13268 17620 13320 17672
rect 9956 17552 10008 17604
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 3424 17527 3476 17536
rect 3424 17493 3433 17527
rect 3433 17493 3467 17527
rect 3467 17493 3476 17527
rect 3424 17484 3476 17493
rect 4160 17484 4212 17536
rect 5356 17527 5408 17536
rect 5356 17493 5365 17527
rect 5365 17493 5399 17527
rect 5399 17493 5408 17527
rect 5356 17484 5408 17493
rect 8208 17527 8260 17536
rect 8208 17493 8217 17527
rect 8217 17493 8251 17527
rect 8251 17493 8260 17527
rect 8208 17484 8260 17493
rect 8484 17484 8536 17536
rect 9588 17484 9640 17536
rect 14004 17620 14056 17672
rect 14096 17663 14148 17672
rect 14096 17629 14105 17663
rect 14105 17629 14139 17663
rect 14139 17629 14148 17663
rect 14096 17620 14148 17629
rect 14280 17663 14332 17672
rect 14280 17629 14289 17663
rect 14289 17629 14323 17663
rect 14323 17629 14332 17663
rect 15936 17756 15988 17808
rect 17500 17824 17552 17876
rect 21364 17824 21416 17876
rect 22928 17824 22980 17876
rect 23296 17824 23348 17876
rect 23480 17824 23532 17876
rect 25136 17867 25188 17876
rect 25136 17833 25145 17867
rect 25145 17833 25179 17867
rect 25179 17833 25188 17867
rect 25136 17824 25188 17833
rect 25964 17824 26016 17876
rect 26332 17824 26384 17876
rect 26608 17867 26660 17876
rect 26608 17833 26617 17867
rect 26617 17833 26651 17867
rect 26651 17833 26660 17867
rect 26608 17824 26660 17833
rect 20996 17756 21048 17808
rect 14280 17620 14332 17629
rect 14372 17552 14424 17604
rect 15476 17620 15528 17672
rect 11244 17484 11296 17536
rect 12348 17527 12400 17536
rect 12348 17493 12357 17527
rect 12357 17493 12391 17527
rect 12391 17493 12400 17527
rect 12348 17484 12400 17493
rect 12992 17484 13044 17536
rect 13176 17484 13228 17536
rect 14096 17484 14148 17536
rect 14740 17484 14792 17536
rect 15016 17527 15068 17536
rect 15016 17493 15025 17527
rect 15025 17493 15059 17527
rect 15059 17493 15068 17527
rect 15016 17484 15068 17493
rect 15384 17484 15436 17536
rect 15476 17484 15528 17536
rect 15936 17663 15988 17672
rect 15936 17629 15945 17663
rect 15945 17629 15979 17663
rect 15979 17629 15988 17663
rect 15936 17620 15988 17629
rect 16672 17688 16724 17740
rect 17684 17688 17736 17740
rect 19708 17688 19760 17740
rect 20352 17731 20404 17740
rect 20352 17697 20361 17731
rect 20361 17697 20395 17731
rect 20395 17697 20404 17731
rect 20352 17688 20404 17697
rect 16120 17595 16172 17604
rect 16120 17561 16129 17595
rect 16129 17561 16163 17595
rect 16163 17561 16172 17595
rect 16120 17552 16172 17561
rect 16580 17620 16632 17672
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 16856 17484 16908 17536
rect 17040 17484 17092 17536
rect 17776 17484 17828 17536
rect 19340 17663 19392 17672
rect 19340 17629 19349 17663
rect 19349 17629 19383 17663
rect 19383 17629 19392 17663
rect 19340 17620 19392 17629
rect 19432 17620 19484 17672
rect 25596 17688 25648 17740
rect 26516 17688 26568 17740
rect 24768 17620 24820 17672
rect 26792 17620 26844 17672
rect 20628 17484 20680 17536
rect 22928 17527 22980 17536
rect 22928 17493 22937 17527
rect 22937 17493 22971 17527
rect 22971 17493 22980 17527
rect 22928 17484 22980 17493
rect 25136 17484 25188 17536
rect 25412 17484 25464 17536
rect 26056 17484 26108 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 2320 17323 2372 17332
rect 2320 17289 2329 17323
rect 2329 17289 2363 17323
rect 2363 17289 2372 17323
rect 2320 17280 2372 17289
rect 3148 17280 3200 17332
rect 4988 17280 5040 17332
rect 5356 17280 5408 17332
rect 6736 17280 6788 17332
rect 8208 17280 8260 17332
rect 940 17144 992 17196
rect 2872 17144 2924 17196
rect 2872 17008 2924 17060
rect 4160 17187 4212 17196
rect 4160 17153 4169 17187
rect 4169 17153 4203 17187
rect 4203 17153 4212 17187
rect 4160 17144 4212 17153
rect 4620 17144 4672 17196
rect 3516 17119 3568 17128
rect 3516 17085 3525 17119
rect 3525 17085 3559 17119
rect 3559 17085 3568 17119
rect 3516 17076 3568 17085
rect 3976 17076 4028 17128
rect 4068 17119 4120 17128
rect 4068 17085 4077 17119
rect 4077 17085 4111 17119
rect 4111 17085 4120 17119
rect 4068 17076 4120 17085
rect 7380 17212 7432 17264
rect 9956 17323 10008 17332
rect 9956 17289 9965 17323
rect 9965 17289 9999 17323
rect 9999 17289 10008 17323
rect 9956 17280 10008 17289
rect 12348 17280 12400 17332
rect 15752 17280 15804 17332
rect 16028 17280 16080 17332
rect 16672 17280 16724 17332
rect 16948 17280 17000 17332
rect 17592 17323 17644 17332
rect 17592 17289 17601 17323
rect 17601 17289 17635 17323
rect 17635 17289 17644 17323
rect 17592 17280 17644 17289
rect 20996 17280 21048 17332
rect 21824 17323 21876 17332
rect 21824 17289 21833 17323
rect 21833 17289 21867 17323
rect 21867 17289 21876 17323
rect 21824 17280 21876 17289
rect 22928 17280 22980 17332
rect 9404 17212 9456 17264
rect 10968 17212 11020 17264
rect 11244 17212 11296 17264
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 9772 17076 9824 17128
rect 8024 17008 8076 17060
rect 8484 17008 8536 17060
rect 13084 17144 13136 17196
rect 13636 17187 13688 17196
rect 13636 17153 13645 17187
rect 13645 17153 13679 17187
rect 13679 17153 13688 17187
rect 13636 17144 13688 17153
rect 14004 17187 14056 17196
rect 14004 17153 14013 17187
rect 14013 17153 14047 17187
rect 14047 17153 14056 17187
rect 14004 17144 14056 17153
rect 11980 17076 12032 17128
rect 12624 17076 12676 17128
rect 14464 17144 14516 17196
rect 12992 17008 13044 17060
rect 3608 16940 3660 16992
rect 4620 16940 4672 16992
rect 14372 16940 14424 16992
rect 15844 17212 15896 17264
rect 14924 17187 14976 17196
rect 14924 17153 14933 17187
rect 14933 17153 14967 17187
rect 14967 17153 14976 17187
rect 14924 17144 14976 17153
rect 15016 17144 15068 17196
rect 16120 17144 16172 17196
rect 14740 17008 14792 17060
rect 15752 17119 15804 17128
rect 15752 17085 15761 17119
rect 15761 17085 15795 17119
rect 15795 17085 15804 17119
rect 15752 17076 15804 17085
rect 16764 17187 16816 17196
rect 16764 17153 16773 17187
rect 16773 17153 16807 17187
rect 16807 17153 16816 17187
rect 16764 17144 16816 17153
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17408 17255 17460 17264
rect 17408 17221 17417 17255
rect 17417 17221 17451 17255
rect 17451 17221 17460 17255
rect 17408 17212 17460 17221
rect 17316 17144 17368 17196
rect 17776 17187 17828 17196
rect 17776 17153 17785 17187
rect 17785 17153 17819 17187
rect 17819 17153 17828 17187
rect 17776 17144 17828 17153
rect 18144 17187 18196 17196
rect 18144 17153 18153 17187
rect 18153 17153 18187 17187
rect 18187 17153 18196 17187
rect 18144 17144 18196 17153
rect 19432 17144 19484 17196
rect 16856 17076 16908 17128
rect 20628 17076 20680 17128
rect 22560 17187 22612 17196
rect 22560 17153 22569 17187
rect 22569 17153 22603 17187
rect 22603 17153 22612 17187
rect 22560 17144 22612 17153
rect 20996 17076 21048 17128
rect 21640 17119 21692 17128
rect 21640 17085 21649 17119
rect 21649 17085 21683 17119
rect 21683 17085 21692 17119
rect 21640 17076 21692 17085
rect 22928 17187 22980 17196
rect 22928 17153 22937 17187
rect 22937 17153 22971 17187
rect 22971 17153 22980 17187
rect 22928 17144 22980 17153
rect 24032 17280 24084 17332
rect 24400 17280 24452 17332
rect 23296 17008 23348 17060
rect 23664 17187 23716 17196
rect 23664 17153 23673 17187
rect 23673 17153 23707 17187
rect 23707 17153 23716 17187
rect 23664 17144 23716 17153
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 23940 17144 23992 17196
rect 25872 17144 25924 17196
rect 26424 17212 26476 17264
rect 26700 17255 26752 17264
rect 26700 17221 26709 17255
rect 26709 17221 26743 17255
rect 26743 17221 26752 17255
rect 26700 17212 26752 17221
rect 26056 17076 26108 17128
rect 26332 17187 26384 17196
rect 26332 17153 26341 17187
rect 26341 17153 26375 17187
rect 26375 17153 26384 17187
rect 26332 17144 26384 17153
rect 26700 17008 26752 17060
rect 15108 16940 15160 16992
rect 17408 16940 17460 16992
rect 17684 16940 17736 16992
rect 24124 16940 24176 16992
rect 24860 16940 24912 16992
rect 26792 16983 26844 16992
rect 26792 16949 26801 16983
rect 26801 16949 26835 16983
rect 26835 16949 26844 16983
rect 26792 16940 26844 16949
rect 27252 16940 27304 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3516 16736 3568 16788
rect 7380 16736 7432 16788
rect 11244 16736 11296 16788
rect 4068 16668 4120 16720
rect 10692 16711 10744 16720
rect 10692 16677 10701 16711
rect 10701 16677 10735 16711
rect 10735 16677 10744 16711
rect 10692 16668 10744 16677
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 9588 16600 9640 16652
rect 11980 16779 12032 16788
rect 11980 16745 11989 16779
rect 11989 16745 12023 16779
rect 12023 16745 12032 16779
rect 11980 16736 12032 16745
rect 14464 16736 14516 16788
rect 14740 16779 14792 16788
rect 14740 16745 14749 16779
rect 14749 16745 14783 16779
rect 14783 16745 14792 16779
rect 14740 16736 14792 16745
rect 16764 16736 16816 16788
rect 16948 16779 17000 16788
rect 16948 16745 16957 16779
rect 16957 16745 16991 16779
rect 16991 16745 17000 16779
rect 16948 16736 17000 16745
rect 18052 16779 18104 16788
rect 18052 16745 18061 16779
rect 18061 16745 18095 16779
rect 18095 16745 18104 16779
rect 18052 16736 18104 16745
rect 18420 16736 18472 16788
rect 19432 16779 19484 16788
rect 19432 16745 19441 16779
rect 19441 16745 19475 16779
rect 19475 16745 19484 16779
rect 19432 16736 19484 16745
rect 22928 16736 22980 16788
rect 24860 16779 24912 16788
rect 24860 16745 24869 16779
rect 24869 16745 24903 16779
rect 24903 16745 24912 16779
rect 24860 16736 24912 16745
rect 25872 16736 25924 16788
rect 26240 16736 26292 16788
rect 4620 16532 4672 16584
rect 4988 16532 5040 16584
rect 8024 16396 8076 16448
rect 8484 16396 8536 16448
rect 11520 16600 11572 16652
rect 13544 16600 13596 16652
rect 13636 16532 13688 16584
rect 12992 16464 13044 16516
rect 14004 16464 14056 16516
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 23296 16668 23348 16720
rect 16580 16643 16632 16652
rect 16580 16609 16589 16643
rect 16589 16609 16623 16643
rect 16623 16609 16632 16643
rect 16580 16600 16632 16609
rect 16672 16532 16724 16584
rect 10508 16396 10560 16448
rect 11796 16396 11848 16448
rect 12440 16439 12492 16448
rect 12440 16405 12449 16439
rect 12449 16405 12483 16439
rect 12483 16405 12492 16439
rect 12440 16396 12492 16405
rect 13176 16396 13228 16448
rect 14096 16396 14148 16448
rect 14740 16464 14792 16516
rect 14924 16464 14976 16516
rect 17408 16532 17460 16584
rect 21640 16600 21692 16652
rect 18144 16532 18196 16584
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19248 16532 19300 16541
rect 22560 16532 22612 16584
rect 14372 16396 14424 16448
rect 17776 16396 17828 16448
rect 18696 16464 18748 16516
rect 23756 16600 23808 16652
rect 25964 16668 26016 16720
rect 23940 16575 23992 16584
rect 23940 16541 23949 16575
rect 23949 16541 23983 16575
rect 23983 16541 23992 16575
rect 23940 16532 23992 16541
rect 24124 16575 24176 16584
rect 24124 16541 24133 16575
rect 24133 16541 24167 16575
rect 24167 16541 24176 16575
rect 24124 16532 24176 16541
rect 24400 16532 24452 16584
rect 25136 16532 25188 16584
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 26056 16600 26108 16652
rect 24032 16464 24084 16516
rect 19432 16396 19484 16448
rect 23572 16396 23624 16448
rect 25412 16396 25464 16448
rect 25964 16575 26016 16584
rect 25964 16541 25973 16575
rect 25973 16541 26007 16575
rect 26007 16541 26016 16575
rect 25964 16532 26016 16541
rect 30012 16643 30064 16652
rect 26240 16575 26292 16584
rect 26240 16541 26249 16575
rect 26249 16541 26283 16575
rect 26283 16541 26292 16575
rect 26240 16532 26292 16541
rect 30012 16609 30021 16643
rect 30021 16609 30055 16643
rect 30055 16609 30064 16643
rect 30012 16600 30064 16609
rect 34612 16464 34664 16516
rect 25872 16396 25924 16448
rect 25964 16396 26016 16448
rect 26240 16439 26292 16448
rect 26240 16405 26249 16439
rect 26249 16405 26283 16439
rect 26283 16405 26292 16439
rect 26240 16396 26292 16405
rect 26516 16396 26568 16448
rect 29644 16439 29696 16448
rect 29644 16405 29653 16439
rect 29653 16405 29687 16439
rect 29687 16405 29696 16439
rect 29644 16396 29696 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11060 16192 11112 16244
rect 3976 16124 4028 16176
rect 3332 16056 3384 16108
rect 4068 16056 4120 16108
rect 4988 16056 5040 16108
rect 5448 16124 5500 16176
rect 13636 16192 13688 16244
rect 14648 16192 14700 16244
rect 15752 16192 15804 16244
rect 18328 16192 18380 16244
rect 18604 16192 18656 16244
rect 18972 16192 19024 16244
rect 19248 16192 19300 16244
rect 19340 16192 19392 16244
rect 19432 16192 19484 16244
rect 20628 16192 20680 16244
rect 8484 15988 8536 16040
rect 10508 15988 10560 16040
rect 11796 15988 11848 16040
rect 12072 16031 12124 16040
rect 12072 15997 12081 16031
rect 12081 15997 12115 16031
rect 12115 15997 12124 16031
rect 12072 15988 12124 15997
rect 4620 15920 4672 15972
rect 12440 16056 12492 16108
rect 12624 16056 12676 16108
rect 13268 16056 13320 16108
rect 4804 15895 4856 15904
rect 4804 15861 4813 15895
rect 4813 15861 4847 15895
rect 4847 15861 4856 15895
rect 4804 15852 4856 15861
rect 9956 15895 10008 15904
rect 9956 15861 9965 15895
rect 9965 15861 9999 15895
rect 9999 15861 10008 15895
rect 9956 15852 10008 15861
rect 11980 15852 12032 15904
rect 13176 16031 13228 16040
rect 13176 15997 13185 16031
rect 13185 15997 13219 16031
rect 13219 15997 13228 16031
rect 14004 16056 14056 16108
rect 14280 16056 14332 16108
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 13176 15988 13228 15997
rect 17776 16099 17828 16108
rect 17776 16065 17785 16099
rect 17785 16065 17819 16099
rect 17819 16065 17828 16099
rect 17776 16056 17828 16065
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 16396 15988 16448 16040
rect 18328 16099 18380 16108
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 18420 16099 18472 16108
rect 18420 16065 18429 16099
rect 18429 16065 18463 16099
rect 18463 16065 18472 16099
rect 18420 16056 18472 16065
rect 18696 16099 18748 16108
rect 18696 16065 18705 16099
rect 18705 16065 18739 16099
rect 18739 16065 18748 16099
rect 18696 16056 18748 16065
rect 19616 16167 19668 16176
rect 19616 16133 19625 16167
rect 19625 16133 19659 16167
rect 19659 16133 19668 16167
rect 19616 16124 19668 16133
rect 23388 16192 23440 16244
rect 23664 16192 23716 16244
rect 18972 16056 19024 16108
rect 19892 16056 19944 16108
rect 19984 16056 20036 16108
rect 21180 16099 21232 16108
rect 16764 15852 16816 15904
rect 17868 15920 17920 15972
rect 17040 15852 17092 15904
rect 17960 15852 18012 15904
rect 19340 15852 19392 15904
rect 19892 15852 19944 15904
rect 20076 15920 20128 15972
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 23848 16124 23900 16176
rect 25228 16192 25280 16244
rect 26148 16192 26200 16244
rect 32404 16192 32456 16244
rect 33048 16235 33100 16244
rect 33048 16201 33057 16235
rect 33057 16201 33091 16235
rect 33091 16201 33100 16235
rect 33048 16192 33100 16201
rect 22560 16056 22612 16108
rect 23296 16099 23348 16108
rect 23296 16065 23305 16099
rect 23305 16065 23339 16099
rect 23339 16065 23348 16099
rect 23296 16056 23348 16065
rect 21640 15988 21692 16040
rect 29644 16124 29696 16176
rect 25412 16099 25464 16108
rect 25412 16065 25421 16099
rect 25421 16065 25455 16099
rect 25455 16065 25464 16099
rect 25412 16056 25464 16065
rect 25872 16056 25924 16108
rect 26240 16099 26292 16108
rect 26240 16065 26249 16099
rect 26249 16065 26283 16099
rect 26283 16065 26292 16099
rect 26240 16056 26292 16065
rect 31944 16056 31996 16108
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 34152 16124 34204 16176
rect 26976 15988 27028 16040
rect 20996 15852 21048 15904
rect 22100 15852 22152 15904
rect 25136 15852 25188 15904
rect 25228 15895 25280 15904
rect 25228 15861 25237 15895
rect 25237 15861 25271 15895
rect 25271 15861 25280 15895
rect 25228 15852 25280 15861
rect 33416 16031 33468 16040
rect 33416 15997 33425 16031
rect 33425 15997 33459 16031
rect 33459 15997 33468 16031
rect 33416 15988 33468 15997
rect 29276 15852 29328 15904
rect 31116 15852 31168 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 3332 15691 3384 15700
rect 3332 15657 3341 15691
rect 3341 15657 3375 15691
rect 3375 15657 3384 15691
rect 3332 15648 3384 15657
rect 4804 15648 4856 15700
rect 5080 15648 5132 15700
rect 12072 15648 12124 15700
rect 12992 15648 13044 15700
rect 13360 15648 13412 15700
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 15200 15691 15252 15700
rect 15200 15657 15209 15691
rect 15209 15657 15243 15691
rect 15243 15657 15252 15691
rect 15200 15648 15252 15657
rect 17500 15691 17552 15700
rect 17500 15657 17509 15691
rect 17509 15657 17543 15691
rect 17543 15657 17552 15691
rect 17500 15648 17552 15657
rect 17868 15648 17920 15700
rect 17960 15648 18012 15700
rect 15108 15580 15160 15632
rect 18328 15580 18380 15632
rect 8484 15512 8536 15564
rect 3608 15487 3660 15496
rect 3608 15453 3617 15487
rect 3617 15453 3651 15487
rect 3651 15453 3660 15487
rect 3608 15444 3660 15453
rect 1860 15419 1912 15428
rect 1860 15385 1869 15419
rect 1869 15385 1903 15419
rect 1903 15385 1912 15419
rect 1860 15376 1912 15385
rect 1676 15308 1728 15360
rect 3792 15308 3844 15360
rect 4712 15444 4764 15496
rect 5908 15444 5960 15496
rect 8024 15487 8076 15496
rect 8024 15453 8033 15487
rect 8033 15453 8067 15487
rect 8067 15453 8076 15487
rect 8024 15444 8076 15453
rect 5448 15376 5500 15428
rect 5632 15376 5684 15428
rect 4896 15308 4948 15360
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 9956 15512 10008 15564
rect 12808 15512 12860 15564
rect 11980 15444 12032 15496
rect 12624 15444 12676 15496
rect 10600 15376 10652 15428
rect 8576 15308 8628 15360
rect 8760 15351 8812 15360
rect 8760 15317 8769 15351
rect 8769 15317 8803 15351
rect 8803 15317 8812 15351
rect 8760 15308 8812 15317
rect 11336 15351 11388 15360
rect 11336 15317 11345 15351
rect 11345 15317 11379 15351
rect 11379 15317 11388 15351
rect 11336 15308 11388 15317
rect 14464 15555 14516 15564
rect 14464 15521 14473 15555
rect 14473 15521 14507 15555
rect 14507 15521 14516 15555
rect 14464 15512 14516 15521
rect 13452 15444 13504 15496
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 14280 15487 14332 15496
rect 14280 15453 14289 15487
rect 14289 15453 14323 15487
rect 14323 15453 14332 15487
rect 14280 15444 14332 15453
rect 14648 15444 14700 15496
rect 15292 15512 15344 15564
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 16672 15512 16724 15564
rect 15016 15444 15068 15453
rect 14740 15308 14792 15360
rect 16120 15487 16172 15496
rect 16120 15453 16129 15487
rect 16129 15453 16163 15487
rect 16163 15453 16172 15487
rect 16120 15444 16172 15453
rect 16856 15376 16908 15428
rect 19524 15648 19576 15700
rect 25872 15648 25924 15700
rect 29276 15691 29328 15700
rect 29276 15657 29285 15691
rect 29285 15657 29319 15691
rect 29319 15657 29328 15691
rect 29276 15648 29328 15657
rect 33416 15648 33468 15700
rect 34152 15691 34204 15700
rect 34152 15657 34161 15691
rect 34161 15657 34195 15691
rect 34195 15657 34204 15691
rect 34152 15648 34204 15657
rect 18972 15580 19024 15632
rect 19156 15444 19208 15496
rect 26976 15512 27028 15564
rect 18604 15376 18656 15428
rect 18972 15419 19024 15428
rect 18972 15385 18981 15419
rect 18981 15385 19015 15419
rect 19015 15385 19024 15419
rect 18972 15376 19024 15385
rect 23388 15444 23440 15496
rect 20076 15419 20128 15428
rect 16672 15308 16724 15360
rect 17040 15351 17092 15360
rect 17040 15317 17049 15351
rect 17049 15317 17083 15351
rect 17083 15317 17092 15351
rect 17040 15308 17092 15317
rect 17224 15308 17276 15360
rect 17868 15351 17920 15360
rect 17868 15317 17877 15351
rect 17877 15317 17911 15351
rect 17911 15317 17920 15351
rect 17868 15308 17920 15317
rect 18420 15308 18472 15360
rect 18880 15308 18932 15360
rect 20076 15385 20085 15419
rect 20085 15385 20119 15419
rect 20119 15385 20128 15419
rect 20076 15376 20128 15385
rect 22744 15376 22796 15428
rect 23480 15376 23532 15428
rect 27528 15444 27580 15496
rect 31208 15444 31260 15496
rect 32312 15580 32364 15632
rect 32588 15580 32640 15632
rect 27160 15376 27212 15428
rect 29000 15376 29052 15428
rect 34336 15444 34388 15496
rect 19340 15308 19392 15360
rect 19984 15308 20036 15360
rect 20996 15351 21048 15360
rect 20996 15317 21005 15351
rect 21005 15317 21039 15351
rect 21039 15317 21048 15351
rect 20996 15308 21048 15317
rect 21088 15308 21140 15360
rect 21916 15308 21968 15360
rect 23204 15308 23256 15360
rect 23664 15308 23716 15360
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 25228 15308 25280 15360
rect 25688 15308 25740 15360
rect 26516 15308 26568 15360
rect 27620 15308 27672 15360
rect 31944 15308 31996 15360
rect 33876 15351 33928 15360
rect 33876 15317 33885 15351
rect 33885 15317 33919 15351
rect 33919 15317 33928 15351
rect 33876 15308 33928 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1860 15104 1912 15156
rect 10600 15104 10652 15156
rect 11336 15104 11388 15156
rect 11980 15036 12032 15088
rect 940 14968 992 15020
rect 7748 14968 7800 15020
rect 10416 14900 10468 14952
rect 3516 14807 3568 14816
rect 3516 14773 3525 14807
rect 3525 14773 3559 14807
rect 3559 14773 3568 14807
rect 3516 14764 3568 14773
rect 5908 14764 5960 14816
rect 10508 14875 10560 14884
rect 10508 14841 10517 14875
rect 10517 14841 10551 14875
rect 10551 14841 10560 14875
rect 11612 15011 11664 15020
rect 11612 14977 11621 15011
rect 11621 14977 11655 15011
rect 11655 14977 11664 15011
rect 11612 14968 11664 14977
rect 14096 15147 14148 15156
rect 14096 15113 14105 15147
rect 14105 15113 14139 15147
rect 14139 15113 14148 15147
rect 14096 15104 14148 15113
rect 14280 15147 14332 15156
rect 14280 15113 14289 15147
rect 14289 15113 14323 15147
rect 14323 15113 14332 15147
rect 14280 15104 14332 15113
rect 15292 15079 15344 15088
rect 15292 15045 15301 15079
rect 15301 15045 15335 15079
rect 15335 15045 15344 15079
rect 15292 15036 15344 15045
rect 17316 15036 17368 15088
rect 19156 15079 19208 15088
rect 19156 15045 19165 15079
rect 19165 15045 19199 15079
rect 19199 15045 19208 15079
rect 19156 15036 19208 15045
rect 13452 14968 13504 15020
rect 13636 14943 13688 14952
rect 13636 14909 13645 14943
rect 13645 14909 13679 14943
rect 13679 14909 13688 14943
rect 13636 14900 13688 14909
rect 14372 15011 14424 15020
rect 14372 14977 14381 15011
rect 14381 14977 14415 15011
rect 14415 14977 14424 15011
rect 14372 14968 14424 14977
rect 14740 14900 14792 14952
rect 14924 15011 14976 15020
rect 14924 14977 14933 15011
rect 14933 14977 14967 15011
rect 14967 14977 14976 15011
rect 14924 14968 14976 14977
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 16120 14968 16172 15020
rect 16580 14900 16632 14952
rect 16856 14968 16908 15020
rect 17500 14968 17552 15020
rect 18972 14968 19024 15020
rect 21916 15079 21968 15088
rect 21916 15045 21925 15079
rect 21925 15045 21959 15079
rect 21959 15045 21968 15079
rect 21916 15036 21968 15045
rect 22284 15104 22336 15156
rect 23204 15036 23256 15088
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 22100 14968 22152 15020
rect 20812 14900 20864 14952
rect 22192 14900 22244 14952
rect 22560 14968 22612 15020
rect 22836 14968 22888 15020
rect 10508 14832 10560 14841
rect 13820 14764 13872 14816
rect 17224 14764 17276 14816
rect 20812 14764 20864 14816
rect 23572 14968 23624 15020
rect 24308 15011 24360 15020
rect 24308 14977 24317 15011
rect 24317 14977 24351 15011
rect 24351 14977 24360 15011
rect 24308 14968 24360 14977
rect 24584 15011 24636 15020
rect 24584 14977 24593 15011
rect 24593 14977 24627 15011
rect 24627 14977 24636 15011
rect 24584 14968 24636 14977
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 24768 14968 24820 14977
rect 25228 14968 25280 15020
rect 23756 14943 23808 14952
rect 23756 14909 23765 14943
rect 23765 14909 23799 14943
rect 23799 14909 23808 14943
rect 23756 14900 23808 14909
rect 24124 14832 24176 14884
rect 26332 14943 26384 14952
rect 26332 14909 26341 14943
rect 26341 14909 26375 14943
rect 26375 14909 26384 14943
rect 26332 14900 26384 14909
rect 27160 15104 27212 15156
rect 26608 14900 26660 14952
rect 26792 15011 26844 15020
rect 26792 14977 26801 15011
rect 26801 14977 26835 15011
rect 26835 14977 26844 15011
rect 26792 14968 26844 14977
rect 27252 15011 27304 15020
rect 27252 14977 27261 15011
rect 27261 14977 27295 15011
rect 27295 14977 27304 15011
rect 27252 14968 27304 14977
rect 27068 14900 27120 14952
rect 27620 15147 27672 15156
rect 27620 15113 27629 15147
rect 27629 15113 27663 15147
rect 27663 15113 27672 15147
rect 27620 15104 27672 15113
rect 32588 15104 32640 15156
rect 27804 14968 27856 15020
rect 27528 14900 27580 14952
rect 29000 14900 29052 14952
rect 26240 14832 26292 14884
rect 22376 14764 22428 14816
rect 22468 14764 22520 14816
rect 22928 14807 22980 14816
rect 22928 14773 22937 14807
rect 22937 14773 22971 14807
rect 22971 14773 22980 14807
rect 22928 14764 22980 14773
rect 23020 14807 23072 14816
rect 23020 14773 23029 14807
rect 23029 14773 23063 14807
rect 23063 14773 23072 14807
rect 23020 14764 23072 14773
rect 23112 14764 23164 14816
rect 28264 14807 28316 14816
rect 28264 14773 28273 14807
rect 28273 14773 28307 14807
rect 28307 14773 28316 14807
rect 28264 14764 28316 14773
rect 29460 14764 29512 14816
rect 30012 14968 30064 15020
rect 30380 14968 30432 15020
rect 31208 15011 31260 15020
rect 31208 14977 31217 15011
rect 31217 14977 31251 15011
rect 31251 14977 31260 15011
rect 31208 14968 31260 14977
rect 31852 14968 31904 15020
rect 32680 15011 32732 15020
rect 32680 14977 32689 15011
rect 32689 14977 32723 15011
rect 32723 14977 32732 15011
rect 32680 14968 32732 14977
rect 29920 14807 29972 14816
rect 29920 14773 29929 14807
rect 29929 14773 29963 14807
rect 29963 14773 29972 14807
rect 29920 14764 29972 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4988 14560 5040 14612
rect 5172 14560 5224 14612
rect 5264 14603 5316 14612
rect 5264 14569 5273 14603
rect 5273 14569 5307 14603
rect 5307 14569 5316 14603
rect 5264 14560 5316 14569
rect 5356 14560 5408 14612
rect 11612 14560 11664 14612
rect 11980 14560 12032 14612
rect 13636 14560 13688 14612
rect 14372 14560 14424 14612
rect 14740 14560 14792 14612
rect 16580 14603 16632 14612
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 13452 14492 13504 14544
rect 14924 14492 14976 14544
rect 5908 14424 5960 14476
rect 16764 14424 16816 14476
rect 4804 14331 4856 14340
rect 4804 14297 4813 14331
rect 4813 14297 4847 14331
rect 4847 14297 4856 14331
rect 4804 14288 4856 14297
rect 5264 14356 5316 14408
rect 5540 14356 5592 14408
rect 8576 14399 8628 14408
rect 8576 14365 8585 14399
rect 8585 14365 8619 14399
rect 8619 14365 8628 14399
rect 8576 14356 8628 14365
rect 8760 14356 8812 14408
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 5080 14220 5132 14272
rect 5356 14220 5408 14272
rect 6552 14220 6604 14272
rect 9128 14288 9180 14340
rect 9772 14288 9824 14340
rect 17224 14399 17276 14408
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17592 14424 17644 14476
rect 18972 14424 19024 14476
rect 21180 14560 21232 14612
rect 20904 14535 20956 14544
rect 20904 14501 20913 14535
rect 20913 14501 20947 14535
rect 20947 14501 20956 14535
rect 20904 14492 20956 14501
rect 22744 14492 22796 14544
rect 11152 14263 11204 14272
rect 11152 14229 11161 14263
rect 11161 14229 11195 14263
rect 11195 14229 11204 14263
rect 11152 14220 11204 14229
rect 15384 14263 15436 14272
rect 15384 14229 15393 14263
rect 15393 14229 15427 14263
rect 15427 14229 15436 14263
rect 15384 14220 15436 14229
rect 15936 14220 15988 14272
rect 20628 14356 20680 14408
rect 22928 14424 22980 14476
rect 20444 14331 20496 14340
rect 20444 14297 20453 14331
rect 20453 14297 20487 14331
rect 20487 14297 20496 14331
rect 20444 14288 20496 14297
rect 21272 14356 21324 14408
rect 21824 14399 21876 14408
rect 21824 14365 21833 14399
rect 21833 14365 21867 14399
rect 21867 14365 21876 14399
rect 21824 14356 21876 14365
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 17040 14263 17092 14272
rect 17040 14229 17049 14263
rect 17049 14229 17083 14263
rect 17083 14229 17092 14263
rect 17040 14220 17092 14229
rect 17408 14220 17460 14272
rect 18972 14220 19024 14272
rect 19340 14220 19392 14272
rect 20076 14263 20128 14272
rect 20076 14229 20085 14263
rect 20085 14229 20119 14263
rect 20119 14229 20128 14263
rect 20076 14220 20128 14229
rect 20352 14263 20404 14272
rect 20352 14229 20354 14263
rect 20354 14229 20388 14263
rect 20388 14229 20404 14263
rect 20352 14220 20404 14229
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 20812 14220 20864 14272
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 21272 14220 21324 14272
rect 22376 14263 22428 14272
rect 22376 14229 22385 14263
rect 22385 14229 22419 14263
rect 22419 14229 22428 14263
rect 22376 14220 22428 14229
rect 22928 14288 22980 14340
rect 23112 14399 23164 14408
rect 23112 14365 23121 14399
rect 23121 14365 23155 14399
rect 23155 14365 23164 14399
rect 23112 14356 23164 14365
rect 23204 14356 23256 14408
rect 23572 14492 23624 14544
rect 24308 14560 24360 14612
rect 26608 14560 26660 14612
rect 31852 14560 31904 14612
rect 26516 14492 26568 14544
rect 26792 14492 26844 14544
rect 27068 14424 27120 14476
rect 23480 14399 23532 14408
rect 23480 14365 23489 14399
rect 23489 14365 23523 14399
rect 23523 14365 23532 14399
rect 23480 14356 23532 14365
rect 23664 14399 23716 14408
rect 23664 14365 23673 14399
rect 23673 14365 23707 14399
rect 23707 14365 23716 14399
rect 23664 14356 23716 14365
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 23756 14356 23808 14365
rect 25504 14399 25556 14408
rect 25504 14365 25513 14399
rect 25513 14365 25547 14399
rect 25547 14365 25556 14399
rect 25504 14356 25556 14365
rect 28264 14492 28316 14544
rect 29276 14535 29328 14544
rect 29276 14501 29285 14535
rect 29285 14501 29319 14535
rect 29319 14501 29328 14535
rect 33048 14560 33100 14612
rect 29276 14492 29328 14501
rect 31852 14467 31904 14476
rect 31852 14433 31861 14467
rect 31861 14433 31895 14467
rect 31895 14433 31904 14467
rect 31852 14424 31904 14433
rect 24584 14288 24636 14340
rect 22836 14220 22888 14272
rect 27988 14399 28040 14408
rect 27988 14365 27997 14399
rect 27997 14365 28031 14399
rect 28031 14365 28040 14399
rect 27988 14356 28040 14365
rect 28172 14356 28224 14408
rect 29460 14356 29512 14408
rect 31300 14356 31352 14408
rect 26424 14220 26476 14272
rect 27436 14220 27488 14272
rect 29920 14288 29972 14340
rect 31760 14220 31812 14272
rect 32220 14220 32272 14272
rect 34612 14288 34664 14340
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4804 14016 4856 14068
rect 5172 14016 5224 14068
rect 2872 13991 2924 14000
rect 2872 13957 2881 13991
rect 2881 13957 2915 13991
rect 2915 13957 2924 13991
rect 2872 13948 2924 13957
rect 3884 13948 3936 14000
rect 5540 13948 5592 14000
rect 5356 13923 5408 13932
rect 5356 13889 5365 13923
rect 5365 13889 5399 13923
rect 5399 13889 5408 13923
rect 5356 13880 5408 13889
rect 3516 13812 3568 13864
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 8760 14016 8812 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10508 14016 10560 14068
rect 11520 14016 11572 14068
rect 13544 14016 13596 14068
rect 14556 14016 14608 14068
rect 16120 14059 16172 14068
rect 16120 14025 16129 14059
rect 16129 14025 16163 14059
rect 16163 14025 16172 14059
rect 16120 14016 16172 14025
rect 20444 14016 20496 14068
rect 21180 14016 21232 14068
rect 21272 14016 21324 14068
rect 21824 14016 21876 14068
rect 23388 14016 23440 14068
rect 23756 14016 23808 14068
rect 25504 14016 25556 14068
rect 11152 13880 11204 13932
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 15384 13880 15436 13932
rect 5172 13787 5224 13796
rect 5172 13753 5181 13787
rect 5181 13753 5215 13787
rect 5215 13753 5224 13787
rect 5172 13744 5224 13753
rect 5264 13787 5316 13796
rect 5264 13753 5273 13787
rect 5273 13753 5307 13787
rect 5307 13753 5316 13787
rect 5264 13744 5316 13753
rect 6920 13744 6972 13796
rect 12900 13744 12952 13796
rect 14924 13744 14976 13796
rect 16856 13923 16908 13932
rect 16856 13889 16865 13923
rect 16865 13889 16899 13923
rect 16899 13889 16908 13923
rect 16856 13880 16908 13889
rect 4896 13719 4948 13728
rect 4896 13685 4905 13719
rect 4905 13685 4939 13719
rect 4939 13685 4948 13719
rect 4896 13676 4948 13685
rect 9128 13676 9180 13728
rect 14188 13676 14240 13728
rect 15844 13812 15896 13864
rect 17408 13923 17460 13932
rect 17408 13889 17417 13923
rect 17417 13889 17451 13923
rect 17451 13889 17460 13923
rect 17408 13880 17460 13889
rect 17684 13880 17736 13932
rect 19248 13923 19300 13932
rect 19248 13889 19257 13923
rect 19257 13889 19291 13923
rect 19291 13889 19300 13923
rect 19248 13880 19300 13889
rect 19340 13880 19392 13932
rect 19432 13923 19484 13932
rect 19432 13889 19441 13923
rect 19441 13889 19475 13923
rect 19475 13889 19484 13923
rect 19432 13880 19484 13889
rect 18880 13812 18932 13864
rect 19524 13855 19576 13864
rect 19524 13821 19533 13855
rect 19533 13821 19567 13855
rect 19567 13821 19576 13855
rect 19524 13812 19576 13821
rect 20076 13948 20128 14000
rect 20536 13880 20588 13932
rect 21088 13948 21140 14000
rect 22376 13948 22428 14000
rect 21548 13923 21600 13932
rect 21548 13889 21557 13923
rect 21557 13889 21591 13923
rect 21591 13889 21600 13923
rect 21548 13880 21600 13889
rect 22928 13880 22980 13932
rect 25228 13991 25280 14000
rect 25228 13957 25237 13991
rect 25237 13957 25271 13991
rect 25271 13957 25280 13991
rect 25228 13948 25280 13957
rect 26148 14016 26200 14068
rect 26240 14016 26292 14068
rect 26332 14016 26384 14068
rect 26424 14016 26476 14068
rect 18420 13787 18472 13796
rect 18420 13753 18429 13787
rect 18429 13753 18463 13787
rect 18463 13753 18472 13787
rect 18420 13744 18472 13753
rect 19340 13744 19392 13796
rect 20352 13744 20404 13796
rect 21272 13855 21324 13864
rect 21272 13821 21281 13855
rect 21281 13821 21315 13855
rect 21315 13821 21324 13855
rect 21272 13812 21324 13821
rect 25228 13812 25280 13864
rect 25596 13880 25648 13932
rect 25780 13923 25832 13932
rect 25780 13889 25789 13923
rect 25789 13889 25823 13923
rect 25823 13889 25832 13923
rect 25780 13880 25832 13889
rect 26056 13923 26108 13932
rect 26056 13889 26065 13923
rect 26065 13889 26099 13923
rect 26099 13889 26108 13923
rect 26056 13880 26108 13889
rect 27252 14016 27304 14068
rect 25504 13744 25556 13796
rect 26240 13744 26292 13796
rect 27528 13880 27580 13932
rect 27988 14016 28040 14068
rect 29276 14059 29328 14068
rect 29276 14025 29285 14059
rect 29285 14025 29319 14059
rect 29319 14025 29328 14059
rect 29276 14016 29328 14025
rect 30472 13948 30524 14000
rect 31760 13948 31812 14000
rect 34060 13948 34112 14000
rect 27252 13787 27304 13796
rect 27252 13753 27261 13787
rect 27261 13753 27295 13787
rect 27295 13753 27304 13787
rect 27252 13744 27304 13753
rect 18788 13676 18840 13728
rect 22836 13676 22888 13728
rect 25780 13676 25832 13728
rect 27436 13744 27488 13796
rect 27620 13744 27672 13796
rect 31300 13744 31352 13796
rect 29368 13676 29420 13728
rect 33048 13923 33100 13932
rect 33048 13889 33057 13923
rect 33057 13889 33091 13923
rect 33091 13889 33100 13923
rect 33048 13880 33100 13889
rect 32220 13855 32272 13864
rect 32220 13821 32229 13855
rect 32229 13821 32263 13855
rect 32263 13821 32272 13855
rect 32220 13812 32272 13821
rect 31944 13744 31996 13796
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 4620 13472 4672 13524
rect 4804 13472 4856 13524
rect 6920 13472 6972 13524
rect 12440 13472 12492 13524
rect 13544 13515 13596 13524
rect 13544 13481 13553 13515
rect 13553 13481 13587 13515
rect 13587 13481 13596 13515
rect 13544 13472 13596 13481
rect 13820 13515 13872 13524
rect 13820 13481 13829 13515
rect 13829 13481 13863 13515
rect 13863 13481 13872 13515
rect 13820 13472 13872 13481
rect 15384 13472 15436 13524
rect 15752 13515 15804 13524
rect 15752 13481 15761 13515
rect 15761 13481 15795 13515
rect 15795 13481 15804 13515
rect 15752 13472 15804 13481
rect 16212 13472 16264 13524
rect 1676 13336 1728 13388
rect 1676 13243 1728 13252
rect 1676 13209 1685 13243
rect 1685 13209 1719 13243
rect 1719 13209 1728 13243
rect 1676 13200 1728 13209
rect 2320 13200 2372 13252
rect 4896 13336 4948 13388
rect 3516 13175 3568 13184
rect 3516 13141 3525 13175
rect 3525 13141 3559 13175
rect 3559 13141 3568 13175
rect 3516 13132 3568 13141
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 7012 13268 7064 13277
rect 9128 13311 9180 13320
rect 9128 13277 9137 13311
rect 9137 13277 9171 13311
rect 9171 13277 9180 13311
rect 9128 13268 9180 13277
rect 11980 13336 12032 13388
rect 10416 13311 10468 13320
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 17592 13447 17644 13456
rect 17592 13413 17601 13447
rect 17601 13413 17635 13447
rect 17635 13413 17644 13447
rect 17592 13404 17644 13413
rect 14924 13336 14976 13388
rect 15844 13336 15896 13388
rect 16304 13311 16356 13320
rect 14280 13200 14332 13252
rect 16304 13277 16313 13311
rect 16313 13277 16347 13311
rect 16347 13277 16356 13311
rect 16304 13268 16356 13277
rect 14556 13243 14608 13252
rect 14556 13209 14565 13243
rect 14565 13209 14599 13243
rect 14599 13209 14608 13243
rect 14556 13200 14608 13209
rect 17040 13268 17092 13320
rect 17684 13268 17736 13320
rect 19248 13472 19300 13524
rect 19984 13472 20036 13524
rect 21548 13472 21600 13524
rect 23112 13472 23164 13524
rect 26332 13515 26384 13524
rect 26332 13481 26341 13515
rect 26341 13481 26375 13515
rect 26375 13481 26384 13515
rect 26332 13472 26384 13481
rect 29368 13472 29420 13524
rect 30380 13515 30432 13524
rect 30380 13481 30389 13515
rect 30389 13481 30423 13515
rect 30423 13481 30432 13515
rect 30380 13472 30432 13481
rect 30472 13472 30524 13524
rect 34060 13472 34112 13524
rect 19340 13404 19392 13456
rect 18512 13336 18564 13388
rect 18880 13311 18932 13320
rect 18880 13277 18889 13311
rect 18889 13277 18923 13311
rect 18923 13277 18932 13311
rect 18880 13268 18932 13277
rect 19064 13311 19116 13320
rect 19064 13277 19073 13311
rect 19073 13277 19107 13311
rect 19107 13277 19116 13311
rect 19064 13268 19116 13277
rect 18328 13200 18380 13252
rect 19432 13268 19484 13320
rect 20076 13268 20128 13320
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 20536 13268 20588 13320
rect 20904 13336 20956 13388
rect 21088 13336 21140 13388
rect 21272 13268 21324 13320
rect 22928 13311 22980 13320
rect 22928 13277 22937 13311
rect 22937 13277 22971 13311
rect 22971 13277 22980 13311
rect 22928 13268 22980 13277
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13544 13132 13596 13184
rect 14188 13132 14240 13184
rect 17408 13175 17460 13184
rect 17408 13141 17417 13175
rect 17417 13141 17451 13175
rect 17451 13141 17460 13175
rect 17408 13132 17460 13141
rect 17500 13132 17552 13184
rect 17960 13132 18012 13184
rect 18512 13132 18564 13184
rect 18788 13132 18840 13184
rect 19156 13132 19208 13184
rect 21364 13200 21416 13252
rect 23204 13268 23256 13320
rect 23388 13311 23440 13320
rect 23388 13277 23397 13311
rect 23397 13277 23431 13311
rect 23431 13277 23440 13311
rect 23388 13268 23440 13277
rect 23848 13268 23900 13320
rect 25044 13404 25096 13456
rect 25596 13336 25648 13388
rect 20260 13175 20312 13184
rect 20260 13141 20269 13175
rect 20269 13141 20303 13175
rect 20303 13141 20312 13175
rect 20260 13132 20312 13141
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20628 13132 20680 13141
rect 20812 13132 20864 13184
rect 23020 13175 23072 13184
rect 23020 13141 23029 13175
rect 23029 13141 23063 13175
rect 23063 13141 23072 13175
rect 23020 13132 23072 13141
rect 23756 13132 23808 13184
rect 25228 13311 25280 13320
rect 25228 13277 25237 13311
rect 25237 13277 25271 13311
rect 25271 13277 25280 13311
rect 25228 13268 25280 13277
rect 25412 13175 25464 13184
rect 25412 13141 25421 13175
rect 25421 13141 25455 13175
rect 25455 13141 25464 13175
rect 25412 13132 25464 13141
rect 27436 13336 27488 13388
rect 27988 13311 28040 13320
rect 27988 13277 27997 13311
rect 27997 13277 28031 13311
rect 28031 13277 28040 13311
rect 27988 13268 28040 13277
rect 31760 13268 31812 13320
rect 31300 13200 31352 13252
rect 32680 13311 32732 13320
rect 32680 13277 32689 13311
rect 32689 13277 32723 13311
rect 32723 13277 32732 13311
rect 32680 13268 32732 13277
rect 33876 13243 33928 13252
rect 33876 13209 33885 13243
rect 33885 13209 33919 13243
rect 33919 13209 33928 13243
rect 33876 13200 33928 13209
rect 26424 13132 26476 13184
rect 27252 13132 27304 13184
rect 32404 13175 32456 13184
rect 32404 13141 32413 13175
rect 32413 13141 32447 13175
rect 32447 13141 32456 13175
rect 32404 13132 32456 13141
rect 34428 13175 34480 13184
rect 34428 13141 34437 13175
rect 34437 13141 34471 13175
rect 34471 13141 34480 13175
rect 34428 13132 34480 13141
rect 34520 13132 34572 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 5264 12928 5316 12980
rect 5540 12928 5592 12980
rect 4988 12860 5040 12912
rect 5448 12903 5500 12912
rect 5448 12869 5457 12903
rect 5457 12869 5491 12903
rect 5491 12869 5500 12903
rect 5448 12860 5500 12869
rect 940 12792 992 12844
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 3516 12588 3568 12640
rect 5632 12631 5684 12640
rect 5632 12597 5641 12631
rect 5641 12597 5675 12631
rect 5675 12597 5684 12631
rect 5632 12588 5684 12597
rect 5816 12631 5868 12640
rect 5816 12597 5825 12631
rect 5825 12597 5859 12631
rect 5859 12597 5868 12631
rect 5816 12588 5868 12597
rect 8300 12588 8352 12640
rect 8760 12656 8812 12708
rect 10416 12928 10468 12980
rect 12992 12928 13044 12980
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 14188 12928 14240 12980
rect 14556 12928 14608 12980
rect 16304 12928 16356 12980
rect 17500 12928 17552 12980
rect 12624 12835 12676 12844
rect 12624 12801 12633 12835
rect 12633 12801 12667 12835
rect 12667 12801 12676 12835
rect 12624 12792 12676 12801
rect 12808 12835 12860 12844
rect 12808 12801 12817 12835
rect 12817 12801 12851 12835
rect 12851 12801 12860 12835
rect 12808 12792 12860 12801
rect 10968 12656 11020 12708
rect 13912 12792 13964 12844
rect 14280 12835 14332 12844
rect 14280 12801 14289 12835
rect 14289 12801 14323 12835
rect 14323 12801 14332 12835
rect 14280 12792 14332 12801
rect 15660 12860 15712 12912
rect 16672 12860 16724 12912
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 15936 12835 15988 12844
rect 14832 12767 14884 12776
rect 14832 12733 14841 12767
rect 14841 12733 14875 12767
rect 14875 12733 14884 12767
rect 14832 12724 14884 12733
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 15568 12724 15620 12776
rect 16212 12792 16264 12844
rect 16856 12792 16908 12844
rect 19064 12928 19116 12980
rect 19156 12971 19208 12980
rect 19156 12937 19165 12971
rect 19165 12937 19199 12971
rect 19199 12937 19208 12971
rect 19156 12928 19208 12937
rect 15660 12699 15712 12708
rect 8668 12588 8720 12640
rect 9128 12588 9180 12640
rect 12440 12588 12492 12640
rect 14280 12588 14332 12640
rect 15108 12588 15160 12640
rect 15660 12665 15669 12699
rect 15669 12665 15703 12699
rect 15703 12665 15712 12699
rect 15660 12656 15712 12665
rect 15936 12656 15988 12708
rect 16856 12656 16908 12708
rect 17500 12724 17552 12776
rect 18972 12860 19024 12912
rect 19340 12903 19392 12912
rect 19340 12869 19349 12903
rect 19349 12869 19383 12903
rect 19383 12869 19392 12903
rect 19340 12860 19392 12869
rect 19524 12971 19576 12980
rect 19524 12937 19549 12971
rect 19549 12937 19576 12971
rect 19524 12928 19576 12937
rect 20444 12928 20496 12980
rect 23664 12928 23716 12980
rect 24584 12928 24636 12980
rect 24676 12928 24728 12980
rect 25044 12928 25096 12980
rect 25228 12928 25280 12980
rect 25320 12928 25372 12980
rect 20904 12860 20956 12912
rect 18420 12792 18472 12844
rect 20168 12792 20220 12844
rect 23388 12835 23440 12844
rect 23388 12801 23397 12835
rect 23397 12801 23431 12835
rect 23431 12801 23440 12835
rect 23388 12792 23440 12801
rect 24400 12792 24452 12844
rect 24492 12792 24544 12844
rect 24952 12835 25004 12844
rect 24952 12801 24961 12835
rect 24961 12801 24995 12835
rect 24995 12801 25004 12835
rect 24952 12792 25004 12801
rect 19340 12724 19392 12776
rect 19524 12724 19576 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 23848 12724 23900 12776
rect 24124 12767 24176 12776
rect 24124 12733 24133 12767
rect 24133 12733 24167 12767
rect 24167 12733 24176 12767
rect 24124 12724 24176 12733
rect 24308 12724 24360 12776
rect 25044 12767 25096 12776
rect 25044 12733 25053 12767
rect 25053 12733 25087 12767
rect 25087 12733 25096 12767
rect 25044 12724 25096 12733
rect 25504 12724 25556 12776
rect 25780 12792 25832 12844
rect 25872 12835 25924 12844
rect 25872 12801 25881 12835
rect 25881 12801 25915 12835
rect 25915 12801 25924 12835
rect 25872 12792 25924 12801
rect 26148 12835 26200 12844
rect 26148 12801 26157 12835
rect 26157 12801 26191 12835
rect 26191 12801 26200 12835
rect 26148 12792 26200 12801
rect 26424 12835 26476 12844
rect 26424 12801 26433 12835
rect 26433 12801 26467 12835
rect 26467 12801 26476 12835
rect 26424 12792 26476 12801
rect 27620 12928 27672 12980
rect 27988 12928 28040 12980
rect 17592 12656 17644 12708
rect 19064 12656 19116 12708
rect 21548 12656 21600 12708
rect 23756 12699 23808 12708
rect 23756 12665 23765 12699
rect 23765 12665 23799 12699
rect 23799 12665 23808 12699
rect 23756 12656 23808 12665
rect 15292 12631 15344 12640
rect 15292 12597 15301 12631
rect 15301 12597 15335 12631
rect 15335 12597 15344 12631
rect 15292 12588 15344 12597
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 17224 12588 17276 12640
rect 17960 12588 18012 12640
rect 18880 12588 18932 12640
rect 19340 12588 19392 12640
rect 20076 12588 20128 12640
rect 20444 12588 20496 12640
rect 24216 12631 24268 12640
rect 24216 12597 24225 12631
rect 24225 12597 24259 12631
rect 24259 12597 24268 12631
rect 24216 12588 24268 12597
rect 24308 12631 24360 12640
rect 24308 12597 24317 12631
rect 24317 12597 24351 12631
rect 24351 12597 24360 12631
rect 24308 12588 24360 12597
rect 24860 12656 24912 12708
rect 25320 12656 25372 12708
rect 25596 12656 25648 12708
rect 26056 12724 26108 12776
rect 27160 12792 27212 12844
rect 29276 12928 29328 12980
rect 32404 12928 32456 12980
rect 33048 12928 33100 12980
rect 29644 12860 29696 12912
rect 25780 12656 25832 12708
rect 27712 12792 27764 12844
rect 28632 12835 28684 12844
rect 28632 12801 28641 12835
rect 28641 12801 28675 12835
rect 28675 12801 28684 12835
rect 28632 12792 28684 12801
rect 33048 12835 33100 12844
rect 33048 12801 33057 12835
rect 33057 12801 33091 12835
rect 33091 12801 33100 12835
rect 33048 12792 33100 12801
rect 34428 12792 34480 12844
rect 30840 12588 30892 12640
rect 34428 12588 34480 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3516 12384 3568 12436
rect 5356 12384 5408 12436
rect 12808 12316 12860 12368
rect 5816 12291 5868 12300
rect 5816 12257 5825 12291
rect 5825 12257 5859 12291
rect 5859 12257 5868 12291
rect 5816 12248 5868 12257
rect 4620 12180 4672 12232
rect 5172 12180 5224 12232
rect 7012 12223 7064 12232
rect 5356 12112 5408 12164
rect 5540 12112 5592 12164
rect 7012 12189 7021 12223
rect 7021 12189 7055 12223
rect 7055 12189 7064 12223
rect 7012 12180 7064 12189
rect 11520 12248 11572 12300
rect 15660 12248 15712 12300
rect 17960 12384 18012 12436
rect 17500 12359 17552 12368
rect 17500 12325 17509 12359
rect 17509 12325 17543 12359
rect 17543 12325 17552 12359
rect 17500 12316 17552 12325
rect 17776 12316 17828 12368
rect 19524 12427 19576 12436
rect 19524 12393 19533 12427
rect 19533 12393 19567 12427
rect 19567 12393 19576 12427
rect 19524 12384 19576 12393
rect 19984 12427 20036 12436
rect 19984 12393 19993 12427
rect 19993 12393 20027 12427
rect 20027 12393 20036 12427
rect 19984 12384 20036 12393
rect 12440 12223 12492 12232
rect 12440 12189 12449 12223
rect 12449 12189 12483 12223
rect 12483 12189 12492 12223
rect 12440 12180 12492 12189
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 14556 12223 14608 12232
rect 14556 12189 14565 12223
rect 14565 12189 14599 12223
rect 14599 12189 14608 12223
rect 14556 12180 14608 12189
rect 14832 12223 14884 12232
rect 14832 12189 14841 12223
rect 14841 12189 14875 12223
rect 14875 12189 14884 12223
rect 14832 12180 14884 12189
rect 7564 12044 7616 12096
rect 8300 12112 8352 12164
rect 8208 12044 8260 12096
rect 8760 12044 8812 12096
rect 9036 12044 9088 12096
rect 15660 12112 15712 12164
rect 17408 12248 17460 12300
rect 18052 12248 18104 12300
rect 17224 12223 17276 12232
rect 17224 12189 17233 12223
rect 17233 12189 17267 12223
rect 17267 12189 17276 12223
rect 17224 12180 17276 12189
rect 17684 12112 17736 12164
rect 15200 12044 15252 12096
rect 15844 12044 15896 12096
rect 15936 12044 15988 12096
rect 16948 12044 17000 12096
rect 17776 12044 17828 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 18236 12223 18288 12232
rect 18236 12189 18245 12223
rect 18245 12189 18279 12223
rect 18279 12189 18288 12223
rect 18236 12180 18288 12189
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 19984 12248 20036 12300
rect 20260 12248 20312 12300
rect 20628 12248 20680 12300
rect 20352 12223 20404 12232
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 20444 12223 20496 12232
rect 20444 12189 20453 12223
rect 20453 12189 20487 12223
rect 20487 12189 20496 12223
rect 20444 12180 20496 12189
rect 21824 12248 21876 12300
rect 25872 12384 25924 12436
rect 29644 12384 29696 12436
rect 25044 12316 25096 12368
rect 21548 12223 21600 12232
rect 21548 12189 21557 12223
rect 21557 12189 21591 12223
rect 21591 12189 21600 12223
rect 21548 12180 21600 12189
rect 21640 12180 21692 12232
rect 25228 12248 25280 12300
rect 20076 12112 20128 12164
rect 19340 12044 19392 12096
rect 19432 12044 19484 12096
rect 22376 12044 22428 12096
rect 24860 12180 24912 12232
rect 25504 12223 25556 12232
rect 25504 12189 25513 12223
rect 25513 12189 25547 12223
rect 25547 12189 25556 12223
rect 25504 12180 25556 12189
rect 26148 12180 26200 12232
rect 29000 12180 29052 12232
rect 29828 12180 29880 12232
rect 30288 12384 30340 12436
rect 31760 12384 31812 12436
rect 32680 12384 32732 12436
rect 31116 12223 31168 12232
rect 31116 12189 31125 12223
rect 31125 12189 31159 12223
rect 31159 12189 31168 12223
rect 31116 12180 31168 12189
rect 31208 12223 31260 12232
rect 31208 12189 31217 12223
rect 31217 12189 31251 12223
rect 31251 12189 31260 12223
rect 31208 12180 31260 12189
rect 34428 12223 34480 12232
rect 34428 12189 34437 12223
rect 34437 12189 34471 12223
rect 34471 12189 34480 12223
rect 34428 12180 34480 12189
rect 34612 12112 34664 12164
rect 25780 12044 25832 12096
rect 27804 12044 27856 12096
rect 28632 12087 28684 12096
rect 28632 12053 28641 12087
rect 28641 12053 28675 12087
rect 28675 12053 28684 12087
rect 28632 12044 28684 12053
rect 31392 12087 31444 12096
rect 31392 12053 31401 12087
rect 31401 12053 31435 12087
rect 31435 12053 31444 12087
rect 31392 12044 31444 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4620 11883 4672 11892
rect 4620 11849 4629 11883
rect 4629 11849 4663 11883
rect 4663 11849 4672 11883
rect 4620 11840 4672 11849
rect 4988 11840 5040 11892
rect 2872 11772 2924 11824
rect 2136 11747 2188 11756
rect 2136 11713 2145 11747
rect 2145 11713 2179 11747
rect 2179 11713 2188 11747
rect 2136 11704 2188 11713
rect 5356 11772 5408 11824
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 2780 11636 2832 11688
rect 2688 11611 2740 11620
rect 2688 11577 2697 11611
rect 2697 11577 2731 11611
rect 2731 11577 2740 11611
rect 3792 11636 3844 11688
rect 6460 11704 6512 11756
rect 7564 11840 7616 11892
rect 8208 11840 8260 11892
rect 8852 11840 8904 11892
rect 11980 11840 12032 11892
rect 10600 11704 10652 11756
rect 12808 11840 12860 11892
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 13912 11883 13964 11892
rect 13912 11849 13921 11883
rect 13921 11849 13955 11883
rect 13955 11849 13964 11883
rect 13912 11840 13964 11849
rect 15108 11840 15160 11892
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 16120 11840 16172 11892
rect 8116 11679 8168 11688
rect 8116 11645 8125 11679
rect 8125 11645 8159 11679
rect 8159 11645 8168 11679
rect 8116 11636 8168 11645
rect 12992 11747 13044 11756
rect 12992 11713 13001 11747
rect 13001 11713 13035 11747
rect 13035 11713 13044 11747
rect 12992 11704 13044 11713
rect 13912 11704 13964 11756
rect 14832 11815 14884 11824
rect 14832 11781 14841 11815
rect 14841 11781 14875 11815
rect 14875 11781 14884 11815
rect 14832 11772 14884 11781
rect 15200 11704 15252 11756
rect 15292 11704 15344 11756
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 16580 11704 16632 11756
rect 16856 11747 16908 11756
rect 16856 11713 16865 11747
rect 16865 11713 16899 11747
rect 16899 11713 16908 11747
rect 16856 11704 16908 11713
rect 16488 11636 16540 11688
rect 17224 11704 17276 11756
rect 18512 11840 18564 11892
rect 18144 11772 18196 11824
rect 17776 11704 17828 11756
rect 18880 11840 18932 11892
rect 19064 11840 19116 11892
rect 19432 11883 19484 11892
rect 19432 11849 19441 11883
rect 19441 11849 19475 11883
rect 19475 11849 19484 11883
rect 19432 11840 19484 11849
rect 2688 11568 2740 11577
rect 9864 11568 9916 11620
rect 2228 11543 2280 11552
rect 2228 11509 2237 11543
rect 2237 11509 2271 11543
rect 2271 11509 2280 11543
rect 2228 11500 2280 11509
rect 6184 11543 6236 11552
rect 6184 11509 6193 11543
rect 6193 11509 6227 11543
rect 6227 11509 6236 11543
rect 6184 11500 6236 11509
rect 12992 11500 13044 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 17592 11500 17644 11552
rect 18512 11636 18564 11688
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 18972 11568 19024 11620
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 19340 11704 19392 11756
rect 19800 11747 19852 11756
rect 19800 11713 19809 11747
rect 19809 11713 19843 11747
rect 19843 11713 19852 11747
rect 19800 11704 19852 11713
rect 19892 11704 19944 11756
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 20168 11568 20220 11620
rect 20628 11840 20680 11892
rect 20996 11840 21048 11892
rect 21640 11840 21692 11892
rect 23572 11840 23624 11892
rect 24216 11840 24268 11892
rect 24492 11883 24544 11892
rect 24492 11849 24501 11883
rect 24501 11849 24535 11883
rect 24535 11849 24544 11883
rect 24492 11840 24544 11849
rect 24584 11883 24636 11892
rect 24584 11849 24593 11883
rect 24593 11849 24627 11883
rect 24627 11849 24636 11883
rect 24584 11840 24636 11849
rect 25596 11840 25648 11892
rect 29000 11840 29052 11892
rect 20536 11704 20588 11756
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 21180 11747 21232 11756
rect 21180 11713 21189 11747
rect 21189 11713 21223 11747
rect 21223 11713 21232 11747
rect 21180 11704 21232 11713
rect 23112 11772 23164 11824
rect 23664 11636 23716 11688
rect 24124 11747 24176 11756
rect 24124 11713 24133 11747
rect 24133 11713 24167 11747
rect 24167 11713 24176 11747
rect 24124 11704 24176 11713
rect 24400 11704 24452 11756
rect 25136 11704 25188 11756
rect 30104 11772 30156 11824
rect 30656 11772 30708 11824
rect 31208 11772 31260 11824
rect 23020 11568 23072 11620
rect 26056 11636 26108 11688
rect 26516 11704 26568 11756
rect 28080 11704 28132 11756
rect 31116 11704 31168 11756
rect 33048 11840 33100 11892
rect 31760 11747 31812 11756
rect 31760 11713 31769 11747
rect 31769 11713 31803 11747
rect 31803 11713 31812 11747
rect 31760 11704 31812 11713
rect 32496 11747 32548 11756
rect 32496 11713 32505 11747
rect 32505 11713 32539 11747
rect 32539 11713 32548 11747
rect 32496 11704 32548 11713
rect 34520 11747 34572 11756
rect 34520 11713 34529 11747
rect 34529 11713 34563 11747
rect 34563 11713 34572 11747
rect 34520 11704 34572 11713
rect 26792 11636 26844 11688
rect 28632 11636 28684 11688
rect 18788 11500 18840 11552
rect 20076 11500 20128 11552
rect 20904 11500 20956 11552
rect 21272 11500 21324 11552
rect 21824 11500 21876 11552
rect 30564 11679 30616 11688
rect 30564 11645 30573 11679
rect 30573 11645 30607 11679
rect 30607 11645 30616 11679
rect 30564 11636 30616 11645
rect 32772 11679 32824 11688
rect 32772 11645 32781 11679
rect 32781 11645 32815 11679
rect 32815 11645 32824 11679
rect 32772 11636 32824 11645
rect 24216 11500 24268 11552
rect 25044 11500 25096 11552
rect 26148 11543 26200 11552
rect 26148 11509 26157 11543
rect 26157 11509 26191 11543
rect 26191 11509 26200 11543
rect 26148 11500 26200 11509
rect 31668 11611 31720 11620
rect 31668 11577 31677 11611
rect 31677 11577 31711 11611
rect 31711 11577 31720 11611
rect 31668 11568 31720 11577
rect 32864 11500 32916 11552
rect 34244 11543 34296 11552
rect 34244 11509 34253 11543
rect 34253 11509 34287 11543
rect 34287 11509 34296 11543
rect 34244 11500 34296 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2780 11296 2832 11348
rect 5448 11296 5500 11348
rect 6184 11296 6236 11348
rect 12992 11296 13044 11348
rect 3516 11271 3568 11280
rect 3516 11237 3525 11271
rect 3525 11237 3559 11271
rect 3559 11237 3568 11271
rect 3516 11228 3568 11237
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 4988 11228 5040 11280
rect 5356 11160 5408 11212
rect 15752 11339 15804 11348
rect 15752 11305 15761 11339
rect 15761 11305 15795 11339
rect 15795 11305 15804 11339
rect 15752 11296 15804 11305
rect 15936 11296 15988 11348
rect 16488 11296 16540 11348
rect 15844 11228 15896 11280
rect 17684 11296 17736 11348
rect 17868 11296 17920 11348
rect 18052 11296 18104 11348
rect 18880 11296 18932 11348
rect 18512 11228 18564 11280
rect 11152 11160 11204 11212
rect 20444 11296 20496 11348
rect 21180 11296 21232 11348
rect 21548 11296 21600 11348
rect 12624 11092 12676 11144
rect 1584 11024 1636 11076
rect 2228 11024 2280 11076
rect 8668 11024 8720 11076
rect 15660 11024 15712 11076
rect 4160 10956 4212 11008
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 17132 11067 17184 11076
rect 17132 11033 17157 11067
rect 17157 11033 17184 11067
rect 17132 11024 17184 11033
rect 17500 11092 17552 11144
rect 17592 11092 17644 11144
rect 18144 11092 18196 11144
rect 18236 11092 18288 11144
rect 18328 11092 18380 11144
rect 18420 11135 18472 11144
rect 18420 11101 18429 11135
rect 18429 11101 18463 11135
rect 18463 11101 18472 11135
rect 18420 11092 18472 11101
rect 18512 11092 18564 11144
rect 18972 11135 19024 11144
rect 18972 11101 18981 11135
rect 18981 11101 19015 11135
rect 19015 11101 19024 11135
rect 18972 11092 19024 11101
rect 19340 11092 19392 11144
rect 19800 11135 19852 11144
rect 19800 11101 19809 11135
rect 19809 11101 19843 11135
rect 19843 11101 19852 11135
rect 19800 11092 19852 11101
rect 19892 11092 19944 11144
rect 20076 11092 20128 11144
rect 20812 11135 20864 11144
rect 20812 11101 20821 11135
rect 20821 11101 20855 11135
rect 20855 11101 20864 11135
rect 20812 11092 20864 11101
rect 20904 11092 20956 11144
rect 21364 11092 21416 11144
rect 17776 10956 17828 11008
rect 22560 11092 22612 11144
rect 23112 11092 23164 11144
rect 23664 11135 23716 11144
rect 23664 11101 23673 11135
rect 23673 11101 23707 11135
rect 23707 11101 23716 11135
rect 23664 11092 23716 11101
rect 23848 11271 23900 11280
rect 23848 11237 23857 11271
rect 23857 11237 23891 11271
rect 23891 11237 23900 11271
rect 23848 11228 23900 11237
rect 24124 11228 24176 11280
rect 25596 11296 25648 11348
rect 26148 11296 26200 11348
rect 29828 11339 29880 11348
rect 29828 11305 29837 11339
rect 29837 11305 29871 11339
rect 29871 11305 29880 11339
rect 29828 11296 29880 11305
rect 30104 11339 30156 11348
rect 30104 11305 30113 11339
rect 30113 11305 30147 11339
rect 30147 11305 30156 11339
rect 30104 11296 30156 11305
rect 30564 11296 30616 11348
rect 30656 11296 30708 11348
rect 31300 11296 31352 11348
rect 31392 11296 31444 11348
rect 32772 11296 32824 11348
rect 32864 11296 32916 11348
rect 34520 11296 34572 11348
rect 26056 11271 26108 11280
rect 26056 11237 26065 11271
rect 26065 11237 26099 11271
rect 26099 11237 26108 11271
rect 26056 11228 26108 11237
rect 26792 11135 26844 11144
rect 26792 11101 26801 11135
rect 26801 11101 26835 11135
rect 26835 11101 26844 11135
rect 26792 11092 26844 11101
rect 22284 11067 22336 11076
rect 22284 11033 22293 11067
rect 22293 11033 22327 11067
rect 22327 11033 22336 11067
rect 22284 11024 22336 11033
rect 24216 11024 24268 11076
rect 27804 11024 27856 11076
rect 30840 11203 30892 11212
rect 30840 11169 30849 11203
rect 30849 11169 30883 11203
rect 30883 11169 30892 11203
rect 32496 11228 32548 11280
rect 30840 11160 30892 11169
rect 31116 11092 31168 11144
rect 31668 11092 31720 11144
rect 34428 11160 34480 11212
rect 30656 11024 30708 11076
rect 18788 10956 18840 11008
rect 20352 10956 20404 11008
rect 21732 10999 21784 11008
rect 21732 10965 21741 10999
rect 21741 10965 21775 10999
rect 21775 10965 21784 10999
rect 21732 10956 21784 10965
rect 28080 10956 28132 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1676 10752 1728 10804
rect 5540 10752 5592 10804
rect 6000 10752 6052 10804
rect 6460 10752 6512 10804
rect 4160 10684 4212 10736
rect 8668 10727 8720 10736
rect 8668 10693 8677 10727
rect 8677 10693 8711 10727
rect 8711 10693 8720 10727
rect 8668 10684 8720 10693
rect 9036 10684 9088 10736
rect 16672 10684 16724 10736
rect 17316 10684 17368 10736
rect 17592 10684 17644 10736
rect 18512 10684 18564 10736
rect 940 10616 992 10668
rect 1400 10480 1452 10532
rect 2780 10480 2832 10532
rect 3148 10591 3200 10600
rect 3148 10557 3157 10591
rect 3157 10557 3191 10591
rect 3191 10557 3200 10591
rect 3148 10548 3200 10557
rect 3884 10548 3936 10600
rect 17132 10616 17184 10668
rect 17500 10616 17552 10668
rect 17776 10659 17828 10668
rect 17776 10625 17785 10659
rect 17785 10625 17819 10659
rect 17819 10625 17828 10659
rect 17776 10616 17828 10625
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 10692 10480 10744 10532
rect 12716 10480 12768 10532
rect 17776 10480 17828 10532
rect 19248 10480 19300 10532
rect 20904 10752 20956 10804
rect 24308 10752 24360 10804
rect 31116 10752 31168 10804
rect 31760 10795 31812 10804
rect 20996 10727 21048 10736
rect 20996 10693 21005 10727
rect 21005 10693 21039 10727
rect 21039 10693 21048 10727
rect 20996 10684 21048 10693
rect 21272 10727 21324 10736
rect 21272 10693 21281 10727
rect 21281 10693 21315 10727
rect 21315 10693 21324 10727
rect 21272 10684 21324 10693
rect 21364 10684 21416 10736
rect 22928 10727 22980 10736
rect 22928 10693 22937 10727
rect 22937 10693 22971 10727
rect 22971 10693 22980 10727
rect 22928 10684 22980 10693
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22284 10616 22336 10625
rect 22560 10659 22612 10668
rect 22560 10625 22569 10659
rect 22569 10625 22603 10659
rect 22603 10625 22612 10659
rect 22560 10616 22612 10625
rect 22652 10659 22704 10668
rect 22652 10625 22661 10659
rect 22661 10625 22695 10659
rect 22695 10625 22704 10659
rect 22652 10616 22704 10625
rect 23112 10616 23164 10668
rect 23480 10659 23532 10668
rect 23480 10625 23489 10659
rect 23489 10625 23523 10659
rect 23523 10625 23532 10659
rect 23480 10616 23532 10625
rect 24216 10659 24268 10668
rect 24216 10625 24225 10659
rect 24225 10625 24259 10659
rect 24259 10625 24268 10659
rect 24216 10616 24268 10625
rect 24400 10616 24452 10668
rect 30656 10616 30708 10668
rect 31760 10761 31769 10795
rect 31769 10761 31803 10795
rect 31803 10761 31812 10795
rect 31760 10752 31812 10761
rect 34520 10795 34572 10804
rect 34520 10761 34529 10795
rect 34529 10761 34563 10795
rect 34563 10761 34572 10795
rect 34520 10752 34572 10761
rect 20812 10412 20864 10464
rect 32404 10480 32456 10532
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 2780 10208 2832 10260
rect 3884 10208 3936 10260
rect 1400 10115 1452 10124
rect 1400 10081 1409 10115
rect 1409 10081 1443 10115
rect 1443 10081 1452 10115
rect 1400 10072 1452 10081
rect 2780 10004 2832 10056
rect 15660 10047 15712 10056
rect 15660 10013 15669 10047
rect 15669 10013 15703 10047
rect 15703 10013 15712 10047
rect 15660 10004 15712 10013
rect 17224 10251 17276 10260
rect 17224 10217 17233 10251
rect 17233 10217 17267 10251
rect 17267 10217 17276 10251
rect 17224 10208 17276 10217
rect 17500 10208 17552 10260
rect 18328 10208 18380 10260
rect 22100 10208 22152 10260
rect 23480 10208 23532 10260
rect 16488 10004 16540 10056
rect 16580 10047 16632 10056
rect 16580 10013 16589 10047
rect 16589 10013 16623 10047
rect 16623 10013 16632 10047
rect 16580 10004 16632 10013
rect 16672 10047 16724 10056
rect 16672 10013 16681 10047
rect 16681 10013 16715 10047
rect 16715 10013 16724 10047
rect 16672 10004 16724 10013
rect 17224 10072 17276 10124
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 17040 10004 17092 10056
rect 17500 10004 17552 10056
rect 17684 10004 17736 10056
rect 17868 10004 17920 10056
rect 20812 10140 20864 10192
rect 20444 10115 20496 10124
rect 20444 10081 20453 10115
rect 20453 10081 20487 10115
rect 20487 10081 20496 10115
rect 20444 10072 20496 10081
rect 20996 10072 21048 10124
rect 21732 10072 21784 10124
rect 18328 10047 18380 10056
rect 18328 10013 18337 10047
rect 18337 10013 18371 10047
rect 18371 10013 18380 10047
rect 18328 10004 18380 10013
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 19984 10004 20036 10056
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 21272 10004 21324 10056
rect 22652 10004 22704 10056
rect 27528 10004 27580 10056
rect 28080 10047 28132 10056
rect 28080 10013 28089 10047
rect 28089 10013 28123 10047
rect 28123 10013 28132 10047
rect 28080 10004 28132 10013
rect 31116 10004 31168 10056
rect 17684 9911 17736 9920
rect 17684 9877 17693 9911
rect 17693 9877 17727 9911
rect 17727 9877 17736 9911
rect 17684 9868 17736 9877
rect 17776 9868 17828 9920
rect 34428 10047 34480 10056
rect 34428 10013 34437 10047
rect 34437 10013 34471 10047
rect 34471 10013 34480 10047
rect 34428 10004 34480 10013
rect 32312 9868 32364 9920
rect 33140 9868 33192 9920
rect 34060 9936 34112 9988
rect 34152 9868 34204 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2780 9664 2832 9716
rect 16672 9596 16724 9648
rect 18420 9664 18472 9716
rect 18328 9596 18380 9648
rect 2688 9528 2740 9580
rect 16488 9528 16540 9580
rect 17224 9571 17276 9580
rect 17224 9537 17233 9571
rect 17233 9537 17267 9571
rect 17267 9537 17276 9571
rect 17224 9528 17276 9537
rect 17868 9571 17920 9580
rect 15660 9460 15712 9512
rect 17684 9503 17736 9512
rect 17684 9469 17693 9503
rect 17693 9469 17727 9503
rect 17727 9469 17736 9503
rect 17684 9460 17736 9469
rect 17868 9537 17897 9571
rect 17897 9537 17920 9571
rect 17868 9528 17920 9537
rect 18144 9460 18196 9512
rect 20996 9596 21048 9648
rect 32404 9639 32456 9648
rect 32404 9605 32413 9639
rect 32413 9605 32447 9639
rect 32447 9605 32456 9639
rect 32404 9596 32456 9605
rect 33140 9596 33192 9648
rect 19432 9571 19484 9580
rect 19432 9537 19441 9571
rect 19441 9537 19475 9571
rect 19475 9537 19484 9571
rect 19432 9528 19484 9537
rect 27344 9528 27396 9580
rect 27528 9528 27580 9580
rect 34152 9571 34204 9580
rect 34152 9537 34161 9571
rect 34161 9537 34195 9571
rect 34195 9537 34204 9571
rect 34152 9528 34204 9537
rect 16580 9324 16632 9376
rect 32036 9460 32088 9512
rect 32496 9460 32548 9512
rect 18604 9324 18656 9376
rect 33876 9367 33928 9376
rect 33876 9333 33885 9367
rect 33885 9333 33919 9367
rect 33919 9333 33928 9367
rect 33876 9324 33928 9333
rect 34060 9367 34112 9376
rect 34060 9333 34069 9367
rect 34069 9333 34103 9367
rect 34103 9333 34112 9367
rect 34060 9324 34112 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2872 9120 2924 9172
rect 16672 9120 16724 9172
rect 17868 9120 17920 9172
rect 18604 9120 18656 9172
rect 19984 9120 20036 9172
rect 32036 9163 32088 9172
rect 32036 9129 32045 9163
rect 32045 9129 32079 9163
rect 32079 9129 32088 9163
rect 32036 9120 32088 9129
rect 940 8916 992 8968
rect 16580 8916 16632 8968
rect 19432 9052 19484 9104
rect 34060 8916 34112 8968
rect 32312 8848 32364 8900
rect 33324 8780 33376 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 34244 7828 34296 7880
rect 34612 7760 34664 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 940 6740 992 6792
rect 1584 6647 1636 6656
rect 1584 6613 1593 6647
rect 1593 6613 1627 6647
rect 1627 6613 1636 6647
rect 1584 6604 1636 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 33876 5652 33928 5704
rect 34336 5627 34388 5636
rect 34336 5593 34345 5627
rect 34345 5593 34379 5627
rect 34379 5593 34388 5627
rect 34336 5584 34388 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2964 4768 3016 4820
rect 940 4564 992 4616
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 33324 3519 33376 3528
rect 33324 3485 33333 3519
rect 33333 3485 33367 3519
rect 33367 3485 33376 3519
rect 33324 3476 33376 3485
rect 34888 3408 34940 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 1492 2592 1544 2644
rect 27344 2635 27396 2644
rect 27344 2601 27353 2635
rect 27353 2601 27387 2635
rect 27387 2601 27396 2635
rect 27344 2592 27396 2601
rect 9036 2456 9088 2508
rect 940 2388 992 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 27252 2388 27304 2440
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 952 36174 980 36751
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 940 36168 992 36174
rect 940 36110 992 36116
rect 33876 36168 33928 36174
rect 33876 36110 33928 36116
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1596 35894 1624 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 1596 35866 1808 35894
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 940 35080 992 35086
rect 940 35022 992 35028
rect 952 34649 980 35022
rect 938 34640 994 34649
rect 938 34575 994 34584
rect 940 32904 992 32910
rect 940 32846 992 32852
rect 952 32473 980 32846
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 938 32464 994 32473
rect 938 32399 994 32408
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30297 1440 30670
rect 1398 30288 1454 30297
rect 1398 30223 1454 30232
rect 1596 29458 1624 32710
rect 1504 29430 1624 29458
rect 940 28552 992 28558
rect 940 28494 992 28500
rect 952 28121 980 28494
rect 938 28112 994 28121
rect 938 28047 994 28056
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 26217 1440 26318
rect 1398 26208 1454 26217
rect 1398 26143 1454 26152
rect 940 24200 992 24206
rect 940 24142 992 24148
rect 952 23769 980 24142
rect 938 23760 994 23769
rect 938 23695 994 23704
rect 1400 23656 1452 23662
rect 1400 23598 1452 23604
rect 1412 23118 1440 23598
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1504 23066 1532 29430
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1596 26234 1624 28358
rect 1596 26206 1716 26234
rect 1688 23186 1716 26206
rect 1676 23180 1728 23186
rect 1676 23122 1728 23128
rect 1504 23038 1716 23066
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21593 980 21966
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1596 21690 1624 21830
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 20942 1440 21422
rect 1688 21010 1716 23038
rect 1676 21004 1728 21010
rect 1676 20946 1728 20952
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 940 19848 992 19854
rect 940 19790 992 19796
rect 952 19417 980 19790
rect 1412 19718 1440 20878
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 938 19408 994 19417
rect 1412 19378 1440 19654
rect 938 19343 994 19352
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1688 17746 1716 19654
rect 1780 19310 1808 35866
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 2872 34944 2924 34950
rect 2872 34886 2924 34892
rect 1860 26240 1912 26246
rect 1860 26182 1912 26188
rect 1872 23798 1900 26182
rect 2044 24064 2096 24070
rect 2044 24006 2096 24012
rect 1860 23792 1912 23798
rect 1860 23734 1912 23740
rect 2056 19922 2084 24006
rect 2228 23044 2280 23050
rect 2228 22986 2280 22992
rect 2240 22778 2268 22986
rect 2596 22976 2648 22982
rect 2596 22918 2648 22924
rect 2228 22772 2280 22778
rect 2228 22714 2280 22720
rect 2608 22574 2636 22918
rect 2884 22710 2912 34886
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 3700 30592 3752 30598
rect 3700 30534 3752 30540
rect 33140 30592 33192 30598
rect 33140 30534 33192 30540
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 3424 24064 3476 24070
rect 3424 24006 3476 24012
rect 2976 23730 3004 24006
rect 3436 23730 3464 24006
rect 3712 23798 3740 30534
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 33152 30326 33180 30534
rect 29276 30320 29328 30326
rect 29276 30262 29328 30268
rect 33140 30320 33192 30326
rect 33140 30262 33192 30268
rect 28816 30184 28868 30190
rect 28816 30126 28868 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 28828 29850 28856 30126
rect 29288 29850 29316 30262
rect 31852 30252 31904 30258
rect 31852 30194 31904 30200
rect 31024 30184 31076 30190
rect 31024 30126 31076 30132
rect 29828 30048 29880 30054
rect 29828 29990 29880 29996
rect 28816 29844 28868 29850
rect 28816 29786 28868 29792
rect 29276 29844 29328 29850
rect 29276 29786 29328 29792
rect 29840 29714 29868 29990
rect 25136 29708 25188 29714
rect 25136 29650 25188 29656
rect 29828 29708 29880 29714
rect 29828 29650 29880 29656
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 24676 29572 24728 29578
rect 24676 29514 24728 29520
rect 23388 29504 23440 29510
rect 23388 29446 23440 29452
rect 24308 29504 24360 29510
rect 24308 29446 24360 29452
rect 24400 29504 24452 29510
rect 24400 29446 24452 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 23400 29186 23428 29446
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 23400 29170 23612 29186
rect 23400 29164 23624 29170
rect 23400 29158 23572 29164
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 21364 27668 21416 27674
rect 21364 27610 21416 27616
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19432 27464 19484 27470
rect 19432 27406 19484 27412
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 20076 27464 20128 27470
rect 20076 27406 20128 27412
rect 18972 27396 19024 27402
rect 18972 27338 19024 27344
rect 17592 27328 17644 27334
rect 17592 27270 17644 27276
rect 17604 27130 17632 27270
rect 18984 27130 19012 27338
rect 19260 27130 19288 27406
rect 17592 27124 17644 27130
rect 17592 27066 17644 27072
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 13360 26988 13412 26994
rect 13360 26930 13412 26936
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 13176 26920 13228 26926
rect 13176 26862 13228 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 13188 26586 13216 26862
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13268 26512 13320 26518
rect 13268 26454 13320 26460
rect 11980 26376 12032 26382
rect 11980 26318 12032 26324
rect 12992 26376 13044 26382
rect 12992 26318 13044 26324
rect 13084 26376 13136 26382
rect 13084 26318 13136 26324
rect 11060 26308 11112 26314
rect 11060 26250 11112 26256
rect 9496 26240 9548 26246
rect 9496 26182 9548 26188
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 8852 25696 8904 25702
rect 8852 25638 8904 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 8864 25158 8892 25638
rect 9416 25294 9444 25842
rect 9508 25702 9536 26182
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 9496 25696 9548 25702
rect 9496 25638 9548 25644
rect 9864 25696 9916 25702
rect 9864 25638 9916 25644
rect 9508 25294 9536 25638
rect 9680 25424 9732 25430
rect 9680 25366 9732 25372
rect 9404 25288 9456 25294
rect 9404 25230 9456 25236
rect 9496 25288 9548 25294
rect 9496 25230 9548 25236
rect 9036 25220 9088 25226
rect 9036 25162 9088 25168
rect 8852 25152 8904 25158
rect 8852 25094 8904 25100
rect 8864 24886 8892 25094
rect 8852 24880 8904 24886
rect 8852 24822 8904 24828
rect 9048 24818 9076 25162
rect 9416 24954 9444 25230
rect 9404 24948 9456 24954
rect 9404 24890 9456 24896
rect 8576 24812 8628 24818
rect 8576 24754 8628 24760
rect 9036 24812 9088 24818
rect 9036 24754 9088 24760
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 8588 24698 8616 24754
rect 8588 24682 8892 24698
rect 8588 24676 8904 24682
rect 8588 24670 8852 24676
rect 8852 24618 8904 24624
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 2964 23724 3016 23730
rect 2964 23666 3016 23672
rect 3424 23724 3476 23730
rect 3424 23666 3476 23672
rect 3436 23322 3464 23666
rect 3424 23316 3476 23322
rect 3424 23258 3476 23264
rect 4080 23202 4108 24142
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6656 23798 6684 24006
rect 4712 23792 4764 23798
rect 4712 23734 4764 23740
rect 6644 23792 6696 23798
rect 6644 23734 6696 23740
rect 8300 23792 8352 23798
rect 8300 23734 8352 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4724 23322 4752 23734
rect 5356 23656 5408 23662
rect 5356 23598 5408 23604
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 4712 23316 4764 23322
rect 4712 23258 4764 23264
rect 4160 23248 4212 23254
rect 4080 23196 4160 23202
rect 4080 23190 4212 23196
rect 4080 23174 4200 23190
rect 2872 22704 2924 22710
rect 2872 22646 2924 22652
rect 3884 22704 3936 22710
rect 3884 22646 3936 22652
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2608 21486 2636 22510
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2700 21894 2728 22374
rect 3896 22234 3924 22646
rect 3884 22228 3936 22234
rect 3884 22170 3936 22176
rect 4080 22030 4108 23174
rect 4816 23118 4844 23462
rect 4804 23112 4856 23118
rect 4804 23054 4856 23060
rect 4712 23044 4764 23050
rect 4712 22986 4764 22992
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 4620 21888 4672 21894
rect 4620 21830 4672 21836
rect 2700 21554 2728 21830
rect 4632 21690 4660 21830
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2700 21350 2728 21490
rect 3148 21480 3200 21486
rect 3148 21422 3200 21428
rect 2228 21344 2280 21350
rect 2228 21286 2280 21292
rect 2688 21344 2740 21350
rect 2688 21286 2740 21292
rect 2872 21344 2924 21350
rect 2872 21286 2924 21292
rect 2240 20874 2268 21286
rect 2228 20868 2280 20874
rect 2228 20810 2280 20816
rect 2884 20262 2912 21286
rect 3160 21146 3188 21422
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 3056 20256 3108 20262
rect 3056 20198 3108 20204
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 2332 19446 2360 20198
rect 2320 19440 2372 19446
rect 2320 19382 2372 19388
rect 1768 19304 1820 19310
rect 1768 19246 1820 19252
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 2320 17604 2372 17610
rect 2320 17546 2372 17552
rect 2332 17338 2360 17546
rect 2320 17332 2372 17338
rect 2320 17274 2372 17280
rect 938 17232 994 17241
rect 2884 17202 2912 20198
rect 3068 19854 3096 20198
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4724 20058 4752 22986
rect 4804 22568 4856 22574
rect 4804 22510 4856 22516
rect 4816 21010 4844 22510
rect 4896 22432 4948 22438
rect 4896 22374 4948 22380
rect 4908 22234 4936 22374
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 5184 22094 5212 23462
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5276 22234 5304 23122
rect 5264 22228 5316 22234
rect 5264 22170 5316 22176
rect 5184 22066 5304 22094
rect 5172 21888 5224 21894
rect 5172 21830 5224 21836
rect 4988 21616 5040 21622
rect 4986 21584 4988 21593
rect 5040 21584 5042 21593
rect 4896 21548 4948 21554
rect 5184 21554 5212 21830
rect 5276 21554 5304 22066
rect 5368 22030 5396 23598
rect 6656 23186 6684 23734
rect 8312 23322 8340 23734
rect 8864 23322 8892 24618
rect 9048 24206 9076 24754
rect 9232 24410 9260 24754
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 8300 23316 8352 23322
rect 8300 23258 8352 23264
rect 8852 23316 8904 23322
rect 8852 23258 8904 23264
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 5448 23112 5500 23118
rect 5448 23054 5500 23060
rect 5460 22234 5488 23054
rect 6656 22438 6684 23122
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 7656 23044 7708 23050
rect 7656 22986 7708 22992
rect 7668 22778 7696 22986
rect 8220 22778 8248 23054
rect 7656 22772 7708 22778
rect 7656 22714 7708 22720
rect 8208 22772 8260 22778
rect 8208 22714 8260 22720
rect 6644 22432 6696 22438
rect 6644 22374 6696 22380
rect 5448 22228 5500 22234
rect 5448 22170 5500 22176
rect 5448 22092 5500 22098
rect 6656 22094 6684 22374
rect 8220 22094 8248 22714
rect 9312 22432 9364 22438
rect 9312 22374 9364 22380
rect 5448 22034 5500 22040
rect 6472 22066 6684 22094
rect 8036 22066 8248 22094
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 5460 21706 5488 22034
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 5368 21678 5488 21706
rect 5368 21554 5396 21678
rect 5736 21554 5764 21966
rect 5920 21690 5948 21966
rect 5908 21684 5960 21690
rect 5908 21626 5960 21632
rect 5816 21616 5868 21622
rect 5814 21584 5816 21593
rect 5868 21584 5870 21593
rect 4986 21519 5042 21528
rect 5172 21548 5224 21554
rect 4896 21490 4948 21496
rect 5172 21490 5224 21496
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5356 21548 5408 21554
rect 5724 21548 5776 21554
rect 5356 21490 5408 21496
rect 5460 21508 5724 21536
rect 4908 21146 4936 21490
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 4988 21344 5040 21350
rect 4988 21286 5040 21292
rect 4896 21140 4948 21146
rect 4896 21082 4948 21088
rect 4804 21004 4856 21010
rect 4804 20946 4856 20952
rect 4712 20052 4764 20058
rect 4712 19994 4764 20000
rect 4436 19984 4488 19990
rect 4436 19926 4488 19932
rect 4252 19916 4304 19922
rect 4252 19858 4304 19864
rect 3056 19848 3108 19854
rect 3056 19790 3108 19796
rect 4160 19712 4212 19718
rect 4160 19654 4212 19660
rect 4172 19446 4200 19654
rect 4264 19514 4292 19858
rect 4252 19508 4304 19514
rect 4252 19450 4304 19456
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4448 19174 4476 19926
rect 4816 19666 4844 20946
rect 5000 19922 5028 21286
rect 4988 19916 5040 19922
rect 4988 19858 5040 19864
rect 4632 19638 4844 19666
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 3056 19168 3108 19174
rect 3056 19110 3108 19116
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 4436 19168 4488 19174
rect 4436 19110 4488 19116
rect 3068 18630 3096 19110
rect 3436 18766 3464 19110
rect 3988 18834 4016 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4632 18850 4660 19638
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4724 18970 4752 19450
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4712 18964 4764 18970
rect 4712 18906 4764 18912
rect 3976 18828 4028 18834
rect 4632 18822 4752 18850
rect 3976 18770 4028 18776
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3056 18624 3108 18630
rect 3056 18566 3108 18572
rect 3068 17610 3096 18566
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 3160 17338 3188 17478
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 938 17167 940 17176
rect 992 17167 994 17176
rect 2872 17196 2924 17202
rect 940 17138 992 17144
rect 2872 17138 2924 17144
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 1860 15428 1912 15434
rect 1860 15370 1912 15376
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 938 15056 994 15065
rect 938 14991 940 15000
rect 992 14991 994 15000
rect 940 14962 992 14968
rect 1688 13394 1716 15302
rect 1872 15162 1900 15370
rect 1860 15156 1912 15162
rect 1860 15098 1912 15104
rect 2884 14006 2912 17002
rect 3332 16108 3384 16114
rect 3332 16050 3384 16056
rect 3344 15706 3372 16050
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3436 14804 3464 17478
rect 4172 17202 4200 17478
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 3516 17128 3568 17134
rect 3516 17070 3568 17076
rect 3976 17128 4028 17134
rect 3976 17070 4028 17076
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3528 16794 3556 17070
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3516 16788 3568 16794
rect 3516 16730 3568 16736
rect 3620 15502 3648 16934
rect 3988 16590 4016 17070
rect 4080 16726 4108 17070
rect 4632 16998 4660 17138
rect 4620 16992 4672 16998
rect 4620 16934 4672 16940
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16720 4120 16726
rect 4068 16662 4120 16668
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 16182 4016 16526
rect 3976 16176 4028 16182
rect 3976 16118 4028 16124
rect 3608 15496 3660 15502
rect 3608 15438 3660 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3516 14816 3568 14822
rect 3436 14776 3516 14804
rect 3516 14758 3568 14764
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 3528 13870 3556 14758
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 1676 13388 1728 13394
rect 1676 13330 1728 13336
rect 1676 13252 1728 13258
rect 1676 13194 1728 13200
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 938 12880 994 12889
rect 938 12815 940 12824
rect 992 12815 994 12824
rect 940 12786 992 12792
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 938 10704 994 10713
rect 938 10639 940 10648
rect 992 10639 994 10648
rect 940 10610 992 10616
rect 1412 10538 1440 11086
rect 1584 11076 1636 11082
rect 1584 11018 1636 11024
rect 1400 10532 1452 10538
rect 1400 10474 1452 10480
rect 1412 10130 1440 10474
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 952 8537 980 8910
rect 1596 8650 1624 11018
rect 1688 10810 1716 13194
rect 2332 12986 2360 13194
rect 3528 13190 3556 13806
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 3528 12646 3556 13126
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 2148 11762 2176 12582
rect 3528 12442 3556 12582
rect 3516 12436 3568 12442
rect 3516 12378 3568 12384
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2780 11688 2832 11694
rect 2780 11630 2832 11636
rect 2688 11620 2740 11626
rect 2688 11562 2740 11568
rect 2228 11552 2280 11558
rect 2228 11494 2280 11500
rect 2240 11082 2268 11494
rect 2228 11076 2280 11082
rect 2228 11018 2280 11024
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1676 9988 1728 9994
rect 1676 9930 1728 9936
rect 1504 8622 1624 8650
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 952 6361 980 6734
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1504 2650 1532 8622
rect 1688 6914 1716 9930
rect 2700 9586 2728 11562
rect 2792 11354 2820 11630
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2792 10538 2820 11290
rect 2780 10532 2832 10538
rect 2780 10474 2832 10480
rect 2792 10266 2820 10474
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9722 2820 9998
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2688 9580 2740 9586
rect 2688 9522 2740 9528
rect 2884 9178 2912 11766
rect 3528 11286 3556 12378
rect 3804 11694 3832 15302
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 14006 3924 14214
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3988 12434 4016 16118
rect 4080 16114 4108 16662
rect 4632 16590 4660 16934
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 4632 15978 4660 16526
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 15914
rect 4724 15502 4752 18822
rect 4816 18290 4844 19246
rect 4908 18970 4936 19654
rect 5000 19446 5028 19654
rect 4988 19440 5040 19446
rect 4988 19382 5040 19388
rect 4988 19168 5040 19174
rect 4988 19110 5040 19116
rect 4896 18964 4948 18970
rect 4896 18906 4948 18912
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4908 17610 4936 18566
rect 5000 18290 5028 19110
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 4804 15904 4856 15910
rect 4804 15846 4856 15852
rect 4816 15706 4844 15846
rect 4804 15700 4856 15706
rect 4804 15642 4856 15648
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4908 15366 4936 17546
rect 5000 17338 5028 18226
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 5000 16114 5028 16526
rect 4988 16108 5040 16114
rect 4988 16050 5040 16056
rect 5092 15706 5120 21354
rect 5356 21140 5408 21146
rect 5356 21082 5408 21088
rect 5264 20800 5316 20806
rect 5264 20742 5316 20748
rect 5276 19854 5304 20742
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5184 19514 5212 19790
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5276 19378 5304 19790
rect 5264 19372 5316 19378
rect 5264 19314 5316 19320
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 18630 5212 19246
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5172 18624 5224 18630
rect 5172 18566 5224 18572
rect 5184 17882 5212 18566
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 5276 17746 5304 19110
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5368 17626 5396 21082
rect 5460 20777 5488 21508
rect 5814 21519 5870 21528
rect 5724 21490 5776 21496
rect 6472 21486 6500 22066
rect 8036 22030 8064 22066
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 9324 21962 9352 22374
rect 9312 21956 9364 21962
rect 9312 21898 9364 21904
rect 7656 21888 7708 21894
rect 7656 21830 7708 21836
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 8024 21888 8076 21894
rect 8024 21830 8076 21836
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6368 21412 6420 21418
rect 6368 21354 6420 21360
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6380 21010 6408 21354
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6368 21004 6420 21010
rect 6368 20946 6420 20952
rect 6564 20942 6592 21286
rect 6656 21146 6684 21354
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 21146 6776 21286
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 6736 21140 6788 21146
rect 6736 21082 6788 21088
rect 6840 21026 6868 21422
rect 6748 20998 6868 21026
rect 6748 20942 6776 20998
rect 6552 20936 6604 20942
rect 6552 20878 6604 20884
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6748 20806 6776 20878
rect 6736 20800 6788 20806
rect 5446 20768 5502 20777
rect 6736 20742 6788 20748
rect 5446 20703 5502 20712
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5460 19174 5488 19858
rect 6748 19446 6776 20742
rect 7668 19854 7696 21830
rect 7760 20874 7788 21830
rect 8036 21622 8064 21830
rect 9324 21690 9352 21898
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 8024 21616 8076 21622
rect 8024 21558 8076 21564
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8864 21146 8892 21490
rect 8852 21140 8904 21146
rect 8852 21082 8904 21088
rect 7748 20868 7800 20874
rect 7748 20810 7800 20816
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20262 8984 20742
rect 8944 20256 8996 20262
rect 8944 20198 8996 20204
rect 8956 19922 8984 20198
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 8576 19848 8628 19854
rect 8576 19790 8628 19796
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 5632 19304 5684 19310
rect 5632 19246 5684 19252
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5644 18970 5672 19246
rect 5632 18964 5684 18970
rect 5632 18906 5684 18912
rect 6564 18766 6592 19314
rect 6552 18760 6604 18766
rect 6552 18702 6604 18708
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5460 18290 5488 18566
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5276 17598 5396 17626
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 4804 14340 4856 14346
rect 4804 14282 4856 14288
rect 4816 14074 4844 14282
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4816 13530 4844 14010
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4908 13394 4936 13670
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5000 12918 5028 14554
rect 5092 14278 5120 15642
rect 5276 15314 5304 17598
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5368 17338 5396 17478
rect 5356 17332 5408 17338
rect 5356 17274 5408 17280
rect 5460 16182 5488 18226
rect 6564 17882 6592 18702
rect 7576 18698 7604 19654
rect 8496 19310 8524 19654
rect 8588 19514 8616 19790
rect 8760 19712 8812 19718
rect 8760 19654 8812 19660
rect 8576 19508 8628 19514
rect 8576 19450 8628 19456
rect 8772 19446 8800 19654
rect 8760 19440 8812 19446
rect 8760 19382 8812 19388
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8312 18766 8340 19110
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 8496 18630 8524 19246
rect 8956 19174 8984 19858
rect 9036 19780 9088 19786
rect 9036 19722 9088 19728
rect 8944 19168 8996 19174
rect 8944 19110 8996 19116
rect 8484 18624 8536 18630
rect 8484 18566 8536 18572
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8312 17882 8340 18090
rect 8496 18086 8524 18566
rect 8956 18086 8984 19110
rect 9048 18970 9076 19722
rect 9036 18964 9088 18970
rect 9036 18906 9088 18912
rect 8484 18080 8536 18086
rect 8484 18022 8536 18028
rect 8944 18080 8996 18086
rect 8944 18022 8996 18028
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 6368 17740 6420 17746
rect 6368 17682 6420 17688
rect 6380 17202 6408 17682
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6748 17338 6776 17546
rect 8496 17542 8524 18022
rect 8956 17678 8984 18022
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8220 17338 8248 17478
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 7392 16794 7420 17206
rect 8496 17066 8524 17478
rect 9416 17270 9444 24890
rect 9508 22438 9536 25230
rect 9692 22642 9720 25366
rect 9876 25362 9904 25638
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 10244 25294 10272 25842
rect 11072 25294 11100 26250
rect 11992 25974 12020 26318
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 11980 25968 12032 25974
rect 11334 25936 11390 25945
rect 11980 25910 12032 25916
rect 11334 25871 11336 25880
rect 11388 25871 11390 25880
rect 11336 25842 11388 25848
rect 11704 25832 11756 25838
rect 11704 25774 11756 25780
rect 11888 25832 11940 25838
rect 11888 25774 11940 25780
rect 11716 25430 11744 25774
rect 11704 25424 11756 25430
rect 11704 25366 11756 25372
rect 11900 25362 11928 25774
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 10232 25288 10284 25294
rect 10232 25230 10284 25236
rect 11060 25288 11112 25294
rect 11704 25288 11756 25294
rect 11112 25248 11192 25276
rect 11060 25230 11112 25236
rect 10416 25220 10468 25226
rect 10416 25162 10468 25168
rect 10876 25220 10928 25226
rect 10876 25162 10928 25168
rect 10428 24274 10456 25162
rect 10508 25152 10560 25158
rect 10508 25094 10560 25100
rect 10416 24268 10468 24274
rect 10416 24210 10468 24216
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 23118 10272 23462
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 10060 22506 10088 23054
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10048 22500 10100 22506
rect 10048 22442 10100 22448
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9508 21894 9536 22374
rect 9784 22098 9812 22374
rect 9772 22092 9824 22098
rect 9772 22034 9824 22040
rect 9680 22024 9732 22030
rect 9600 21984 9680 22012
rect 9600 21894 9628 21984
rect 10060 22012 10088 22442
rect 10232 22024 10284 22030
rect 10060 21984 10232 22012
rect 9680 21966 9732 21972
rect 10232 21966 10284 21972
rect 9496 21888 9548 21894
rect 9496 21830 9548 21836
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 10140 21888 10192 21894
rect 10140 21830 10192 21836
rect 9508 21486 9536 21830
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9508 20602 9536 21422
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9496 20256 9548 20262
rect 10152 20244 10180 21830
rect 10244 21554 10272 21966
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 10336 21486 10364 22578
rect 10520 21690 10548 25094
rect 10888 24698 10916 25162
rect 10888 24682 11100 24698
rect 10888 24676 11112 24682
rect 10888 24670 11060 24676
rect 11060 24618 11112 24624
rect 10784 24608 10836 24614
rect 10784 24550 10836 24556
rect 10692 24268 10744 24274
rect 10692 24210 10744 24216
rect 10704 24138 10732 24210
rect 10796 24188 10824 24550
rect 11164 24410 11192 25248
rect 11704 25230 11756 25236
rect 11336 25220 11388 25226
rect 11336 25162 11388 25168
rect 11244 25152 11296 25158
rect 11244 25094 11296 25100
rect 11152 24404 11204 24410
rect 11152 24346 11204 24352
rect 11060 24200 11112 24206
rect 10796 24160 11060 24188
rect 10692 24132 10744 24138
rect 10692 24074 10744 24080
rect 10980 23798 11008 24160
rect 11060 24142 11112 24148
rect 10968 23792 11020 23798
rect 10968 23734 11020 23740
rect 10600 23724 10652 23730
rect 10600 23666 10652 23672
rect 10612 23526 10640 23666
rect 10600 23520 10652 23526
rect 10600 23462 10652 23468
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 10612 22438 10640 23462
rect 10796 22506 10824 23462
rect 10784 22500 10836 22506
rect 10784 22442 10836 22448
rect 10600 22432 10652 22438
rect 10600 22374 10652 22380
rect 10980 22166 11008 23734
rect 11164 23050 11192 24346
rect 11256 24206 11284 25094
rect 11348 24954 11376 25162
rect 11716 24954 11744 25230
rect 11336 24948 11388 24954
rect 11336 24890 11388 24896
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11716 23866 11744 24890
rect 11888 24336 11940 24342
rect 11888 24278 11940 24284
rect 11900 24206 11928 24278
rect 11888 24200 11940 24206
rect 11888 24142 11940 24148
rect 11992 24070 12020 25910
rect 12544 25906 12572 26250
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 12256 25152 12308 25158
rect 12256 25094 12308 25100
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12084 24342 12112 25094
rect 12072 24336 12124 24342
rect 12124 24296 12204 24324
rect 12072 24278 12124 24284
rect 12176 24138 12204 24296
rect 12164 24132 12216 24138
rect 12164 24074 12216 24080
rect 11980 24064 12032 24070
rect 11980 24006 12032 24012
rect 11992 23866 12020 24006
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11980 23860 12032 23866
rect 11980 23802 12032 23808
rect 12164 23588 12216 23594
rect 12164 23530 12216 23536
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 11888 22568 11940 22574
rect 11940 22528 12112 22556
rect 11888 22510 11940 22516
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10876 22024 10928 22030
rect 10876 21966 10928 21972
rect 10508 21684 10560 21690
rect 10508 21626 10560 21632
rect 10324 21480 10376 21486
rect 10324 21422 10376 21428
rect 10336 21146 10364 21422
rect 10324 21140 10376 21146
rect 10324 21082 10376 21088
rect 10520 20262 10548 21626
rect 10888 21146 10916 21966
rect 10980 21536 11008 22102
rect 11072 21894 11100 22374
rect 11796 22094 11848 22098
rect 11796 22092 12020 22094
rect 11848 22066 12020 22092
rect 11796 22034 11848 22040
rect 11888 22024 11940 22030
rect 11888 21966 11940 21972
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11060 21548 11112 21554
rect 10980 21508 11060 21536
rect 11060 21490 11112 21496
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10980 21010 11008 21286
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11336 20936 11388 20942
rect 11336 20878 11388 20884
rect 11716 20924 11744 21830
rect 11808 21690 11836 21830
rect 11900 21690 11928 21966
rect 11796 21684 11848 21690
rect 11796 21626 11848 21632
rect 11888 21684 11940 21690
rect 11888 21626 11940 21632
rect 11900 21146 11928 21626
rect 11992 21554 12020 22066
rect 12084 21690 12112 22528
rect 12176 21690 12204 23530
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12164 21684 12216 21690
rect 12164 21626 12216 21632
rect 11980 21548 12032 21554
rect 11980 21490 12032 21496
rect 11980 21344 12032 21350
rect 11980 21286 12032 21292
rect 11992 21146 12020 21286
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11980 21140 12032 21146
rect 11980 21082 12032 21088
rect 11888 20936 11940 20942
rect 11716 20896 11888 20924
rect 10692 20528 10744 20534
rect 10692 20470 10744 20476
rect 10232 20256 10284 20262
rect 10152 20216 10232 20244
rect 9496 20198 9548 20204
rect 10232 20198 10284 20204
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 9508 19854 9536 20198
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 10152 19446 10180 19654
rect 10140 19440 10192 19446
rect 10140 19382 10192 19388
rect 10244 18970 10272 20198
rect 10704 20058 10732 20470
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11072 20058 11100 20402
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11256 19854 11284 20198
rect 11348 20058 11376 20878
rect 11716 20602 11744 20896
rect 11888 20878 11940 20884
rect 11980 20868 12032 20874
rect 11980 20810 12032 20816
rect 11796 20800 11848 20806
rect 11796 20742 11848 20748
rect 11704 20596 11756 20602
rect 11704 20538 11756 20544
rect 11808 20534 11836 20742
rect 11520 20528 11572 20534
rect 11520 20470 11572 20476
rect 11796 20528 11848 20534
rect 11796 20470 11848 20476
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11532 19854 11560 20470
rect 11992 20058 12020 20810
rect 12084 20466 12112 21626
rect 12268 20874 12296 25094
rect 12360 24954 12388 25094
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 12440 24880 12492 24886
rect 12440 24822 12492 24828
rect 12452 24614 12480 24822
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12544 24206 12572 25842
rect 12728 25838 12756 26182
rect 13004 25906 13032 26318
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12992 25900 13044 25906
rect 12992 25842 13044 25848
rect 12716 25832 12768 25838
rect 12716 25774 12768 25780
rect 12820 25430 12848 25842
rect 12900 25764 12952 25770
rect 12900 25706 12952 25712
rect 12808 25424 12860 25430
rect 12808 25366 12860 25372
rect 12808 25152 12860 25158
rect 12912 25140 12940 25706
rect 13004 25294 13032 25842
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 12992 25152 13044 25158
rect 12912 25112 12992 25140
rect 12808 25094 12860 25100
rect 12992 25094 13044 25100
rect 12716 24608 12768 24614
rect 12716 24550 12768 24556
rect 12728 24410 12756 24550
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12820 24274 12848 25094
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12348 24132 12400 24138
rect 12348 24074 12400 24080
rect 12360 23866 12388 24074
rect 12348 23860 12400 23866
rect 12348 23802 12400 23808
rect 12544 23730 12572 24142
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12820 23730 12848 24006
rect 12532 23724 12584 23730
rect 12532 23666 12584 23672
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 22778 12480 23462
rect 12716 22976 12768 22982
rect 12716 22918 12768 22924
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12728 22642 12756 22918
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12532 22092 12584 22098
rect 12532 22034 12584 22040
rect 12544 21486 12572 22034
rect 12728 22030 12756 22578
rect 13004 22506 13032 25094
rect 13096 24682 13124 26318
rect 13280 25786 13308 26454
rect 13372 26042 13400 26930
rect 13544 26784 13596 26790
rect 13544 26726 13596 26732
rect 15936 26784 15988 26790
rect 15936 26726 15988 26732
rect 16120 26784 16172 26790
rect 16120 26726 16172 26732
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 13556 26586 13584 26726
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 15948 26314 15976 26726
rect 15936 26308 15988 26314
rect 15936 26250 15988 26256
rect 13636 26240 13688 26246
rect 13636 26182 13688 26188
rect 13912 26240 13964 26246
rect 13912 26182 13964 26188
rect 13360 26036 13412 26042
rect 13360 25978 13412 25984
rect 13648 25906 13676 26182
rect 13728 26036 13780 26042
rect 13728 25978 13780 25984
rect 13452 25900 13504 25906
rect 13452 25842 13504 25848
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13280 25758 13400 25786
rect 13176 25696 13228 25702
rect 13176 25638 13228 25644
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13188 25498 13216 25638
rect 13176 25492 13228 25498
rect 13176 25434 13228 25440
rect 13280 25294 13308 25638
rect 13372 25498 13400 25758
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13464 25430 13492 25842
rect 13452 25424 13504 25430
rect 13452 25366 13504 25372
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13648 25226 13676 25842
rect 13740 25498 13768 25978
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13832 25702 13860 25842
rect 13820 25696 13872 25702
rect 13820 25638 13872 25644
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13924 25430 13952 26182
rect 15948 25956 15976 26250
rect 16028 25968 16080 25974
rect 14094 25936 14150 25945
rect 15948 25928 16028 25956
rect 16028 25910 16080 25916
rect 16132 25906 16160 26726
rect 16396 26580 16448 26586
rect 16396 26522 16448 26528
rect 16304 26240 16356 26246
rect 16304 26182 16356 26188
rect 14094 25871 14096 25880
rect 14148 25871 14150 25880
rect 15568 25900 15620 25906
rect 14096 25842 14148 25848
rect 15568 25842 15620 25848
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 16120 25900 16172 25906
rect 16120 25842 16172 25848
rect 14108 25498 14136 25842
rect 14462 25800 14518 25809
rect 14462 25735 14464 25744
rect 14516 25735 14518 25744
rect 14464 25706 14516 25712
rect 14096 25492 14148 25498
rect 14096 25434 14148 25440
rect 13912 25424 13964 25430
rect 13912 25366 13964 25372
rect 14096 25288 14148 25294
rect 14096 25230 14148 25236
rect 13636 25220 13688 25226
rect 13636 25162 13688 25168
rect 13728 25152 13780 25158
rect 13728 25094 13780 25100
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13740 24818 13768 25094
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13084 24676 13136 24682
rect 13084 24618 13136 24624
rect 13096 24342 13124 24618
rect 13740 24614 13768 24754
rect 13832 24750 13860 25094
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13084 24336 13136 24342
rect 13136 24284 13216 24290
rect 13084 24278 13216 24284
rect 13096 24262 13216 24278
rect 13188 24206 13216 24262
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12532 21480 12584 21486
rect 12532 21422 12584 21428
rect 12636 21146 12664 21830
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12256 20868 12308 20874
rect 12256 20810 12308 20816
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11520 19848 11572 19854
rect 11520 19790 11572 19796
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11256 19446 11284 19790
rect 11808 19514 11836 19790
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11992 19446 12020 19858
rect 12084 19514 12112 20402
rect 12164 20392 12216 20398
rect 12164 20334 12216 20340
rect 12176 19922 12204 20334
rect 12268 19922 12296 20402
rect 12164 19916 12216 19922
rect 12164 19858 12216 19864
rect 12256 19916 12308 19922
rect 12256 19858 12308 19864
rect 12176 19718 12204 19858
rect 12452 19854 12480 21082
rect 12728 21010 12756 21626
rect 12820 21418 12848 21966
rect 13096 21554 13124 24142
rect 13188 23866 13216 24142
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13464 22438 13492 22578
rect 13268 22432 13320 22438
rect 13268 22374 13320 22380
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13280 22098 13308 22374
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 12808 21412 12860 21418
rect 12808 21354 12860 21360
rect 12900 21344 12952 21350
rect 12900 21286 12952 21292
rect 12912 21010 12940 21286
rect 13096 21146 13124 21490
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12900 21004 12952 21010
rect 12900 20946 12952 20952
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 12532 20800 12584 20806
rect 12532 20742 12584 20748
rect 12544 20466 12572 20742
rect 13280 20534 13308 20878
rect 13268 20528 13320 20534
rect 13268 20470 13320 20476
rect 12532 20460 12584 20466
rect 12532 20402 12584 20408
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 12072 19508 12124 19514
rect 12072 19450 12124 19456
rect 11244 19440 11296 19446
rect 11244 19382 11296 19388
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9588 18624 9640 18630
rect 9588 18566 9640 18572
rect 9600 17542 9628 18566
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9404 17264 9456 17270
rect 9404 17206 9456 17212
rect 8024 17060 8076 17066
rect 8024 17002 8076 17008
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 8036 16454 8064 17002
rect 9600 16658 9628 17478
rect 9784 17134 9812 18838
rect 11256 18834 11284 19382
rect 11520 19372 11572 19378
rect 11572 19320 11652 19334
rect 11520 19314 11652 19320
rect 11532 19306 11652 19314
rect 10692 18828 10744 18834
rect 10692 18770 10744 18776
rect 11244 18828 11296 18834
rect 11244 18770 11296 18776
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 9956 17604 10008 17610
rect 9956 17546 10008 17552
rect 9968 17338 9996 17546
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9772 17128 9824 17134
rect 9824 17088 9904 17116
rect 9772 17070 9824 17076
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 8484 16448 8536 16454
rect 8484 16390 8536 16396
rect 5448 16176 5500 16182
rect 5448 16118 5500 16124
rect 8036 15502 8064 16390
rect 8496 16046 8524 16390
rect 8484 16040 8536 16046
rect 8484 15982 8536 15988
rect 8496 15570 8524 15982
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 5448 15428 5500 15434
rect 5448 15370 5500 15376
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5276 15286 5396 15314
rect 5262 15192 5318 15201
rect 5262 15127 5318 15136
rect 5276 14618 5304 15127
rect 5368 14618 5396 15286
rect 5172 14612 5224 14618
rect 5172 14554 5224 14560
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5356 14612 5408 14618
rect 5356 14554 5408 14560
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 5184 14074 5212 14554
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5184 13802 5212 14010
rect 5276 13802 5304 14350
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13938 5396 14214
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 5264 13796 5316 13802
rect 5264 13738 5316 13744
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3896 12406 4016 12434
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3896 10606 3924 12406
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4632 11898 4660 12174
rect 5000 11898 5028 12854
rect 5184 12238 5212 13738
rect 5276 12986 5304 13738
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5460 12918 5488 15370
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5552 14006 5580 14350
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5552 12986 5580 13942
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5448 12912 5500 12918
rect 5448 12854 5500 12860
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5368 12170 5396 12378
rect 5356 12164 5408 12170
rect 5356 12106 5408 12112
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 5000 11286 5028 11834
rect 5368 11830 5396 12106
rect 5356 11824 5408 11830
rect 5356 11766 5408 11772
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5368 11218 5396 11766
rect 5460 11354 5488 12854
rect 5552 12170 5580 12922
rect 5644 12646 5672 15370
rect 5920 14822 5948 15438
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 7760 15026 7788 15302
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 14482 5948 14758
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 8588 14414 8616 15302
rect 8772 14414 8800 15302
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 6552 14272 6604 14278
rect 6552 14214 6604 14220
rect 6564 13938 6592 14214
rect 8772 14074 8800 14350
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9772 14340 9824 14346
rect 9772 14282 9824 14288
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6920 13796 6972 13802
rect 6920 13738 6972 13744
rect 6932 13530 6960 13738
rect 6920 13524 6972 13530
rect 6920 13466 6972 13472
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5828 12306 5856 12582
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 7024 12238 7052 13262
rect 8772 12714 8800 14010
rect 9140 13734 9168 14282
rect 9784 14074 9812 14282
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9128 13728 9180 13734
rect 9128 13670 9180 13676
rect 9140 13326 9168 13670
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8760 12708 8812 12714
rect 8760 12650 8812 12656
rect 8300 12640 8352 12646
rect 8300 12582 8352 12588
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 8312 12170 8340 12582
rect 5540 12164 5592 12170
rect 5540 12106 5592 12112
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5356 11212 5408 11218
rect 5356 11154 5408 11160
rect 4160 11008 4212 11014
rect 4160 10950 4212 10956
rect 4172 10742 4200 10950
rect 5552 10810 5580 12106
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 7576 11898 7604 12038
rect 8220 11898 8248 12038
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8680 11880 8708 12582
rect 8772 12102 8800 12650
rect 9140 12646 9168 13262
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8852 11892 8904 11898
rect 8680 11852 8852 11880
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6012 10810 6040 11698
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6196 11354 6224 11494
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 6472 10810 6500 11698
rect 8116 11688 8168 11694
rect 8114 11656 8116 11665
rect 8168 11656 8170 11665
rect 8114 11591 8170 11600
rect 8680 11082 8708 11852
rect 8852 11834 8904 11840
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 8680 10742 8708 11018
rect 9048 10742 9076 12038
rect 9876 11626 9904 17088
rect 9956 15904 10008 15910
rect 9956 15846 10008 15852
rect 9968 15570 9996 15846
rect 9956 15564 10008 15570
rect 9956 15506 10008 15512
rect 10428 14958 10456 18702
rect 10704 18290 10732 18770
rect 11624 18766 11652 19306
rect 11612 18760 11664 18766
rect 11612 18702 11664 18708
rect 12268 18714 12296 19722
rect 12544 19446 12572 20402
rect 12716 20256 12768 20262
rect 12716 20198 12768 20204
rect 12728 20058 12756 20198
rect 13188 20058 13216 20402
rect 13358 20088 13414 20097
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 13176 20052 13228 20058
rect 13358 20023 13360 20032
rect 13176 19994 13228 20000
rect 13412 20023 13414 20032
rect 13360 19994 13412 20000
rect 13464 19786 13492 22374
rect 13832 21962 13860 24686
rect 14004 24268 14056 24274
rect 14004 24210 14056 24216
rect 14016 23662 14044 24210
rect 14004 23656 14056 23662
rect 14004 23598 14056 23604
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13924 22642 13952 23258
rect 14108 22778 14136 25230
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14292 23730 14320 24006
rect 14280 23724 14332 23730
rect 14280 23666 14332 23672
rect 14384 23322 14412 24006
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14372 22976 14424 22982
rect 14372 22918 14424 22924
rect 14096 22772 14148 22778
rect 14096 22714 14148 22720
rect 14280 22772 14332 22778
rect 14280 22714 14332 22720
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13648 21010 13676 21558
rect 13832 21010 13860 21626
rect 13924 21146 13952 22578
rect 14188 22568 14240 22574
rect 14188 22510 14240 22516
rect 14004 22228 14056 22234
rect 14004 22170 14056 22176
rect 14016 21622 14044 22170
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14004 21616 14056 21622
rect 14004 21558 14056 21564
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13648 20330 13676 20946
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13832 19854 13860 20742
rect 13924 20602 13952 21082
rect 13912 20596 13964 20602
rect 13912 20538 13964 20544
rect 13924 20466 13952 20538
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 14108 19922 14136 21830
rect 14200 20602 14228 22510
rect 14292 22438 14320 22714
rect 14384 22574 14412 22918
rect 14476 22778 14504 25706
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14936 25498 14964 25638
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 15580 25362 15608 25842
rect 15660 25696 15712 25702
rect 15660 25638 15712 25644
rect 15568 25356 15620 25362
rect 15568 25298 15620 25304
rect 15292 25288 15344 25294
rect 15292 25230 15344 25236
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15212 24410 15240 24686
rect 15304 24410 15332 25230
rect 15384 24676 15436 24682
rect 15384 24618 15436 24624
rect 15200 24404 15252 24410
rect 15200 24346 15252 24352
rect 15292 24404 15344 24410
rect 15292 24346 15344 24352
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14568 23798 14596 24142
rect 14556 23792 14608 23798
rect 14556 23734 14608 23740
rect 15304 23730 15332 24210
rect 15396 23730 15424 24618
rect 15476 24200 15528 24206
rect 15476 24142 15528 24148
rect 15488 23866 15516 24142
rect 15476 23860 15528 23866
rect 15476 23802 15528 23808
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15384 23724 15436 23730
rect 15384 23666 15436 23672
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23050 15240 23462
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 14464 22772 14516 22778
rect 14464 22714 14516 22720
rect 14372 22568 14424 22574
rect 14372 22510 14424 22516
rect 14280 22432 14332 22438
rect 14280 22374 14332 22380
rect 14292 22030 14320 22374
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14372 21956 14424 21962
rect 14372 21898 14424 21904
rect 14384 21332 14412 21898
rect 14476 21690 14504 22714
rect 15304 22234 15332 23258
rect 15396 23186 15424 23666
rect 15384 23180 15436 23186
rect 15384 23122 15436 23128
rect 15580 23118 15608 25298
rect 15672 24954 15700 25638
rect 15764 25294 15792 25842
rect 16212 25832 16264 25838
rect 15856 25780 16212 25786
rect 15856 25774 16264 25780
rect 15856 25758 16252 25774
rect 15856 25498 15884 25758
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 16028 25696 16080 25702
rect 16080 25644 16252 25650
rect 16028 25638 16252 25644
rect 15844 25492 15896 25498
rect 15844 25434 15896 25440
rect 15948 25378 15976 25638
rect 16040 25622 16252 25638
rect 16120 25424 16172 25430
rect 15948 25372 16120 25378
rect 15948 25366 16172 25372
rect 15948 25350 16160 25366
rect 16224 25362 16252 25622
rect 16316 25362 16344 26182
rect 16408 25906 16436 26522
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 16488 26376 16540 26382
rect 16488 26318 16540 26324
rect 16500 26042 16528 26318
rect 16580 26308 16632 26314
rect 16580 26250 16632 26256
rect 16592 26042 16620 26250
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16580 26036 16632 26042
rect 16580 25978 16632 25984
rect 17052 25906 17080 26454
rect 17236 26382 17264 26726
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17408 26376 17460 26382
rect 17512 26364 17540 26930
rect 18800 26790 18828 26930
rect 18880 26920 18932 26926
rect 18880 26862 18932 26868
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18788 26784 18840 26790
rect 18788 26726 18840 26732
rect 18144 26444 18196 26450
rect 18144 26386 18196 26392
rect 17460 26336 17540 26364
rect 17408 26318 17460 26324
rect 17132 26240 17184 26246
rect 17132 26182 17184 26188
rect 17144 25906 17172 26182
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 16212 25356 16264 25362
rect 15752 25288 15804 25294
rect 15752 25230 15804 25236
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15660 24812 15712 24818
rect 15764 24800 15792 25230
rect 15948 24818 15976 25350
rect 16212 25298 16264 25304
rect 16304 25356 16356 25362
rect 16304 25298 16356 25304
rect 16212 25152 16264 25158
rect 16212 25094 16264 25100
rect 16224 24954 16252 25094
rect 16212 24948 16264 24954
rect 16212 24890 16264 24896
rect 15712 24772 15792 24800
rect 15936 24812 15988 24818
rect 15660 24754 15712 24760
rect 15936 24754 15988 24760
rect 15844 24744 15896 24750
rect 15844 24686 15896 24692
rect 15752 24676 15804 24682
rect 15752 24618 15804 24624
rect 15764 24342 15792 24618
rect 15856 24410 15884 24686
rect 15844 24404 15896 24410
rect 15844 24346 15896 24352
rect 15752 24336 15804 24342
rect 15752 24278 15804 24284
rect 15752 24200 15804 24206
rect 15752 24142 15804 24148
rect 15764 23866 15792 24142
rect 15856 23866 15884 24346
rect 16316 24342 16344 25298
rect 16408 24682 16436 25842
rect 16672 25764 16724 25770
rect 16672 25706 16724 25712
rect 16488 25696 16540 25702
rect 16488 25638 16540 25644
rect 16580 25696 16632 25702
rect 16580 25638 16632 25644
rect 16500 24682 16528 25638
rect 16592 25498 16620 25638
rect 16580 25492 16632 25498
rect 16580 25434 16632 25440
rect 16684 25362 16712 25706
rect 17052 25498 17080 25842
rect 17144 25809 17172 25842
rect 17130 25800 17186 25809
rect 17130 25735 17186 25744
rect 17040 25492 17092 25498
rect 17040 25434 17092 25440
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16396 24676 16448 24682
rect 16396 24618 16448 24624
rect 16488 24676 16540 24682
rect 16488 24618 16540 24624
rect 16304 24336 16356 24342
rect 16304 24278 16356 24284
rect 15752 23860 15804 23866
rect 15752 23802 15804 23808
rect 15844 23860 15896 23866
rect 15844 23802 15896 23808
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 15764 23322 15792 23666
rect 16316 23662 16344 24278
rect 16408 24274 16436 24618
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16500 23730 16528 24618
rect 17144 24410 17172 25735
rect 17132 24404 17184 24410
rect 17132 24346 17184 24352
rect 16488 23724 16540 23730
rect 16488 23666 16540 23672
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 17132 23520 17184 23526
rect 17132 23462 17184 23468
rect 15752 23316 15804 23322
rect 15752 23258 15804 23264
rect 17144 23186 17172 23462
rect 17132 23180 17184 23186
rect 17132 23122 17184 23128
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 15580 22778 15608 23054
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 14648 22160 14700 22166
rect 14648 22102 14700 22108
rect 14660 21690 14688 22102
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15660 22024 15712 22030
rect 15660 21966 15712 21972
rect 14464 21684 14516 21690
rect 14464 21626 14516 21632
rect 14648 21684 14700 21690
rect 14648 21626 14700 21632
rect 14660 21486 14688 21626
rect 15028 21554 15056 21966
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15304 21554 15332 21830
rect 15672 21554 15700 21966
rect 15016 21548 15068 21554
rect 15016 21490 15068 21496
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 16672 21548 16724 21554
rect 16672 21490 16724 21496
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14292 21304 14412 21332
rect 14188 20596 14240 20602
rect 14188 20538 14240 20544
rect 14200 20466 14228 20538
rect 14292 20466 14320 21304
rect 16684 20942 16712 21490
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16672 20936 16724 20942
rect 16672 20878 16724 20884
rect 14372 20868 14424 20874
rect 14372 20810 14424 20816
rect 14384 20534 14412 20810
rect 14372 20528 14424 20534
rect 14372 20470 14424 20476
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14188 20256 14240 20262
rect 14188 20198 14240 20204
rect 14200 20058 14228 20198
rect 14188 20052 14240 20058
rect 14188 19994 14240 20000
rect 14096 19916 14148 19922
rect 14096 19858 14148 19864
rect 13820 19848 13872 19854
rect 13820 19790 13872 19796
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13464 19514 13492 19722
rect 14476 19718 14504 20402
rect 14924 20256 14976 20262
rect 14924 20198 14976 20204
rect 14936 19786 14964 20198
rect 15120 19922 15148 20470
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15384 20392 15436 20398
rect 15384 20334 15436 20340
rect 15396 20058 15424 20334
rect 15488 20058 15516 20402
rect 16684 20398 16712 20878
rect 16960 20806 16988 21422
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16856 20528 16908 20534
rect 16856 20470 16908 20476
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16868 20058 16896 20470
rect 16960 20466 16988 20742
rect 17144 20602 17172 20878
rect 17132 20596 17184 20602
rect 17132 20538 17184 20544
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 16960 20058 16988 20402
rect 17420 20330 17448 26318
rect 18156 25974 18184 26386
rect 18524 26382 18552 26726
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18788 26376 18840 26382
rect 18892 26364 18920 26862
rect 19076 26382 19104 26930
rect 19352 26858 19380 27406
rect 19340 26852 19392 26858
rect 19340 26794 19392 26800
rect 19248 26784 19300 26790
rect 19248 26726 19300 26732
rect 18840 26336 18920 26364
rect 19064 26376 19116 26382
rect 18788 26318 18840 26324
rect 19064 26318 19116 26324
rect 19156 26376 19208 26382
rect 19156 26318 19208 26324
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18248 26042 18276 26182
rect 18236 26036 18288 26042
rect 18236 25978 18288 25984
rect 17592 25968 17644 25974
rect 17592 25910 17644 25916
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 17604 23730 17632 25910
rect 18800 25838 18828 26318
rect 19076 25974 19104 26318
rect 19064 25968 19116 25974
rect 19064 25910 19116 25916
rect 18328 25832 18380 25838
rect 18328 25774 18380 25780
rect 18788 25832 18840 25838
rect 18788 25774 18840 25780
rect 18340 24818 18368 25774
rect 18328 24812 18380 24818
rect 18328 24754 18380 24760
rect 17960 24676 18012 24682
rect 17960 24618 18012 24624
rect 17972 23798 18000 24618
rect 18236 24268 18288 24274
rect 18236 24210 18288 24216
rect 18248 23866 18276 24210
rect 18236 23860 18288 23866
rect 18236 23802 18288 23808
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 17592 23724 17644 23730
rect 17592 23666 17644 23672
rect 17604 22778 17632 23666
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 18052 22568 18104 22574
rect 18052 22510 18104 22516
rect 18064 22166 18092 22510
rect 18052 22160 18104 22166
rect 18052 22102 18104 22108
rect 17592 22092 17644 22098
rect 17592 22034 17644 22040
rect 17604 21690 17632 22034
rect 17684 22024 17736 22030
rect 17684 21966 17736 21972
rect 17592 21684 17644 21690
rect 17592 21626 17644 21632
rect 17592 20936 17644 20942
rect 17696 20924 17724 21966
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17644 20896 17724 20924
rect 17592 20878 17644 20884
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 15108 19916 15160 19922
rect 15108 19858 15160 19864
rect 16856 19916 16908 19922
rect 16960 19904 16988 19994
rect 16908 19876 16988 19904
rect 16856 19858 16908 19864
rect 14924 19780 14976 19786
rect 14924 19722 14976 19728
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 12808 19508 12860 19514
rect 12808 19450 12860 19456
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 12532 19440 12584 19446
rect 12532 19382 12584 19388
rect 10876 18692 10928 18698
rect 10876 18634 10928 18640
rect 11796 18692 11848 18698
rect 12268 18686 12388 18714
rect 11796 18634 11848 18640
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10704 16726 10732 18226
rect 10888 18154 10916 18634
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10876 18148 10928 18154
rect 10876 18090 10928 18096
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10520 16046 10548 16390
rect 10508 16040 10560 16046
rect 10508 15982 10560 15988
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10520 14890 10548 15982
rect 10600 15428 10652 15434
rect 10600 15370 10652 15376
rect 10612 15162 10640 15370
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10508 14884 10560 14890
rect 10508 14826 10560 14832
rect 10520 14074 10548 14826
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 12986 10456 13262
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10980 12714 11008 17206
rect 11072 16250 11100 18566
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11348 17746 11376 18226
rect 11808 18222 11836 18634
rect 12360 18340 12388 18686
rect 12820 18408 12848 19450
rect 13464 18970 13492 19450
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 14556 18964 14608 18970
rect 14556 18906 14608 18912
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13268 18624 13320 18630
rect 13268 18566 13320 18572
rect 12820 18380 12940 18408
rect 12532 18352 12584 18358
rect 12360 18312 12532 18340
rect 12532 18294 12584 18300
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11336 17740 11388 17746
rect 11336 17682 11388 17688
rect 11808 17678 11836 18158
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 12348 17536 12400 17542
rect 12348 17478 12400 17484
rect 11256 17270 11284 17478
rect 12360 17338 12388 17478
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11256 16794 11284 17206
rect 11980 17128 12032 17134
rect 11980 17070 12032 17076
rect 11992 16794 12020 17070
rect 11244 16788 11296 16794
rect 11244 16730 11296 16736
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11348 15162 11376 15302
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11164 13938 11192 14214
rect 11532 14074 11560 16594
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11808 16046 11836 16390
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11992 15910 12020 16730
rect 12452 16454 12480 18022
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16114 12480 16390
rect 12636 16114 12664 17070
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12072 16040 12124 16046
rect 12072 15982 12124 15988
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15502 12020 15846
rect 12084 15706 12112 15982
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12636 15502 12664 16050
rect 12820 15570 12848 18226
rect 12808 15564 12860 15570
rect 12808 15506 12860 15512
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 12624 15496 12676 15502
rect 12624 15438 12676 15444
rect 11992 15094 12020 15438
rect 11980 15088 12032 15094
rect 11980 15030 12032 15036
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11624 14618 11652 14962
rect 11992 14618 12020 15030
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 10612 10996 10640 11698
rect 11164 11218 11192 13874
rect 11532 12306 11560 14010
rect 11992 13394 12020 14554
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12452 13530 12480 13874
rect 12820 13870 12848 15506
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11520 12300 11572 12306
rect 11520 12242 11572 12248
rect 11992 11898 12020 13330
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12624 12844 12676 12850
rect 12624 12786 12676 12792
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12452 12238 12480 12582
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 12636 11150 12664 12786
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 10692 11008 10744 11014
rect 10612 10968 10692 10996
rect 10692 10950 10744 10956
rect 4160 10736 4212 10742
rect 4160 10678 4212 10684
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 3148 10600 3200 10606
rect 3148 10542 3200 10548
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 3160 6914 3188 10542
rect 3896 10266 3924 10542
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 1596 6886 1716 6914
rect 2976 6886 3188 6914
rect 1596 6662 1624 6886
rect 1584 6656 1636 6662
rect 1584 6598 1636 6604
rect 2976 4826 3004 6886
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 9048 2514 9076 10678
rect 10704 10538 10732 10950
rect 12728 10538 12756 13126
rect 12820 12850 12848 13806
rect 12912 13802 12940 18380
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13084 18284 13136 18290
rect 13084 18226 13136 18232
rect 13004 17542 13032 18226
rect 13096 18086 13124 18226
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12992 17536 13044 17542
rect 12992 17478 13044 17484
rect 13004 17066 13032 17478
rect 13096 17202 13124 18022
rect 13188 17542 13216 18566
rect 13280 18290 13308 18566
rect 14016 18358 14044 18634
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 13280 17678 13308 18226
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12992 17060 13044 17066
rect 12992 17002 13044 17008
rect 13004 16522 13032 17002
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 13004 15706 13032 16458
rect 13176 16448 13228 16454
rect 13176 16390 13228 16396
rect 13188 16046 13216 16390
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13176 16040 13228 16046
rect 13176 15982 13228 15988
rect 12992 15700 13044 15706
rect 12992 15642 13044 15648
rect 13280 15484 13308 16050
rect 13360 15700 13412 15706
rect 13464 15688 13492 18226
rect 13728 18148 13780 18154
rect 13728 18090 13780 18096
rect 13740 17814 13768 18090
rect 13832 17882 13860 18226
rect 14292 17882 14320 18226
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 14280 17876 14332 17882
rect 14280 17818 14332 17824
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 14004 17672 14056 17678
rect 14004 17614 14056 17620
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14280 17672 14332 17678
rect 14280 17614 14332 17620
rect 14016 17202 14044 17614
rect 14108 17542 14136 17614
rect 14096 17536 14148 17542
rect 14096 17478 14148 17484
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13556 15706 13584 16594
rect 13648 16590 13676 17138
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13648 16250 13676 16526
rect 14016 16522 14044 17138
rect 14004 16516 14056 16522
rect 14004 16458 14056 16464
rect 14108 16454 14136 17478
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 14004 16108 14056 16114
rect 14108 16096 14136 16390
rect 14292 16114 14320 17614
rect 14384 17610 14412 18158
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14384 16590 14412 16934
rect 14476 16794 14504 17138
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 14372 16448 14424 16454
rect 14424 16408 14504 16436
rect 14372 16390 14424 16396
rect 14056 16068 14136 16096
rect 14004 16050 14056 16056
rect 13412 15660 13492 15688
rect 13544 15700 13596 15706
rect 13360 15642 13412 15648
rect 13544 15642 13596 15648
rect 14108 15586 14136 16068
rect 14280 16108 14332 16114
rect 14280 16050 14332 16056
rect 14108 15558 14228 15586
rect 14476 15570 14504 16408
rect 13452 15496 13504 15502
rect 13280 15456 13452 15484
rect 13452 15438 13504 15444
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13464 15026 13492 15438
rect 14108 15162 14136 15438
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13464 14550 13492 14962
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13648 14618 13676 14894
rect 13820 14816 13872 14822
rect 13820 14758 13872 14764
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13452 14544 13504 14550
rect 13452 14486 13504 14492
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12912 13274 12940 13738
rect 13556 13530 13584 14010
rect 13832 13530 13860 14758
rect 14200 13734 14228 15558
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 14280 15496 14332 15502
rect 14280 15438 14332 15444
rect 14292 15162 14320 15438
rect 14280 15156 14332 15162
rect 14280 15098 14332 15104
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14618 14412 14962
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14568 14074 14596 18906
rect 14660 17882 14688 19246
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17066 14780 17478
rect 14936 17202 14964 19722
rect 15120 18766 15148 19858
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 15396 19718 15424 19790
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15396 19310 15424 19654
rect 15672 19514 15700 19790
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15384 19304 15436 19310
rect 15384 19246 15436 19252
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 16132 18698 16160 19790
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 16224 19514 16252 19654
rect 16212 19508 16264 19514
rect 16212 19450 16264 19456
rect 16396 19440 16448 19446
rect 16396 19382 16448 19388
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16224 18290 16252 18566
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15936 18284 15988 18290
rect 15936 18226 15988 18232
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 15212 17882 15240 18226
rect 15304 17882 15332 18226
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15200 17876 15252 17882
rect 15200 17818 15252 17824
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15396 17542 15424 18022
rect 15476 17672 15528 17678
rect 15476 17614 15528 17620
rect 15488 17542 15516 17614
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15384 17536 15436 17542
rect 15384 17478 15436 17484
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15028 17202 15056 17478
rect 15764 17338 15792 18226
rect 15856 17882 15884 18226
rect 15948 18086 15976 18226
rect 15936 18080 15988 18086
rect 15988 18040 16068 18068
rect 15936 18022 15988 18028
rect 15844 17876 15896 17882
rect 15844 17818 15896 17824
rect 15936 17808 15988 17814
rect 15936 17750 15988 17756
rect 15948 17678 15976 17750
rect 15936 17672 15988 17678
rect 15936 17614 15988 17620
rect 15948 17524 15976 17614
rect 15856 17496 15976 17524
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15856 17270 15884 17496
rect 16040 17338 16068 18040
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 16028 17332 16080 17338
rect 16028 17274 16080 17280
rect 15844 17264 15896 17270
rect 15844 17206 15896 17212
rect 16132 17202 16160 17546
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 16120 17196 16172 17202
rect 16120 17138 16172 17144
rect 14740 17060 14792 17066
rect 14740 17002 14792 17008
rect 14752 16794 14780 17002
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14936 16522 14964 17138
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14660 15502 14688 16186
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14752 15450 14780 16458
rect 15120 15638 15148 16934
rect 15764 16250 15792 17070
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15212 15706 15240 16050
rect 16408 16046 16436 19382
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17316 18760 17368 18766
rect 17316 18702 17368 18708
rect 17236 18630 17264 18702
rect 17224 18624 17276 18630
rect 17224 18566 17276 18572
rect 17040 18284 17092 18290
rect 17040 18226 17092 18232
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16488 18080 16540 18086
rect 16488 18022 16540 18028
rect 16500 17882 16528 18022
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16684 17746 16712 18158
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16592 16658 16620 17614
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16672 17332 16724 17338
rect 16672 17274 16724 17280
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16684 16590 16712 17274
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16776 16794 16804 17138
rect 16868 17134 16896 17478
rect 16960 17338 16988 17614
rect 17052 17542 17080 18226
rect 17236 18154 17264 18566
rect 17328 18358 17356 18702
rect 17604 18426 17632 20878
rect 17880 20806 17908 21014
rect 18340 20806 18368 24754
rect 19076 24750 19104 25910
rect 19168 25906 19196 26318
rect 19156 25900 19208 25906
rect 19156 25842 19208 25848
rect 19260 25838 19288 26726
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19352 25974 19380 26386
rect 19444 26382 19472 27406
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27130 20024 27406
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 20088 26994 20116 27406
rect 20260 27328 20312 27334
rect 20260 27270 20312 27276
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 20272 27062 20300 27270
rect 20456 27130 20484 27270
rect 20444 27124 20496 27130
rect 20444 27066 20496 27072
rect 20260 27056 20312 27062
rect 20260 26998 20312 27004
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20076 26988 20128 26994
rect 20076 26930 20128 26936
rect 21008 26586 21036 26998
rect 21376 26994 21404 27610
rect 23400 27606 23428 29158
rect 23572 29106 23624 29112
rect 23480 28960 23532 28966
rect 23480 28902 23532 28908
rect 23492 28558 23520 28902
rect 23480 28552 23532 28558
rect 23480 28494 23532 28500
rect 23676 28490 23704 29242
rect 24320 29238 24348 29446
rect 23940 29232 23992 29238
rect 23940 29174 23992 29180
rect 24308 29232 24360 29238
rect 24308 29174 24360 29180
rect 23952 28762 23980 29174
rect 24412 29170 24440 29446
rect 24400 29164 24452 29170
rect 24400 29106 24452 29112
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 24412 28642 24440 29106
rect 24412 28626 24532 28642
rect 24412 28620 24544 28626
rect 24412 28614 24492 28620
rect 24492 28562 24544 28568
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 23584 28014 23612 28358
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23388 27600 23440 27606
rect 23388 27542 23440 27548
rect 22468 27532 22520 27538
rect 22468 27474 22520 27480
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22100 27056 22152 27062
rect 22100 26998 22152 27004
rect 21272 26988 21324 26994
rect 21272 26930 21324 26936
rect 21364 26988 21416 26994
rect 21364 26930 21416 26936
rect 20996 26580 21048 26586
rect 20996 26522 21048 26528
rect 21086 26480 21142 26489
rect 21086 26415 21088 26424
rect 21140 26415 21142 26424
rect 21088 26386 21140 26392
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19444 26042 19472 26318
rect 20720 26240 20772 26246
rect 20720 26182 20772 26188
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 26036 19484 26042
rect 19432 25978 19484 25984
rect 19340 25968 19392 25974
rect 19340 25910 19392 25916
rect 19248 25832 19300 25838
rect 19300 25792 19380 25820
rect 19248 25774 19300 25780
rect 19352 24818 19380 25792
rect 20732 25430 20760 26182
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20916 25294 20944 25638
rect 20904 25288 20956 25294
rect 20904 25230 20956 25236
rect 20076 25152 20128 25158
rect 20076 25094 20128 25100
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19340 24812 19392 24818
rect 19340 24754 19392 24760
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 18420 23112 18472 23118
rect 18420 23054 18472 23060
rect 18432 22574 18460 23054
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18616 22778 18644 22918
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18420 22568 18472 22574
rect 18420 22510 18472 22516
rect 19260 21690 19288 23462
rect 19996 23322 20024 24754
rect 20088 24070 20116 25094
rect 20456 24818 20484 25094
rect 20824 24954 20852 25094
rect 20812 24948 20864 24954
rect 20812 24890 20864 24896
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20076 24064 20128 24070
rect 20076 24006 20128 24012
rect 20272 23730 20300 24278
rect 20444 24064 20496 24070
rect 20496 24024 20576 24052
rect 20444 24006 20496 24012
rect 20548 23866 20576 24024
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20548 23730 20576 23802
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20272 23322 20300 23666
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19984 23316 20036 23322
rect 19984 23258 20036 23264
rect 20260 23316 20312 23322
rect 20260 23258 20312 23264
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 19352 22098 19380 22918
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19248 21684 19300 21690
rect 19076 21644 19248 21672
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 18328 20800 18380 20806
rect 18328 20742 18380 20748
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17696 20058 17724 20538
rect 17776 20256 17828 20262
rect 17776 20198 17828 20204
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17696 19854 17724 19994
rect 17788 19854 17816 20198
rect 17880 20058 17908 20742
rect 17958 20088 18014 20097
rect 17868 20052 17920 20058
rect 17958 20023 17960 20032
rect 17868 19994 17920 20000
rect 18012 20023 18014 20032
rect 17960 19994 18012 20000
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 17684 19848 17736 19854
rect 17684 19790 17736 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17960 19780 18012 19786
rect 17960 19722 18012 19728
rect 17972 19514 18000 19722
rect 18800 19514 18828 19926
rect 19076 19922 19104 21644
rect 19248 21626 19300 21632
rect 19444 21486 19472 23258
rect 20916 23202 20944 25230
rect 21008 24886 21036 25842
rect 21100 24886 21128 26386
rect 21284 26042 21312 26930
rect 22112 26330 22140 26998
rect 22204 26858 22232 27270
rect 22480 26994 22508 27474
rect 23204 27328 23256 27334
rect 23204 27270 23256 27276
rect 23216 26994 23244 27270
rect 22468 26988 22520 26994
rect 22468 26930 22520 26936
rect 23204 26988 23256 26994
rect 23204 26930 23256 26936
rect 22192 26852 22244 26858
rect 22192 26794 22244 26800
rect 22204 26586 22232 26794
rect 22480 26586 22508 26930
rect 22928 26784 22980 26790
rect 22928 26726 22980 26732
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 22192 26580 22244 26586
rect 22192 26522 22244 26528
rect 22468 26580 22520 26586
rect 22468 26522 22520 26528
rect 22940 26489 22968 26726
rect 22926 26480 22982 26489
rect 22926 26415 22928 26424
rect 22980 26415 22982 26424
rect 22928 26386 22980 26392
rect 23584 26382 23612 26726
rect 23296 26376 23348 26382
rect 21456 26308 21508 26314
rect 22112 26302 22232 26330
rect 23572 26376 23624 26382
rect 23296 26318 23348 26324
rect 23400 26324 23572 26330
rect 23400 26318 23624 26324
rect 21456 26250 21508 26256
rect 21364 26240 21416 26246
rect 21364 26182 21416 26188
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21376 25922 21404 26182
rect 21284 25894 21404 25922
rect 21284 25702 21312 25894
rect 21272 25696 21324 25702
rect 21272 25638 21324 25644
rect 21284 25158 21312 25638
rect 21272 25152 21324 25158
rect 21272 25094 21324 25100
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 21088 24880 21140 24886
rect 21088 24822 21140 24828
rect 21008 24206 21036 24822
rect 21100 24342 21128 24822
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 21100 23798 21128 24278
rect 21088 23792 21140 23798
rect 21140 23752 21220 23780
rect 21088 23734 21140 23740
rect 20916 23174 21128 23202
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20916 22778 20944 23174
rect 21100 23118 21128 23174
rect 20996 23112 21048 23118
rect 20994 23080 20996 23089
rect 21088 23112 21140 23118
rect 21048 23080 21050 23089
rect 21088 23054 21140 23060
rect 20994 23015 21050 23024
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 19524 22500 19576 22506
rect 19524 22442 19576 22448
rect 19536 22030 19564 22442
rect 20916 22234 20944 22714
rect 21008 22642 21036 23015
rect 21192 22778 21220 23752
rect 21284 23526 21312 25094
rect 21364 24676 21416 24682
rect 21468 24664 21496 26250
rect 22204 26246 22232 26302
rect 22192 26240 22244 26246
rect 22192 26182 22244 26188
rect 23308 25770 23336 26318
rect 23400 26302 23612 26318
rect 23296 25764 23348 25770
rect 23296 25706 23348 25712
rect 23400 25702 23428 26302
rect 22376 25696 22428 25702
rect 22376 25638 22428 25644
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22928 25696 22980 25702
rect 22928 25638 22980 25644
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21416 24636 21496 24664
rect 21364 24618 21416 24624
rect 21376 24138 21404 24618
rect 21744 24206 21772 25094
rect 21836 24954 21864 25298
rect 22388 24954 22416 25638
rect 22664 25430 22692 25638
rect 22652 25424 22704 25430
rect 22652 25366 22704 25372
rect 21824 24948 21876 24954
rect 21824 24890 21876 24896
rect 22376 24948 22428 24954
rect 22376 24890 22428 24896
rect 22100 24676 22152 24682
rect 22100 24618 22152 24624
rect 21732 24200 21784 24206
rect 21732 24142 21784 24148
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21744 23866 21772 24142
rect 22112 24052 22140 24618
rect 22388 24410 22416 24890
rect 22664 24886 22692 25366
rect 22940 25294 22968 25638
rect 23400 25514 23428 25638
rect 23308 25486 23428 25514
rect 23676 25498 23704 28426
rect 24400 27668 24452 27674
rect 24400 27610 24452 27616
rect 24412 27130 24440 27610
rect 24504 27470 24532 28562
rect 24492 27464 24544 27470
rect 24492 27406 24544 27412
rect 24504 27130 24532 27406
rect 24400 27124 24452 27130
rect 24400 27066 24452 27072
rect 24492 27124 24544 27130
rect 24492 27066 24544 27072
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24320 26518 24348 26930
rect 24688 26586 24716 29514
rect 24872 29306 24900 29582
rect 25148 29306 25176 29650
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 28356 29640 28408 29646
rect 28356 29582 28408 29588
rect 29184 29640 29236 29646
rect 29184 29582 29236 29588
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 25136 29300 25188 29306
rect 25136 29242 25188 29248
rect 24872 29170 24900 29242
rect 24860 29164 24912 29170
rect 24860 29106 24912 29112
rect 25044 29164 25096 29170
rect 25044 29106 25096 29112
rect 25136 29164 25188 29170
rect 25136 29106 25188 29112
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24780 27674 24808 28630
rect 24872 28422 24900 29106
rect 25056 28490 25084 29106
rect 25148 28626 25176 29106
rect 26988 29034 27016 29582
rect 27068 29572 27120 29578
rect 27068 29514 27120 29520
rect 26976 29028 27028 29034
rect 26976 28970 27028 28976
rect 26240 28960 26292 28966
rect 26240 28902 26292 28908
rect 25136 28620 25188 28626
rect 25136 28562 25188 28568
rect 26252 28558 26280 28902
rect 26516 28688 26568 28694
rect 26516 28630 26568 28636
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 26332 28552 26384 28558
rect 26332 28494 26384 28500
rect 25044 28484 25096 28490
rect 25044 28426 25096 28432
rect 25412 28484 25464 28490
rect 25412 28426 25464 28432
rect 24860 28416 24912 28422
rect 24860 28358 24912 28364
rect 24768 27668 24820 27674
rect 24768 27610 24820 27616
rect 24768 26988 24820 26994
rect 24768 26930 24820 26936
rect 24676 26580 24728 26586
rect 24676 26522 24728 26528
rect 24308 26512 24360 26518
rect 24308 26454 24360 26460
rect 23756 26444 23808 26450
rect 23756 26386 23808 26392
rect 23768 25498 23796 26386
rect 23664 25492 23716 25498
rect 23308 25430 23336 25486
rect 23664 25434 23716 25440
rect 23756 25492 23808 25498
rect 23756 25434 23808 25440
rect 23296 25424 23348 25430
rect 23296 25366 23348 25372
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 22468 24880 22520 24886
rect 22468 24822 22520 24828
rect 22652 24880 22704 24886
rect 22652 24822 22704 24828
rect 22480 24614 22508 24822
rect 22468 24608 22520 24614
rect 22468 24550 22520 24556
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22376 24404 22428 24410
rect 22376 24346 22428 24352
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 22204 24206 22232 24346
rect 22192 24200 22244 24206
rect 22192 24142 22244 24148
rect 22192 24064 22244 24070
rect 22112 24024 22192 24052
rect 22192 24006 22244 24012
rect 21732 23860 21784 23866
rect 21732 23802 21784 23808
rect 22204 23730 22232 24006
rect 22848 23730 22876 24346
rect 22940 24070 22968 25230
rect 23216 24954 23244 25230
rect 23308 25226 23336 25366
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23296 25220 23348 25226
rect 23296 25162 23348 25168
rect 23204 24948 23256 24954
rect 23204 24890 23256 24896
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 22928 24064 22980 24070
rect 22928 24006 22980 24012
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22468 23724 22520 23730
rect 22468 23666 22520 23672
rect 22652 23724 22704 23730
rect 22652 23666 22704 23672
rect 22744 23724 22796 23730
rect 22744 23666 22796 23672
rect 22836 23724 22888 23730
rect 22836 23666 22888 23672
rect 21824 23656 21876 23662
rect 21824 23598 21876 23604
rect 21272 23520 21324 23526
rect 21272 23462 21324 23468
rect 21836 23322 21864 23598
rect 22112 23322 22140 23666
rect 21824 23316 21876 23322
rect 21824 23258 21876 23264
rect 22100 23316 22152 23322
rect 22100 23258 22152 23264
rect 21456 22976 21508 22982
rect 21456 22918 21508 22924
rect 21548 22976 21600 22982
rect 21548 22918 21600 22924
rect 21180 22772 21232 22778
rect 21180 22714 21232 22720
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 21468 22506 21496 22918
rect 21560 22778 21588 22918
rect 21548 22772 21600 22778
rect 21548 22714 21600 22720
rect 22204 22642 22232 23666
rect 22480 23322 22508 23666
rect 22664 23322 22692 23666
rect 22756 23526 22784 23666
rect 22744 23520 22796 23526
rect 22744 23462 22796 23468
rect 22468 23316 22520 23322
rect 22468 23258 22520 23264
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22848 23118 22876 23666
rect 22836 23112 22888 23118
rect 22756 23060 22836 23066
rect 22756 23054 22888 23060
rect 22756 23038 22876 23054
rect 22940 23050 22968 24006
rect 23216 23526 23244 24550
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23204 23520 23256 23526
rect 23204 23462 23256 23468
rect 23032 23186 23060 23462
rect 23216 23322 23244 23462
rect 23204 23316 23256 23322
rect 23204 23258 23256 23264
rect 23020 23180 23072 23186
rect 23020 23122 23072 23128
rect 22928 23044 22980 23050
rect 22756 22982 22784 23038
rect 22928 22986 22980 22992
rect 22468 22976 22520 22982
rect 22468 22918 22520 22924
rect 22744 22976 22796 22982
rect 22744 22918 22796 22924
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 22376 22568 22428 22574
rect 22376 22510 22428 22516
rect 21456 22500 21508 22506
rect 21456 22442 21508 22448
rect 20904 22228 20956 22234
rect 20904 22170 20956 22176
rect 21744 22098 21772 22510
rect 21732 22092 21784 22098
rect 22388 22094 22416 22510
rect 21732 22034 21784 22040
rect 22204 22066 22416 22094
rect 19524 22024 19576 22030
rect 19524 21966 19576 21972
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19432 21480 19484 21486
rect 19432 21422 19484 21428
rect 19708 21412 19760 21418
rect 19708 21354 19760 21360
rect 19720 20942 19748 21354
rect 20088 21078 20116 21966
rect 21744 21690 21772 22034
rect 22204 21962 22232 22066
rect 22480 21962 22508 22918
rect 22848 22778 22876 22918
rect 22836 22772 22888 22778
rect 22836 22714 22888 22720
rect 22940 22658 22968 22986
rect 23032 22778 23060 23122
rect 23112 23112 23164 23118
rect 23216 23089 23244 23258
rect 23112 23054 23164 23060
rect 23202 23080 23258 23089
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 22664 22630 22968 22658
rect 22572 22098 22600 22578
rect 22560 22092 22612 22098
rect 22560 22034 22612 22040
rect 22192 21956 22244 21962
rect 22192 21898 22244 21904
rect 22468 21956 22520 21962
rect 22468 21898 22520 21904
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 20628 21548 20680 21554
rect 20628 21490 20680 21496
rect 20444 21140 20496 21146
rect 20444 21082 20496 21088
rect 20076 21072 20128 21078
rect 20076 21014 20128 21020
rect 19708 20936 19760 20942
rect 19708 20878 19760 20884
rect 20260 20936 20312 20942
rect 20260 20878 20312 20884
rect 20168 20800 20220 20806
rect 20168 20742 20220 20748
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 20180 20330 20208 20742
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 19076 19446 19104 19858
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 17684 19440 17736 19446
rect 19064 19440 19116 19446
rect 17684 19382 17736 19388
rect 17696 19242 17724 19382
rect 17868 19372 17920 19378
rect 18340 19366 18552 19394
rect 19064 19382 19116 19388
rect 17920 19320 18000 19334
rect 17868 19314 18000 19320
rect 17880 19306 18000 19314
rect 18340 19310 18368 19366
rect 18524 19334 18552 19366
rect 19076 19334 19104 19382
rect 19352 19378 19380 19790
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19984 19712 20036 19718
rect 19984 19654 20036 19660
rect 19444 19394 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19444 19378 19656 19394
rect 19996 19378 20024 19654
rect 20180 19514 20208 20266
rect 20272 20262 20300 20878
rect 20456 20398 20484 21082
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 19922 20300 20198
rect 20260 19916 20312 19922
rect 20260 19858 20312 19864
rect 20640 19854 20668 21490
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 20732 19854 20760 21286
rect 21836 21146 21864 21286
rect 21824 21140 21876 21146
rect 21824 21082 21876 21088
rect 22480 20058 22508 21898
rect 22572 21690 22600 22034
rect 22560 21684 22612 21690
rect 22560 21626 22612 21632
rect 22560 20936 22612 20942
rect 22664 20924 22692 22630
rect 22836 22568 22888 22574
rect 22836 22510 22888 22516
rect 22848 21706 22876 22510
rect 23124 22438 23152 23054
rect 23202 23015 23258 23024
rect 23112 22432 23164 22438
rect 23112 22374 23164 22380
rect 22612 20896 22692 20924
rect 22756 21678 22876 21706
rect 22560 20878 22612 20884
rect 22572 20602 22600 20878
rect 22756 20602 22784 21678
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 22848 20942 22876 21558
rect 23124 21350 23152 22374
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 21010 23152 21286
rect 23112 21004 23164 21010
rect 23112 20946 23164 20952
rect 23216 20942 23244 23015
rect 23308 22710 23336 25162
rect 23676 24682 23704 25230
rect 23768 24954 23796 25434
rect 24780 25362 24808 26930
rect 24872 25498 24900 28358
rect 25424 27470 25452 28426
rect 26240 28416 26292 28422
rect 26240 28358 26292 28364
rect 26252 27674 26280 28358
rect 26344 27674 26372 28494
rect 26240 27668 26292 27674
rect 26240 27610 26292 27616
rect 26332 27668 26384 27674
rect 26332 27610 26384 27616
rect 25412 27464 25464 27470
rect 25412 27406 25464 27412
rect 25964 27464 26016 27470
rect 25964 27406 26016 27412
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 25044 27328 25096 27334
rect 25044 27270 25096 27276
rect 25872 27328 25924 27334
rect 25872 27270 25924 27276
rect 25056 26790 25084 27270
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25148 27033 25176 27066
rect 25884 27062 25912 27270
rect 25228 27056 25280 27062
rect 25134 27024 25190 27033
rect 25412 27056 25464 27062
rect 25280 27016 25412 27044
rect 25228 26998 25280 27004
rect 25412 26998 25464 27004
rect 25872 27056 25924 27062
rect 25872 26998 25924 27004
rect 25134 26959 25136 26968
rect 25188 26959 25190 26968
rect 25136 26930 25188 26936
rect 25688 26920 25740 26926
rect 25686 26888 25688 26897
rect 25740 26888 25742 26897
rect 25686 26823 25742 26832
rect 25044 26784 25096 26790
rect 25044 26726 25096 26732
rect 25700 26382 25728 26823
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25884 26382 25912 26726
rect 25976 26586 26004 27406
rect 26160 27130 26188 27406
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26424 27396 26476 27402
rect 26424 27338 26476 27344
rect 26344 27130 26372 27338
rect 26148 27124 26200 27130
rect 26148 27066 26200 27072
rect 26240 27124 26292 27130
rect 26240 27066 26292 27072
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26056 26988 26108 26994
rect 26056 26930 26108 26936
rect 25964 26580 26016 26586
rect 25964 26522 26016 26528
rect 26068 26382 26096 26930
rect 25688 26376 25740 26382
rect 25688 26318 25740 26324
rect 25872 26376 25924 26382
rect 25872 26318 25924 26324
rect 26056 26376 26108 26382
rect 26056 26318 26108 26324
rect 26252 26314 26280 27066
rect 26330 27024 26386 27033
rect 26436 27010 26464 27338
rect 26386 26982 26464 27010
rect 26330 26959 26332 26968
rect 26384 26959 26386 26968
rect 26332 26930 26384 26936
rect 26528 26858 26556 28630
rect 26988 28626 27016 28970
rect 26976 28620 27028 28626
rect 26976 28562 27028 28568
rect 27080 28558 27108 29514
rect 27988 28960 28040 28966
rect 27988 28902 28040 28908
rect 28000 28558 28028 28902
rect 28368 28762 28396 29582
rect 29196 29510 29224 29582
rect 29184 29504 29236 29510
rect 29184 29446 29236 29452
rect 29840 29306 29868 29650
rect 30380 29572 30432 29578
rect 30380 29514 30432 29520
rect 30196 29504 30248 29510
rect 30196 29446 30248 29452
rect 29828 29300 29880 29306
rect 29828 29242 29880 29248
rect 28540 28960 28592 28966
rect 28540 28902 28592 28908
rect 28356 28756 28408 28762
rect 28356 28698 28408 28704
rect 28264 28688 28316 28694
rect 28184 28648 28264 28676
rect 28184 28642 28212 28648
rect 28092 28626 28212 28642
rect 28264 28630 28316 28636
rect 28080 28620 28212 28626
rect 28132 28614 28212 28620
rect 28080 28562 28132 28568
rect 27068 28552 27120 28558
rect 27068 28494 27120 28500
rect 27988 28552 28040 28558
rect 27988 28494 28040 28500
rect 28172 28552 28224 28558
rect 28172 28494 28224 28500
rect 28080 28484 28132 28490
rect 28080 28426 28132 28432
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27724 28218 27752 28358
rect 28092 28218 28120 28426
rect 27712 28212 27764 28218
rect 27712 28154 27764 28160
rect 28080 28212 28132 28218
rect 28080 28154 28132 28160
rect 27528 28076 27580 28082
rect 27528 28018 27580 28024
rect 27712 28076 27764 28082
rect 27712 28018 27764 28024
rect 27540 27402 27568 28018
rect 27724 27538 27752 28018
rect 28184 28014 28212 28494
rect 28552 28490 28580 28902
rect 29840 28626 29868 29242
rect 30208 28966 30236 29446
rect 30392 29306 30420 29514
rect 30380 29300 30432 29306
rect 30380 29242 30432 29248
rect 30196 28960 30248 28966
rect 30196 28902 30248 28908
rect 29828 28620 29880 28626
rect 29828 28562 29880 28568
rect 28540 28484 28592 28490
rect 28540 28426 28592 28432
rect 28172 28008 28224 28014
rect 28172 27950 28224 27956
rect 27712 27532 27764 27538
rect 27712 27474 27764 27480
rect 28552 27470 28580 28426
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 27528 27396 27580 27402
rect 27528 27338 27580 27344
rect 28552 27130 28580 27406
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 29104 27130 29132 27270
rect 29840 27130 29868 28562
rect 30208 28082 30236 28902
rect 31036 28762 31064 30126
rect 31864 30054 31892 30194
rect 33888 30122 33916 36110
rect 34336 36100 34388 36106
rect 34336 36042 34388 36048
rect 34348 35737 34376 36042
rect 34334 35728 34390 35737
rect 34334 35663 34390 35672
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34612 33924 34664 33930
rect 34612 33866 34664 33872
rect 34624 33561 34652 33866
rect 34704 33856 34756 33862
rect 34704 33798 34756 33804
rect 34610 33552 34666 33561
rect 34610 33487 34666 33496
rect 34520 31816 34572 31822
rect 34520 31758 34572 31764
rect 34060 31680 34112 31686
rect 34060 31622 34112 31628
rect 34072 31385 34100 31622
rect 34058 31376 34114 31385
rect 34058 31311 34114 31320
rect 34428 30592 34480 30598
rect 34428 30534 34480 30540
rect 33876 30116 33928 30122
rect 33876 30058 33928 30064
rect 34440 30054 34468 30534
rect 31852 30048 31904 30054
rect 31852 29990 31904 29996
rect 34244 30048 34296 30054
rect 34244 29990 34296 29996
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 31668 29640 31720 29646
rect 31668 29582 31720 29588
rect 31024 28756 31076 28762
rect 31024 28698 31076 28704
rect 31680 28694 31708 29582
rect 31864 29578 31892 29990
rect 34256 29782 34284 29990
rect 34244 29776 34296 29782
rect 34244 29718 34296 29724
rect 32220 29708 32272 29714
rect 32220 29650 32272 29656
rect 31852 29572 31904 29578
rect 31852 29514 31904 29520
rect 32232 28694 32260 29650
rect 32588 29640 32640 29646
rect 32588 29582 32640 29588
rect 32600 29306 32628 29582
rect 32588 29300 32640 29306
rect 32588 29242 32640 29248
rect 31668 28688 31720 28694
rect 31668 28630 31720 28636
rect 32220 28688 32272 28694
rect 32220 28630 32272 28636
rect 30288 28484 30340 28490
rect 30288 28426 30340 28432
rect 30300 28218 30328 28426
rect 30288 28212 30340 28218
rect 30288 28154 30340 28160
rect 31680 28082 31708 28630
rect 32312 28620 32364 28626
rect 32312 28562 32364 28568
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 32036 28552 32088 28558
rect 32036 28494 32088 28500
rect 31772 28422 31800 28494
rect 31760 28416 31812 28422
rect 31760 28358 31812 28364
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 31668 28076 31720 28082
rect 31668 28018 31720 28024
rect 31772 27878 31800 28358
rect 32048 28014 32076 28494
rect 32324 28218 32352 28562
rect 32312 28212 32364 28218
rect 32312 28154 32364 28160
rect 32036 28008 32088 28014
rect 32036 27950 32088 27956
rect 31300 27872 31352 27878
rect 31300 27814 31352 27820
rect 31760 27872 31812 27878
rect 31760 27814 31812 27820
rect 32312 27872 32364 27878
rect 32312 27814 32364 27820
rect 28540 27124 28592 27130
rect 28540 27066 28592 27072
rect 29092 27124 29144 27130
rect 29092 27066 29144 27072
rect 29644 27124 29696 27130
rect 29644 27066 29696 27072
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 26792 26988 26844 26994
rect 26792 26930 26844 26936
rect 27068 26988 27120 26994
rect 27068 26930 27120 26936
rect 27252 26988 27304 26994
rect 27252 26930 27304 26936
rect 26804 26897 26832 26930
rect 26790 26888 26846 26897
rect 26516 26852 26568 26858
rect 26790 26823 26846 26832
rect 26516 26794 26568 26800
rect 27080 26314 27108 26930
rect 27264 26382 27292 26930
rect 29656 26926 29684 27066
rect 31312 26994 31340 27814
rect 31772 27674 31800 27814
rect 31760 27668 31812 27674
rect 31760 27610 31812 27616
rect 31668 27532 31720 27538
rect 31668 27474 31720 27480
rect 32128 27532 32180 27538
rect 32128 27474 32180 27480
rect 31484 27328 31536 27334
rect 31484 27270 31536 27276
rect 31496 27130 31524 27270
rect 31484 27124 31536 27130
rect 31484 27066 31536 27072
rect 31680 26994 31708 27474
rect 32140 27130 32168 27474
rect 32128 27124 32180 27130
rect 32128 27066 32180 27072
rect 32324 26994 32352 27814
rect 32600 27538 32628 29242
rect 34058 29200 34114 29209
rect 34058 29135 34114 29144
rect 33048 28960 33100 28966
rect 33048 28902 33100 28908
rect 33060 28762 33088 28902
rect 33048 28756 33100 28762
rect 33048 28698 33100 28704
rect 34072 28626 34100 29135
rect 34060 28620 34112 28626
rect 34060 28562 34112 28568
rect 34440 28422 34468 29990
rect 34532 29850 34560 31758
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 34716 29306 34744 33798
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34704 29300 34756 29306
rect 34704 29242 34756 29248
rect 34796 29232 34848 29238
rect 34796 29174 34848 29180
rect 34808 28762 34836 29174
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28756 34848 28762
rect 34796 28698 34848 28704
rect 34520 28552 34572 28558
rect 34520 28494 34572 28500
rect 32772 28416 32824 28422
rect 32772 28358 32824 28364
rect 34428 28416 34480 28422
rect 34428 28358 34480 28364
rect 32784 28014 32812 28358
rect 32772 28008 32824 28014
rect 32772 27950 32824 27956
rect 34440 27878 34468 28358
rect 34428 27872 34480 27878
rect 34428 27814 34480 27820
rect 34440 27554 34468 27814
rect 34532 27674 34560 28494
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34520 27668 34572 27674
rect 34520 27610 34572 27616
rect 32588 27532 32640 27538
rect 34440 27526 34560 27554
rect 32588 27474 32640 27480
rect 32600 27130 32628 27474
rect 34532 27470 34560 27526
rect 34520 27464 34572 27470
rect 34520 27406 34572 27412
rect 32588 27124 32640 27130
rect 32588 27066 32640 27072
rect 31300 26988 31352 26994
rect 31300 26930 31352 26936
rect 31668 26988 31720 26994
rect 31668 26930 31720 26936
rect 32312 26988 32364 26994
rect 32312 26930 32364 26936
rect 29644 26920 29696 26926
rect 29644 26862 29696 26868
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 27068 26308 27120 26314
rect 27068 26250 27120 26256
rect 26332 26240 26384 26246
rect 26332 26182 26384 26188
rect 26344 25974 26372 26182
rect 26332 25968 26384 25974
rect 26332 25910 26384 25916
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 24860 25492 24912 25498
rect 24860 25434 24912 25440
rect 26160 25362 26188 25842
rect 24768 25356 24820 25362
rect 24768 25298 24820 25304
rect 26148 25356 26200 25362
rect 26148 25298 26200 25304
rect 24032 25288 24084 25294
rect 24032 25230 24084 25236
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24860 25288 24912 25294
rect 24860 25230 24912 25236
rect 25780 25288 25832 25294
rect 25780 25230 25832 25236
rect 25964 25288 26016 25294
rect 25964 25230 26016 25236
rect 23756 24948 23808 24954
rect 23756 24890 23808 24896
rect 24044 24818 24072 25230
rect 24308 25152 24360 25158
rect 24308 25094 24360 25100
rect 24320 24818 24348 25094
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 24032 24812 24084 24818
rect 24032 24754 24084 24760
rect 24308 24812 24360 24818
rect 24308 24754 24360 24760
rect 23664 24676 23716 24682
rect 23664 24618 23716 24624
rect 23388 24064 23440 24070
rect 23388 24006 23440 24012
rect 23400 23798 23428 24006
rect 23676 23866 23704 24618
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23296 22704 23348 22710
rect 23296 22646 23348 22652
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23400 22234 23428 22374
rect 23388 22228 23440 22234
rect 23388 22170 23440 22176
rect 23296 21344 23348 21350
rect 23296 21286 23348 21292
rect 22836 20936 22888 20942
rect 22836 20878 22888 20884
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 22848 20602 22876 20878
rect 22928 20868 22980 20874
rect 22928 20810 22980 20816
rect 22560 20596 22612 20602
rect 22560 20538 22612 20544
rect 22744 20596 22796 20602
rect 22744 20538 22796 20544
rect 22836 20596 22888 20602
rect 22836 20538 22888 20544
rect 20996 20052 21048 20058
rect 20996 19994 21048 20000
rect 22468 20052 22520 20058
rect 22468 19994 22520 20000
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20720 19848 20772 19854
rect 20720 19790 20772 19796
rect 20640 19514 20668 19790
rect 20824 19530 20852 19858
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20168 19508 20220 19514
rect 20168 19450 20220 19456
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20732 19502 20852 19530
rect 20732 19446 20760 19502
rect 20720 19440 20772 19446
rect 20720 19382 20772 19388
rect 20916 19378 20944 19790
rect 18524 19310 18736 19334
rect 17684 19236 17736 19242
rect 17736 19196 17908 19224
rect 17684 19178 17736 19184
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 17316 18352 17368 18358
rect 17316 18294 17368 18300
rect 17406 18320 17462 18329
rect 17406 18255 17408 18264
rect 17460 18255 17462 18264
rect 17500 18284 17552 18290
rect 17408 18226 17460 18232
rect 17500 18226 17552 18232
rect 17592 18284 17644 18290
rect 17592 18226 17644 18232
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17408 18148 17460 18154
rect 17408 18090 17460 18096
rect 17040 17536 17092 17542
rect 17040 17478 17092 17484
rect 16948 17332 17000 17338
rect 16948 17274 17000 17280
rect 17420 17270 17448 18090
rect 17512 17882 17540 18226
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17604 17338 17632 18226
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17592 17332 17644 17338
rect 17592 17274 17644 17280
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16960 16794 16988 17138
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16396 16040 16448 16046
rect 16396 15982 16448 15988
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15016 15496 15068 15502
rect 14752 15444 15016 15450
rect 14752 15438 15068 15444
rect 14752 15422 15056 15438
rect 14752 15366 14780 15422
rect 14740 15360 14792 15366
rect 14740 15302 14792 15308
rect 15120 15026 15148 15574
rect 16684 15570 16712 16526
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 16672 15564 16724 15570
rect 16672 15506 16724 15512
rect 15304 15094 15332 15506
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 16132 15026 16160 15438
rect 16672 15360 16724 15366
rect 16672 15302 16724 15308
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 14618 14780 14894
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 14936 14550 14964 14962
rect 16580 14952 16632 14958
rect 16580 14894 16632 14900
rect 16592 14618 16620 14894
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 14924 14544 14976 14550
rect 14924 14486 14976 14492
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 14556 14068 14608 14074
rect 14556 14010 14608 14016
rect 15396 13938 15424 14214
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 14924 13796 14976 13802
rect 14924 13738 14976 13744
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 12912 13246 13032 13274
rect 13004 12986 13032 13246
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 12992 12980 13044 12986
rect 12992 12922 13044 12928
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12820 12374 12848 12786
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12820 11898 12848 12174
rect 13556 11898 13584 13126
rect 13832 12986 13860 13466
rect 14200 13190 14228 13670
rect 14936 13394 14964 13738
rect 15396 13530 15424 13874
rect 15844 13864 15896 13870
rect 15844 13806 15896 13812
rect 15384 13524 15436 13530
rect 15384 13466 15436 13472
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14280 13252 14332 13258
rect 14280 13194 14332 13200
rect 14556 13252 14608 13258
rect 14556 13194 14608 13200
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14200 12986 14228 13126
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 14188 12980 14240 12986
rect 14188 12922 14240 12928
rect 14292 12850 14320 13194
rect 14568 12986 14596 13194
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 14280 12844 14332 12850
rect 14280 12786 14332 12792
rect 13924 11898 13952 12786
rect 14292 12646 14320 12786
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 14568 12238 14596 12922
rect 14936 12850 14964 13330
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14832 12776 14884 12782
rect 14832 12718 14884 12724
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 14844 12238 14872 12718
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15292 12640 15344 12646
rect 15292 12582 15344 12588
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 12808 11892 12860 11898
rect 12808 11834 12860 11840
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13924 11762 13952 11834
rect 14844 11830 14872 12174
rect 15120 11898 15148 12582
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15108 11892 15160 11898
rect 15108 11834 15160 11840
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 15212 11762 15240 12038
rect 15304 11762 15332 12582
rect 15580 11898 15608 12718
rect 15672 12714 15700 12854
rect 15660 12708 15712 12714
rect 15660 12650 15712 12656
rect 15672 12306 15700 12650
rect 15660 12300 15712 12306
rect 15660 12242 15712 12248
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 13912 11756 13964 11762
rect 13912 11698 13964 11704
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 13004 11558 13032 11698
rect 12992 11552 13044 11558
rect 12992 11494 13044 11500
rect 13004 11354 13032 11494
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 15672 11082 15700 12106
rect 15764 11354 15792 13466
rect 15856 13394 15884 13806
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15948 12850 15976 14214
rect 16120 14068 16172 14074
rect 16120 14010 16172 14016
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15948 12714 15976 12786
rect 15936 12708 15988 12714
rect 15936 12650 15988 12656
rect 15948 12102 15976 12650
rect 16132 12434 16160 14010
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 16224 12850 16252 13466
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16316 12986 16344 13262
rect 16304 12980 16356 12986
rect 16304 12922 16356 12928
rect 16684 12918 16712 15302
rect 16776 14482 16804 15846
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16868 15026 16896 15370
rect 17052 15366 17080 15846
rect 17040 15360 17092 15366
rect 17040 15302 17092 15308
rect 17224 15360 17276 15366
rect 17224 15302 17276 15308
rect 16856 15020 16908 15026
rect 16856 14962 16908 14968
rect 16764 14476 16816 14482
rect 16764 14418 16816 14424
rect 16868 13938 16896 14962
rect 17236 14822 17264 15302
rect 17328 15094 17356 17138
rect 17696 16998 17724 17682
rect 17776 17536 17828 17542
rect 17776 17478 17828 17484
rect 17788 17202 17816 17478
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17408 16992 17460 16998
rect 17408 16934 17460 16940
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17420 16590 17448 16934
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17788 16114 17816 16390
rect 17776 16108 17828 16114
rect 17776 16050 17828 16056
rect 17880 15978 17908 19196
rect 17972 16114 18000 19306
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18420 19304 18472 19310
rect 18524 19306 18748 19310
rect 18420 19246 18472 19252
rect 18696 19304 18748 19306
rect 18696 19246 18748 19252
rect 18984 19306 19104 19334
rect 19340 19372 19392 19378
rect 19444 19372 19668 19378
rect 19444 19366 19616 19372
rect 19340 19314 19392 19320
rect 19616 19314 19668 19320
rect 19984 19372 20036 19378
rect 19984 19314 20036 19320
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 18064 16794 18092 19246
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18052 16788 18104 16794
rect 18052 16730 18104 16736
rect 18156 16590 18184 17138
rect 18144 16584 18196 16590
rect 18144 16526 18196 16532
rect 18340 16250 18368 19110
rect 18432 18748 18460 19246
rect 18984 18902 19012 19306
rect 19064 19236 19116 19242
rect 19064 19178 19116 19184
rect 18604 18896 18656 18902
rect 18604 18838 18656 18844
rect 18972 18896 19024 18902
rect 18972 18838 19024 18844
rect 18512 18760 18564 18766
rect 18432 18720 18512 18748
rect 18512 18702 18564 18708
rect 18524 18222 18552 18702
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18340 16114 18368 16186
rect 18432 16114 18460 16730
rect 18616 16250 18644 18838
rect 19076 18766 19104 19178
rect 19352 18834 19380 19314
rect 19628 18970 19656 19314
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 20916 18766 20944 19314
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20720 18692 20772 18698
rect 20720 18634 20772 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19338 18320 19394 18329
rect 19338 18255 19394 18264
rect 19708 18284 19760 18290
rect 19352 17678 19380 18255
rect 19708 18226 19760 18232
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 19720 17746 19748 18226
rect 20364 17746 20392 18226
rect 20732 18154 20760 18634
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 21008 17814 21036 19994
rect 22756 19854 22784 20538
rect 22836 20256 22888 20262
rect 22940 20244 22968 20810
rect 22888 20216 22968 20244
rect 22836 20198 22888 20204
rect 21916 19848 21968 19854
rect 21916 19790 21968 19796
rect 22744 19848 22796 19854
rect 22744 19790 22796 19796
rect 21088 19780 21140 19786
rect 21088 19722 21140 19728
rect 21100 19378 21128 19722
rect 21548 19508 21600 19514
rect 21548 19450 21600 19456
rect 21560 19394 21588 19450
rect 21560 19378 21680 19394
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 21560 19372 21692 19378
rect 21560 19366 21640 19372
rect 21100 18698 21128 19314
rect 21364 18760 21416 18766
rect 21364 18702 21416 18708
rect 21088 18692 21140 18698
rect 21088 18634 21140 18640
rect 21376 18290 21404 18702
rect 21560 18698 21588 19366
rect 21640 19314 21692 19320
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21744 18426 21772 19110
rect 21928 18902 21956 19790
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22112 19310 22140 19654
rect 22756 19514 22784 19790
rect 22848 19718 22876 20198
rect 22928 19916 22980 19922
rect 22928 19858 22980 19864
rect 22836 19712 22888 19718
rect 22836 19654 22888 19660
rect 22744 19508 22796 19514
rect 22744 19450 22796 19456
rect 22940 19378 22968 19858
rect 23308 19786 23336 21286
rect 23400 20482 23428 22170
rect 23768 22094 23796 24754
rect 24308 23520 24360 23526
rect 24308 23462 24360 23468
rect 24320 23118 24348 23462
rect 24412 23322 24440 25230
rect 24872 24954 24900 25230
rect 24860 24948 24912 24954
rect 24860 24890 24912 24896
rect 25792 24886 25820 25230
rect 25780 24880 25832 24886
rect 25780 24822 25832 24828
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 24492 23724 24544 23730
rect 24492 23666 24544 23672
rect 24400 23316 24452 23322
rect 24400 23258 24452 23264
rect 24504 23118 24532 23666
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24872 23322 24900 23462
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24872 23202 24900 23258
rect 24780 23174 24900 23202
rect 24780 23118 24808 23174
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24308 23112 24360 23118
rect 24308 23054 24360 23060
rect 24492 23112 24544 23118
rect 24492 23054 24544 23060
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 23584 22066 23796 22094
rect 23584 21690 23612 22066
rect 23572 21684 23624 21690
rect 23572 21626 23624 21632
rect 23584 21146 23612 21626
rect 24044 21146 24072 23054
rect 24504 22982 24532 23054
rect 24492 22976 24544 22982
rect 24492 22918 24544 22924
rect 24504 22778 24532 22918
rect 24872 22778 24900 23054
rect 24492 22772 24544 22778
rect 24492 22714 24544 22720
rect 24860 22772 24912 22778
rect 24860 22714 24912 22720
rect 24964 21146 24992 24754
rect 25596 24676 25648 24682
rect 25596 24618 25648 24624
rect 25608 24206 25636 24618
rect 25596 24200 25648 24206
rect 25596 24142 25648 24148
rect 25608 23798 25636 24142
rect 25044 23792 25096 23798
rect 25044 23734 25096 23740
rect 25596 23792 25648 23798
rect 25596 23734 25648 23740
rect 25056 22574 25084 23734
rect 25792 23186 25820 24822
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25884 24410 25912 24754
rect 25976 24750 26004 25230
rect 25964 24744 26016 24750
rect 25964 24686 26016 24692
rect 25872 24404 25924 24410
rect 25872 24346 25924 24352
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25044 22568 25096 22574
rect 25044 22510 25096 22516
rect 26056 22094 26108 22098
rect 26160 22094 26188 25298
rect 27080 24342 27108 26250
rect 27264 26042 27292 26318
rect 27252 26036 27304 26042
rect 27252 25978 27304 25984
rect 29552 25968 29604 25974
rect 29656 25956 29684 26862
rect 31312 26246 31340 26930
rect 30656 26240 30708 26246
rect 30656 26182 30708 26188
rect 31300 26240 31352 26246
rect 31300 26182 31352 26188
rect 29604 25928 29684 25956
rect 29552 25910 29604 25916
rect 27160 25900 27212 25906
rect 27160 25842 27212 25848
rect 27172 24614 27200 25842
rect 27344 25832 27396 25838
rect 27344 25774 27396 25780
rect 27356 25362 27384 25774
rect 28080 25764 28132 25770
rect 28080 25706 28132 25712
rect 27344 25356 27396 25362
rect 27344 25298 27396 25304
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27344 25152 27396 25158
rect 27344 25094 27396 25100
rect 27160 24608 27212 24614
rect 27160 24550 27212 24556
rect 27068 24336 27120 24342
rect 27068 24278 27120 24284
rect 26976 24200 27028 24206
rect 26976 24142 27028 24148
rect 26988 23866 27016 24142
rect 27172 23866 27200 24550
rect 27356 24274 27384 25094
rect 27632 24274 27660 25230
rect 27344 24268 27396 24274
rect 27344 24210 27396 24216
rect 27620 24268 27672 24274
rect 27620 24210 27672 24216
rect 27436 24200 27488 24206
rect 27436 24142 27488 24148
rect 26976 23860 27028 23866
rect 26976 23802 27028 23808
rect 27160 23860 27212 23866
rect 27160 23802 27212 23808
rect 27448 23798 27476 24142
rect 27816 24138 27844 25230
rect 28092 24410 28120 25706
rect 29656 24954 29684 25928
rect 30564 25968 30616 25974
rect 30564 25910 30616 25916
rect 30576 25498 30604 25910
rect 30564 25492 30616 25498
rect 30564 25434 30616 25440
rect 30668 25158 30696 26182
rect 31680 26042 31708 26930
rect 31668 26036 31720 26042
rect 31668 25978 31720 25984
rect 31852 25832 31904 25838
rect 31852 25774 31904 25780
rect 32220 25832 32272 25838
rect 32220 25774 32272 25780
rect 31760 25764 31812 25770
rect 31760 25706 31812 25712
rect 31772 25294 31800 25706
rect 31864 25294 31892 25774
rect 32232 25498 32260 25774
rect 32220 25492 32272 25498
rect 32220 25434 32272 25440
rect 32324 25362 32352 26930
rect 32600 26586 32628 27066
rect 32588 26580 32640 26586
rect 32588 26522 32640 26528
rect 34532 26382 34560 27406
rect 34794 27024 34850 27033
rect 34704 26988 34756 26994
rect 34794 26959 34796 26968
rect 34704 26930 34756 26936
rect 34848 26959 34850 26968
rect 34796 26930 34848 26936
rect 34716 26586 34744 26930
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34704 26580 34756 26586
rect 34704 26522 34756 26528
rect 34520 26376 34572 26382
rect 34520 26318 34572 26324
rect 33048 26308 33100 26314
rect 33048 26250 33100 26256
rect 33060 26042 33088 26250
rect 33048 26036 33100 26042
rect 33048 25978 33100 25984
rect 34532 25702 34560 26318
rect 34520 25696 34572 25702
rect 34520 25638 34572 25644
rect 32312 25356 32364 25362
rect 32312 25298 32364 25304
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31852 25288 31904 25294
rect 31852 25230 31904 25236
rect 32956 25288 33008 25294
rect 32956 25230 33008 25236
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 29644 24948 29696 24954
rect 29644 24890 29696 24896
rect 28080 24404 28132 24410
rect 28080 24346 28132 24352
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 28632 24200 28684 24206
rect 28632 24142 28684 24148
rect 27804 24132 27856 24138
rect 27804 24074 27856 24080
rect 27988 24132 28040 24138
rect 27988 24074 28040 24080
rect 27528 24064 27580 24070
rect 27528 24006 27580 24012
rect 27436 23792 27488 23798
rect 27436 23734 27488 23740
rect 27540 23526 27568 24006
rect 27816 23798 27844 24074
rect 27804 23792 27856 23798
rect 27804 23734 27856 23740
rect 28000 23662 28028 24074
rect 28644 23866 28672 24142
rect 28736 23866 28764 24278
rect 29656 24274 29684 24890
rect 29092 24268 29144 24274
rect 29092 24210 29144 24216
rect 29644 24268 29696 24274
rect 29644 24210 29696 24216
rect 29000 24200 29052 24206
rect 29000 24142 29052 24148
rect 28908 24064 28960 24070
rect 28908 24006 28960 24012
rect 28920 23866 28948 24006
rect 29012 23866 29040 24142
rect 29104 23866 29132 24210
rect 29368 24200 29420 24206
rect 29368 24142 29420 24148
rect 28632 23860 28684 23866
rect 28632 23802 28684 23808
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 28908 23860 28960 23866
rect 28908 23802 28960 23808
rect 29000 23860 29052 23866
rect 29000 23802 29052 23808
rect 29092 23860 29144 23866
rect 29092 23802 29144 23808
rect 28356 23792 28408 23798
rect 28408 23740 29132 23746
rect 28356 23734 29132 23740
rect 28368 23730 29132 23734
rect 29380 23730 29408 24142
rect 28368 23724 29144 23730
rect 28368 23718 29092 23724
rect 29092 23666 29144 23672
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 27988 23656 28040 23662
rect 27988 23598 28040 23604
rect 27252 23520 27304 23526
rect 27252 23462 27304 23468
rect 27528 23520 27580 23526
rect 27528 23462 27580 23468
rect 26240 22636 26292 22642
rect 26240 22578 26292 22584
rect 26252 22166 26280 22578
rect 26240 22160 26292 22166
rect 26240 22102 26292 22108
rect 26332 22160 26384 22166
rect 26384 22108 26464 22114
rect 26332 22102 26464 22108
rect 26056 22092 26188 22094
rect 26108 22066 26188 22092
rect 26344 22086 26464 22102
rect 27264 22098 27292 23462
rect 29656 22778 29684 24210
rect 30668 23526 30696 25094
rect 31772 24818 31800 25230
rect 31944 25152 31996 25158
rect 31944 25094 31996 25100
rect 31956 24818 31984 25094
rect 32968 24818 32996 25230
rect 34060 25220 34112 25226
rect 34060 25162 34112 25168
rect 34072 24857 34100 25162
rect 34152 24880 34204 24886
rect 34058 24848 34114 24857
rect 31760 24812 31812 24818
rect 31760 24754 31812 24760
rect 31944 24812 31996 24818
rect 31944 24754 31996 24760
rect 32956 24812 33008 24818
rect 34152 24822 34204 24828
rect 34058 24783 34114 24792
rect 32956 24754 33008 24760
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30852 23866 30880 24074
rect 30840 23860 30892 23866
rect 30840 23802 30892 23808
rect 30656 23520 30708 23526
rect 30656 23462 30708 23468
rect 29644 22772 29696 22778
rect 29644 22714 29696 22720
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 27620 22568 27672 22574
rect 27620 22510 27672 22516
rect 27528 22432 27580 22438
rect 27528 22374 27580 22380
rect 26056 22034 26108 22040
rect 26332 21480 26384 21486
rect 26332 21422 26384 21428
rect 26344 21146 26372 21422
rect 26436 21350 26464 22086
rect 26608 22092 26660 22098
rect 27252 22092 27304 22098
rect 26660 22052 26740 22080
rect 26608 22034 26660 22040
rect 26516 21888 26568 21894
rect 26516 21830 26568 21836
rect 26608 21888 26660 21894
rect 26608 21830 26660 21836
rect 26528 21554 26556 21830
rect 26620 21622 26648 21830
rect 26608 21616 26660 21622
rect 26608 21558 26660 21564
rect 26516 21548 26568 21554
rect 26516 21490 26568 21496
rect 26712 21418 26740 22052
rect 27252 22034 27304 22040
rect 26884 22024 26936 22030
rect 26884 21966 26936 21972
rect 27344 22024 27396 22030
rect 27540 22012 27568 22374
rect 27396 21984 27568 22012
rect 27344 21966 27396 21972
rect 26792 21956 26844 21962
rect 26792 21898 26844 21904
rect 26804 21690 26832 21898
rect 26896 21894 26924 21966
rect 27160 21956 27212 21962
rect 27160 21898 27212 21904
rect 26884 21888 26936 21894
rect 26884 21830 26936 21836
rect 27172 21690 27200 21898
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 26792 21684 26844 21690
rect 26792 21626 26844 21632
rect 27160 21684 27212 21690
rect 27160 21626 27212 21632
rect 26804 21554 26832 21626
rect 27540 21554 27568 21830
rect 26792 21548 26844 21554
rect 26792 21490 26844 21496
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 26700 21412 26752 21418
rect 26700 21354 26752 21360
rect 26424 21344 26476 21350
rect 26424 21286 26476 21292
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 24952 21140 25004 21146
rect 24952 21082 25004 21088
rect 26332 21140 26384 21146
rect 26332 21082 26384 21088
rect 23480 21004 23532 21010
rect 23480 20946 23532 20952
rect 23492 20602 23520 20946
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23400 20454 23520 20482
rect 23492 19836 23520 20454
rect 23584 20330 23612 21082
rect 25320 21072 25372 21078
rect 25320 21014 25372 21020
rect 24492 21004 24544 21010
rect 24492 20946 24544 20952
rect 23664 20936 23716 20942
rect 23664 20878 23716 20884
rect 23848 20936 23900 20942
rect 23848 20878 23900 20884
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 23676 20466 23704 20878
rect 23756 20868 23808 20874
rect 23756 20810 23808 20816
rect 23664 20460 23716 20466
rect 23664 20402 23716 20408
rect 23768 20398 23796 20810
rect 23860 20534 23888 20878
rect 23848 20528 23900 20534
rect 23848 20470 23900 20476
rect 23756 20392 23808 20398
rect 23756 20334 23808 20340
rect 23572 20324 23624 20330
rect 23572 20266 23624 20272
rect 24136 20058 24164 20878
rect 24504 20602 24532 20946
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24492 20596 24544 20602
rect 24492 20538 24544 20544
rect 24872 20262 24900 20878
rect 25332 20602 25360 21014
rect 25780 20936 25832 20942
rect 25780 20878 25832 20884
rect 25872 20936 25924 20942
rect 25872 20878 25924 20884
rect 25504 20800 25556 20806
rect 25504 20742 25556 20748
rect 25320 20596 25372 20602
rect 25320 20538 25372 20544
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24124 20052 24176 20058
rect 24124 19994 24176 20000
rect 25516 19922 25544 20742
rect 25792 20466 25820 20878
rect 25884 20806 25912 20878
rect 26436 20806 26464 21286
rect 26712 21146 26740 21354
rect 27540 21350 27568 21490
rect 27632 21350 27660 22510
rect 27896 22432 27948 22438
rect 27896 22374 27948 22380
rect 27908 22166 27936 22374
rect 27896 22160 27948 22166
rect 27896 22102 27948 22108
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27804 22024 27856 22030
rect 27804 21966 27856 21972
rect 27724 21690 27752 21966
rect 27712 21684 27764 21690
rect 27712 21626 27764 21632
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27620 21344 27672 21350
rect 27620 21286 27672 21292
rect 26700 21140 26752 21146
rect 26700 21082 26752 21088
rect 25872 20800 25924 20806
rect 25872 20742 25924 20748
rect 26424 20800 26476 20806
rect 26424 20742 26476 20748
rect 25780 20460 25832 20466
rect 25780 20402 25832 20408
rect 25884 20346 25912 20742
rect 25964 20460 26016 20466
rect 25964 20402 26016 20408
rect 25700 20318 25912 20346
rect 25596 20256 25648 20262
rect 25596 20198 25648 20204
rect 25504 19916 25556 19922
rect 25504 19858 25556 19864
rect 25608 19854 25636 20198
rect 23664 19848 23716 19854
rect 23492 19808 23664 19836
rect 23296 19780 23348 19786
rect 23296 19722 23348 19728
rect 23492 19514 23520 19808
rect 23664 19790 23716 19796
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 22928 19372 22980 19378
rect 22928 19314 22980 19320
rect 22100 19304 22152 19310
rect 22100 19246 22152 19252
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22560 19168 22612 19174
rect 22560 19110 22612 19116
rect 22204 18970 22232 19110
rect 22192 18964 22244 18970
rect 22192 18906 22244 18912
rect 21916 18896 21968 18902
rect 21916 18838 21968 18844
rect 22572 18834 22600 19110
rect 22560 18828 22612 18834
rect 22560 18770 22612 18776
rect 21824 18760 21876 18766
rect 21824 18702 21876 18708
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 21732 18420 21784 18426
rect 21732 18362 21784 18368
rect 21836 18290 21864 18702
rect 21364 18284 21416 18290
rect 21364 18226 21416 18232
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21376 17882 21404 18226
rect 21364 17876 21416 17882
rect 21364 17818 21416 17824
rect 20996 17808 21048 17814
rect 20996 17750 21048 17756
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 20352 17740 20404 17746
rect 20352 17682 20404 17688
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19432 17672 19484 17678
rect 19432 17614 19484 17620
rect 19444 17202 19472 17614
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19444 16794 19472 17138
rect 20640 17134 20668 17478
rect 21008 17338 21036 17750
rect 21836 17338 21864 18226
rect 20996 17332 21048 17338
rect 20996 17274 21048 17280
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21008 17134 21036 17274
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20996 17128 21048 17134
rect 20996 17070 21048 17076
rect 21640 17128 21692 17134
rect 21640 17070 21692 17076
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18604 16244 18656 16250
rect 18604 16186 18656 16192
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18420 16108 18472 16114
rect 18420 16050 18472 16056
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17880 15706 17908 15914
rect 17972 15910 18000 16050
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17972 15706 18000 15846
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 17316 15088 17368 15094
rect 17316 15030 17368 15036
rect 17512 15026 17540 15642
rect 18340 15638 18368 16050
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 17866 15464 17922 15473
rect 17866 15399 17922 15408
rect 17880 15366 17908 15399
rect 18432 15366 18460 16050
rect 18616 15434 18644 16186
rect 18708 16114 18736 16458
rect 19260 16250 19288 16526
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 19444 16250 19472 16390
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20640 16250 20668 17070
rect 21652 16658 21680 17070
rect 21640 16652 21692 16658
rect 21640 16594 21692 16600
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19340 16244 19392 16250
rect 19340 16186 19392 16192
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 18984 16114 19012 16186
rect 19352 16130 19380 16186
rect 19616 16176 19668 16182
rect 19536 16136 19616 16164
rect 19536 16130 19564 16136
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18972 16108 19024 16114
rect 19352 16102 19564 16130
rect 19616 16118 19668 16124
rect 18972 16050 19024 16056
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18984 15434 19012 15574
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 18604 15428 18656 15434
rect 18604 15370 18656 15376
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 14414 17264 14758
rect 18892 14618 18920 15302
rect 18984 15026 19012 15370
rect 19168 15094 19196 15438
rect 19352 15366 19380 15846
rect 19536 15706 19564 16102
rect 19892 16108 19944 16114
rect 19892 16050 19944 16056
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 19904 15910 19932 16050
rect 19892 15904 19944 15910
rect 19892 15846 19944 15852
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19996 15366 20024 16050
rect 20076 15972 20128 15978
rect 20076 15914 20128 15920
rect 20088 15434 20116 15914
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 21008 15366 21036 15846
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19156 15088 19208 15094
rect 19156 15030 19208 15036
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17224 14408 17276 14414
rect 17224 14350 17276 14356
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 17052 13326 17080 14214
rect 17420 13938 17448 14214
rect 17408 13932 17460 13938
rect 17408 13874 17460 13880
rect 17604 13462 17632 14418
rect 17684 13932 17736 13938
rect 17684 13874 17736 13880
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 12714 16896 12786
rect 16856 12708 16908 12714
rect 16856 12650 16908 12656
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 17224 12640 17276 12646
rect 17224 12582 17276 12588
rect 16040 12406 16160 12434
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 15752 11348 15804 11354
rect 15752 11290 15804 11296
rect 15856 11286 15884 12038
rect 15948 11354 15976 12038
rect 16040 11778 16068 12406
rect 16224 12186 16252 12582
rect 17236 12238 17264 12582
rect 17420 12306 17448 13126
rect 17512 12986 17540 13126
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17512 12782 17540 12922
rect 17500 12776 17552 12782
rect 17500 12718 17552 12724
rect 17604 12714 17632 13398
rect 17696 13326 17724 13874
rect 18892 13870 18920 14554
rect 18984 14482 19012 14962
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18972 14272 19024 14278
rect 18972 14214 19024 14220
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 17960 13184 18012 13190
rect 17880 13144 17960 13172
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17500 12368 17552 12374
rect 17500 12310 17552 12316
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 16132 12158 16252 12186
rect 17224 12232 17276 12238
rect 17276 12192 17356 12220
rect 17224 12174 17276 12180
rect 16132 11898 16160 12158
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16854 11792 16910 11801
rect 16040 11762 16160 11778
rect 16040 11756 16172 11762
rect 16040 11750 16120 11756
rect 16120 11698 16172 11704
rect 16580 11756 16632 11762
rect 16854 11727 16856 11736
rect 16580 11698 16632 11704
rect 16908 11727 16910 11736
rect 16856 11698 16908 11704
rect 16488 11688 16540 11694
rect 16488 11630 16540 11636
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11393 16344 11494
rect 16302 11384 16358 11393
rect 15936 11348 15988 11354
rect 16500 11354 16528 11630
rect 16302 11319 16358 11328
rect 16488 11348 16540 11354
rect 15936 11290 15988 11296
rect 16488 11290 16540 11296
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 12716 10532 12768 10538
rect 12716 10474 12768 10480
rect 15672 10062 15700 11018
rect 16500 10062 16528 11290
rect 16592 10062 16620 11698
rect 16672 10736 16724 10742
rect 16672 10678 16724 10684
rect 16684 10062 16712 10678
rect 16960 10146 16988 12038
rect 17224 11756 17276 11762
rect 17224 11698 17276 11704
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17144 10674 17172 11018
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 17236 10266 17264 11698
rect 17328 10742 17356 12192
rect 17512 11150 17540 12310
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17592 11552 17644 11558
rect 17592 11494 17644 11500
rect 17604 11257 17632 11494
rect 17696 11354 17724 12106
rect 17788 12102 17816 12310
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17590 11248 17646 11257
rect 17590 11183 17646 11192
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17604 10742 17632 11086
rect 17316 10736 17368 10742
rect 17316 10678 17368 10684
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17512 10266 17540 10610
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17500 10260 17552 10266
rect 17500 10202 17552 10208
rect 16960 10118 17080 10146
rect 17236 10130 17264 10202
rect 17052 10062 17080 10118
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16580 10056 16632 10062
rect 16580 9998 16632 10004
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 15672 9518 15700 9998
rect 16500 9586 16528 9998
rect 16488 9580 16540 9586
rect 16488 9522 16540 9528
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 16592 9382 16620 9998
rect 16684 9654 16712 9998
rect 16672 9648 16724 9654
rect 16672 9590 16724 9596
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8974 16620 9318
rect 16684 9178 16712 9590
rect 17236 9586 17264 10066
rect 17512 10062 17540 10202
rect 17696 10062 17724 11290
rect 17788 11014 17816 11698
rect 17880 11354 17908 13144
rect 17960 13126 18012 13132
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17972 12442 18000 12582
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18340 12322 18368 13194
rect 18432 12850 18460 13738
rect 18788 13728 18840 13734
rect 18788 13670 18840 13676
rect 18512 13388 18564 13394
rect 18512 13330 18564 13336
rect 18524 13190 18552 13330
rect 18800 13190 18828 13670
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18788 13184 18840 13190
rect 18788 13126 18840 13132
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18156 12294 18368 12322
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17776 11008 17828 11014
rect 17776 10950 17828 10956
rect 17788 10674 17816 10950
rect 17972 10674 18000 12038
rect 18064 11354 18092 12242
rect 18156 11830 18184 12294
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18144 11824 18196 11830
rect 18144 11766 18196 11772
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17776 10668 17828 10674
rect 17776 10610 17828 10616
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 18064 10554 18092 11290
rect 18142 11248 18198 11257
rect 18142 11183 18198 11192
rect 18156 11150 18184 11183
rect 18248 11150 18276 12174
rect 18340 11150 18368 12294
rect 18432 11150 18460 12786
rect 18892 12646 18920 13262
rect 18984 12918 19012 14214
rect 19352 13938 19380 14214
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19248 13932 19300 13938
rect 19248 13874 19300 13880
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19260 13530 19288 13874
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 19076 12986 19104 13262
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19168 12986 19196 13126
rect 19260 13002 19288 13466
rect 19352 13462 19380 13738
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19444 13326 19472 13874
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13410 19564 13806
rect 19996 13530 20024 15302
rect 20812 14952 20864 14958
rect 20812 14894 20864 14900
rect 20824 14822 20852 14894
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20074 14512 20130 14521
rect 20074 14447 20130 14456
rect 20456 14470 20760 14498
rect 20088 14278 20116 14447
rect 20456 14346 20484 14470
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20088 14006 20116 14214
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 20364 13802 20392 14214
rect 20456 14074 20484 14282
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 20548 13938 20576 14214
rect 20536 13932 20588 13938
rect 20536 13874 20588 13880
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19536 13382 20024 13410
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19338 13016 19394 13025
rect 19574 13019 19882 13028
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19156 12980 19208 12986
rect 19260 12974 19338 13002
rect 19338 12951 19394 12960
rect 19524 12980 19576 12986
rect 19156 12922 19208 12928
rect 19524 12922 19576 12928
rect 18972 12912 19024 12918
rect 18972 12854 19024 12860
rect 19076 12714 19104 12922
rect 19340 12912 19392 12918
rect 19536 12889 19564 12922
rect 19340 12854 19392 12860
rect 19522 12880 19578 12889
rect 19352 12782 19380 12854
rect 19522 12815 19578 12824
rect 19340 12776 19392 12782
rect 19340 12718 19392 12724
rect 19524 12776 19576 12782
rect 19524 12718 19576 12724
rect 19064 12708 19116 12714
rect 19064 12650 19116 12656
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12102 19380 12582
rect 19536 12442 19564 12718
rect 19996 12442 20024 13382
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20088 12646 20116 13262
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20168 12844 20220 12850
rect 20168 12786 20220 12792
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 19524 12436 19576 12442
rect 19524 12378 19576 12384
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 19996 12306 20024 12378
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 18524 11898 18552 12038
rect 19444 11898 19472 12038
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18880 11892 18932 11898
rect 19064 11892 19116 11898
rect 18932 11852 19064 11880
rect 18880 11834 18932 11840
rect 19064 11834 19116 11840
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18524 11286 18552 11630
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18512 11280 18564 11286
rect 18564 11228 18644 11234
rect 18512 11222 18644 11228
rect 18524 11206 18644 11222
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 18236 11144 18288 11150
rect 18236 11086 18288 11092
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18420 11144 18472 11150
rect 18420 11086 18472 11092
rect 18512 11144 18564 11150
rect 18512 11086 18564 11092
rect 17776 10532 17828 10538
rect 17776 10474 17828 10480
rect 17880 10526 18092 10554
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17788 9926 17816 10474
rect 17880 10062 17908 10526
rect 17868 10056 17920 10062
rect 17868 9998 17920 10004
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17224 9580 17276 9586
rect 17224 9522 17276 9528
rect 17696 9518 17724 9862
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17684 9512 17736 9518
rect 17684 9454 17736 9460
rect 17880 9178 17908 9522
rect 18156 9518 18184 11086
rect 18340 10266 18368 11086
rect 18524 10742 18552 11086
rect 18616 10826 18644 11206
rect 18800 11014 18828 11494
rect 18892 11354 18920 11698
rect 18972 11620 19024 11626
rect 18972 11562 19024 11568
rect 18984 11529 19012 11562
rect 18970 11520 19026 11529
rect 18970 11455 19026 11464
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18984 10826 19012 11086
rect 18616 10798 19012 10826
rect 18512 10736 18564 10742
rect 18512 10678 18564 10684
rect 19260 10538 19288 11698
rect 19352 11150 19380 11698
rect 19812 11150 19840 11698
rect 19904 11529 19932 11698
rect 20088 11642 20116 12106
rect 20180 11762 20208 12786
rect 20272 12306 20300 13126
rect 20456 12986 20484 13262
rect 20444 12980 20496 12986
rect 20444 12922 20496 12928
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20456 12238 20484 12582
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20088 11626 20208 11642
rect 20088 11620 20220 11626
rect 20088 11614 20168 11620
rect 20168 11562 20220 11568
rect 20076 11552 20128 11558
rect 19890 11520 19946 11529
rect 20076 11494 20128 11500
rect 19890 11455 19946 11464
rect 19904 11150 19932 11455
rect 20088 11150 20116 11494
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19800 11144 19852 11150
rect 19800 11086 19852 11092
rect 19892 11144 19944 11150
rect 20076 11144 20128 11150
rect 19944 11104 20024 11132
rect 19892 11086 19944 11092
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19248 10532 19300 10538
rect 19248 10474 19300 10480
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 19996 10062 20024 11104
rect 20076 11086 20128 11092
rect 20364 11014 20392 12174
rect 20456 11354 20484 12174
rect 20548 11762 20576 13262
rect 20640 13190 20668 14350
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20640 12306 20668 13126
rect 20732 12434 20760 14470
rect 20824 14278 20852 14758
rect 20904 14544 20956 14550
rect 20902 14512 20904 14521
rect 20956 14512 20958 14521
rect 20902 14447 20958 14456
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20824 13190 20852 14214
rect 21008 13988 21036 15302
rect 21100 15026 21128 15302
rect 21088 15020 21140 15026
rect 21088 14962 21140 14968
rect 21192 14618 21220 16050
rect 21652 16046 21680 16594
rect 21640 16040 21692 16046
rect 21640 15982 21692 15988
rect 22100 15904 22152 15910
rect 22100 15846 22152 15852
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21928 15094 21956 15302
rect 21916 15088 21968 15094
rect 21916 15030 21968 15036
rect 22112 15026 22140 15846
rect 22284 15156 22336 15162
rect 22284 15098 22336 15104
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 22100 15020 22152 15026
rect 22100 14962 22152 14968
rect 21180 14612 21232 14618
rect 21180 14554 21232 14560
rect 21284 14414 21312 14962
rect 22192 14952 22244 14958
rect 22192 14894 22244 14900
rect 22204 14657 22232 14894
rect 22190 14648 22246 14657
rect 22190 14583 22246 14592
rect 22296 14414 22324 15098
rect 22480 15042 22508 18702
rect 22940 17882 22968 19314
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 22928 17876 22980 17882
rect 22928 17818 22980 17824
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22940 17338 22968 17478
rect 22928 17332 22980 17338
rect 22928 17274 22980 17280
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22928 17196 22980 17202
rect 22928 17138 22980 17144
rect 22572 16590 22600 17138
rect 22940 16794 22968 17138
rect 22928 16788 22980 16794
rect 22928 16730 22980 16736
rect 22560 16584 22612 16590
rect 22560 16526 22612 16532
rect 22572 16114 22600 16526
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 23216 15473 23244 18702
rect 23388 18420 23440 18426
rect 23388 18362 23440 18368
rect 23296 17876 23348 17882
rect 23296 17818 23348 17824
rect 23308 17066 23336 17818
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23308 16726 23336 17002
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23308 16114 23336 16662
rect 23400 16250 23428 18362
rect 23492 18358 23520 19450
rect 25608 19310 25636 19790
rect 25596 19304 25648 19310
rect 25596 19246 25648 19252
rect 24584 19236 24636 19242
rect 24584 19178 24636 19184
rect 24492 18760 24544 18766
rect 24492 18702 24544 18708
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23480 18352 23532 18358
rect 23480 18294 23532 18300
rect 23492 17882 23520 18294
rect 23756 18148 23808 18154
rect 23756 18090 23808 18096
rect 23480 17876 23532 17882
rect 23480 17818 23532 17824
rect 23768 17202 23796 18090
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23572 16448 23624 16454
rect 23572 16390 23624 16396
rect 23388 16244 23440 16250
rect 23388 16186 23440 16192
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23388 15496 23440 15502
rect 23202 15464 23258 15473
rect 22744 15428 22796 15434
rect 22744 15370 22796 15376
rect 23124 15422 23202 15450
rect 22388 15014 22508 15042
rect 22560 15020 22612 15026
rect 22388 14822 22416 15014
rect 22560 14962 22612 14968
rect 22376 14816 22428 14822
rect 22376 14758 22428 14764
rect 22468 14816 22520 14822
rect 22572 14804 22600 14962
rect 22520 14776 22600 14804
rect 22468 14758 22520 14764
rect 21272 14408 21324 14414
rect 21272 14350 21324 14356
rect 21824 14408 21876 14414
rect 21824 14350 21876 14356
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 21284 14278 21312 14350
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21192 14074 21220 14214
rect 21284 14074 21312 14214
rect 21836 14074 21864 14350
rect 22376 14272 22428 14278
rect 22480 14260 22508 14758
rect 22756 14550 22784 15370
rect 22836 15020 22888 15026
rect 22836 14962 22888 14968
rect 22744 14544 22796 14550
rect 22744 14486 22796 14492
rect 22848 14278 22876 14962
rect 23124 14822 23152 15422
rect 23388 15438 23440 15444
rect 23202 15399 23258 15408
rect 23204 15360 23256 15366
rect 23204 15302 23256 15308
rect 23216 15094 23244 15302
rect 23204 15088 23256 15094
rect 23204 15030 23256 15036
rect 22928 14816 22980 14822
rect 22928 14758 22980 14764
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23112 14816 23164 14822
rect 23112 14758 23164 14764
rect 22940 14482 22968 14758
rect 22928 14476 22980 14482
rect 22928 14418 22980 14424
rect 22928 14340 22980 14346
rect 23032 14328 23060 14758
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23204 14408 23256 14414
rect 23204 14350 23256 14356
rect 22980 14300 23060 14328
rect 22928 14282 22980 14288
rect 22428 14232 22508 14260
rect 22836 14272 22888 14278
rect 22376 14214 22428 14220
rect 22836 14214 22888 14220
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21824 14068 21876 14074
rect 21824 14010 21876 14016
rect 22388 14006 22416 14214
rect 21088 14000 21140 14006
rect 21008 13960 21088 13988
rect 21088 13942 21140 13948
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 21100 13394 21128 13942
rect 21548 13932 21600 13938
rect 21548 13874 21600 13880
rect 21272 13864 21324 13870
rect 21272 13806 21324 13812
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 20812 13184 20864 13190
rect 20812 13126 20864 13132
rect 20824 12782 20852 13126
rect 20916 12918 20944 13330
rect 21284 13326 21312 13806
rect 21560 13530 21588 13874
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 20904 12912 20956 12918
rect 20904 12854 20956 12860
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20732 12406 20852 12434
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20640 11898 20668 12242
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20444 11348 20496 11354
rect 20444 11290 20496 11296
rect 20352 11008 20404 11014
rect 20352 10950 20404 10956
rect 20364 10062 20392 10950
rect 20456 10130 20484 11290
rect 20824 11150 20852 12406
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21008 11762 21036 11834
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20916 11150 20944 11494
rect 20812 11144 20864 11150
rect 20812 11086 20864 11092
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20916 10810 20944 11086
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21008 10742 21036 11698
rect 21192 11354 21220 11698
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21284 10742 21312 11494
rect 21376 11150 21404 13194
rect 21548 12708 21600 12714
rect 21548 12650 21600 12656
rect 21560 12238 21588 12650
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 21548 12232 21600 12238
rect 21548 12174 21600 12180
rect 21640 12232 21692 12238
rect 21640 12174 21692 12180
rect 21560 11354 21588 12174
rect 21652 11898 21680 12174
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21836 11558 21864 12242
rect 22388 12102 22416 13942
rect 22848 13734 22876 14214
rect 22940 13938 22968 14282
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22836 13728 22888 13734
rect 22836 13670 22888 13676
rect 22848 12434 22876 13670
rect 22940 13326 22968 13874
rect 23124 13530 23152 14350
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23216 13326 23244 14350
rect 23400 14074 23428 15438
rect 23480 15428 23532 15434
rect 23480 15370 23532 15376
rect 23492 14414 23520 15370
rect 23584 15026 23612 16390
rect 23676 16250 23704 17138
rect 23768 16658 23796 17138
rect 23756 16652 23808 16658
rect 23756 16594 23808 16600
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23860 16182 23888 18566
rect 24504 18426 24532 18702
rect 24596 18426 24624 19178
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24688 18766 24716 19110
rect 25700 18834 25728 20318
rect 25780 19848 25832 19854
rect 25976 19836 26004 20402
rect 26056 19984 26108 19990
rect 26056 19926 26108 19932
rect 25832 19808 26004 19836
rect 25780 19790 25832 19796
rect 25976 19514 26004 19808
rect 25964 19508 26016 19514
rect 25964 19450 26016 19456
rect 25780 19168 25832 19174
rect 25780 19110 25832 19116
rect 25792 18970 25820 19110
rect 25780 18964 25832 18970
rect 25780 18906 25832 18912
rect 25688 18828 25740 18834
rect 25688 18770 25740 18776
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 25872 18692 25924 18698
rect 25872 18634 25924 18640
rect 25412 18624 25464 18630
rect 25412 18566 25464 18572
rect 25596 18624 25648 18630
rect 25596 18566 25648 18572
rect 25688 18624 25740 18630
rect 25688 18566 25740 18572
rect 24492 18420 24544 18426
rect 24492 18362 24544 18368
rect 24584 18420 24636 18426
rect 24584 18362 24636 18368
rect 24308 18284 24360 18290
rect 24596 18272 24624 18362
rect 24360 18244 24624 18272
rect 24308 18226 24360 18232
rect 25424 18222 25452 18566
rect 25608 18358 25636 18566
rect 25596 18352 25648 18358
rect 25596 18294 25648 18300
rect 25228 18216 25280 18222
rect 25228 18158 25280 18164
rect 25412 18216 25464 18222
rect 25412 18158 25464 18164
rect 25136 18148 25188 18154
rect 25136 18090 25188 18096
rect 24400 18080 24452 18086
rect 24400 18022 24452 18028
rect 24412 17338 24440 18022
rect 25148 17882 25176 18090
rect 25240 18086 25268 18158
rect 25228 18080 25280 18086
rect 25228 18022 25280 18028
rect 25136 17876 25188 17882
rect 25136 17818 25188 17824
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24032 17332 24084 17338
rect 24032 17274 24084 17280
rect 24400 17332 24452 17338
rect 24400 17274 24452 17280
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 23952 16590 23980 17138
rect 23940 16584 23992 16590
rect 23940 16526 23992 16532
rect 24044 16522 24072 17274
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24136 16590 24164 16934
rect 24412 16590 24440 17274
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24400 16584 24452 16590
rect 24400 16526 24452 16532
rect 24032 16516 24084 16522
rect 24032 16458 24084 16464
rect 23848 16176 23900 16182
rect 23848 16118 23900 16124
rect 23664 15360 23716 15366
rect 23664 15302 23716 15308
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23572 15020 23624 15026
rect 23572 14962 23624 14968
rect 23584 14550 23612 14962
rect 23572 14544 23624 14550
rect 23572 14486 23624 14492
rect 23676 14414 23704 15302
rect 23768 14958 23796 15302
rect 24780 15026 24808 17614
rect 25424 17542 25452 18158
rect 25608 17746 25636 18294
rect 25700 18290 25728 18566
rect 25884 18290 25912 18634
rect 25976 18358 26004 19450
rect 26068 18850 26096 19926
rect 27540 19922 27568 21286
rect 27632 21146 27660 21286
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27632 20398 27660 21082
rect 27620 20392 27672 20398
rect 27620 20334 27672 20340
rect 27528 19916 27580 19922
rect 27528 19858 27580 19864
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 26424 19440 26476 19446
rect 26424 19382 26476 19388
rect 26068 18834 26188 18850
rect 26068 18828 26200 18834
rect 26068 18822 26148 18828
rect 26148 18770 26200 18776
rect 26240 18760 26292 18766
rect 26240 18702 26292 18708
rect 26252 18426 26280 18702
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 25688 18284 25740 18290
rect 25688 18226 25740 18232
rect 25872 18284 25924 18290
rect 25872 18226 25924 18232
rect 26056 18080 26108 18086
rect 26056 18022 26108 18028
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25596 17740 25648 17746
rect 25596 17682 25648 17688
rect 25136 17536 25188 17542
rect 25136 17478 25188 17484
rect 25412 17536 25464 17542
rect 25412 17478 25464 17484
rect 24860 16992 24912 16998
rect 24860 16934 24912 16940
rect 24872 16794 24900 16934
rect 24860 16788 24912 16794
rect 24860 16730 24912 16736
rect 25148 16590 25176 17478
rect 25872 17196 25924 17202
rect 25872 17138 25924 17144
rect 25884 16794 25912 17138
rect 25872 16788 25924 16794
rect 25872 16730 25924 16736
rect 25976 16726 26004 17818
rect 26068 17542 26096 18022
rect 26332 17876 26384 17882
rect 26332 17818 26384 17824
rect 26056 17536 26108 17542
rect 26056 17478 26108 17484
rect 26068 17134 26096 17478
rect 26344 17202 26372 17818
rect 26436 17270 26464 19382
rect 26620 17882 26648 19722
rect 26700 19372 26752 19378
rect 26700 19314 26752 19320
rect 26712 18970 26740 19314
rect 26700 18964 26752 18970
rect 26700 18906 26752 18912
rect 27632 18902 27660 19722
rect 27724 19666 27752 21626
rect 27816 21554 27844 21966
rect 27908 21690 27936 22102
rect 28460 22030 28488 22578
rect 28448 22024 28500 22030
rect 28448 21966 28500 21972
rect 27988 21956 28040 21962
rect 27988 21898 28040 21904
rect 29092 21956 29144 21962
rect 29092 21898 29144 21904
rect 27896 21684 27948 21690
rect 27896 21626 27948 21632
rect 28000 21570 28028 21898
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28828 21622 28856 21830
rect 29104 21690 29132 21898
rect 29092 21684 29144 21690
rect 29092 21626 29144 21632
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27908 21542 28028 21570
rect 28724 21616 28776 21622
rect 28724 21558 28776 21564
rect 28816 21616 28868 21622
rect 28816 21558 28868 21564
rect 28172 21548 28224 21554
rect 27816 19854 27844 21490
rect 27908 20806 27936 21542
rect 28172 21490 28224 21496
rect 27896 20800 27948 20806
rect 27896 20742 27948 20748
rect 27804 19848 27856 19854
rect 27804 19790 27856 19796
rect 27908 19786 27936 20742
rect 28184 20466 28212 21490
rect 28736 21434 28764 21558
rect 29000 21480 29052 21486
rect 28736 21428 29000 21434
rect 28736 21422 29052 21428
rect 28736 21406 29040 21422
rect 28736 20602 28764 21406
rect 28724 20596 28776 20602
rect 28724 20538 28776 20544
rect 28172 20460 28224 20466
rect 28172 20402 28224 20408
rect 28172 20256 28224 20262
rect 28172 20198 28224 20204
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28184 20058 28212 20198
rect 28172 20052 28224 20058
rect 28172 19994 28224 20000
rect 28460 19854 28488 20198
rect 29656 19922 29684 22714
rect 30380 22568 30432 22574
rect 30380 22510 30432 22516
rect 30392 22234 30420 22510
rect 30380 22228 30432 22234
rect 30380 22170 30432 22176
rect 29920 21956 29972 21962
rect 29920 21898 29972 21904
rect 29932 21690 29960 21898
rect 30668 21894 30696 23462
rect 30932 22704 30984 22710
rect 30932 22646 30984 22652
rect 30944 22234 30972 22646
rect 30932 22228 30984 22234
rect 30932 22170 30984 22176
rect 31772 22098 31800 24754
rect 31956 24410 31984 24754
rect 31944 24404 31996 24410
rect 31944 24346 31996 24352
rect 32680 24064 32732 24070
rect 32680 24006 32732 24012
rect 32036 22636 32088 22642
rect 32036 22578 32088 22584
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 31760 22092 31812 22098
rect 31760 22034 31812 22040
rect 32048 22030 32076 22578
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32508 21962 32536 22578
rect 32588 22500 32640 22506
rect 32588 22442 32640 22448
rect 32496 21956 32548 21962
rect 32496 21898 32548 21904
rect 30656 21888 30708 21894
rect 30656 21830 30708 21836
rect 29920 21684 29972 21690
rect 29920 21626 29972 21632
rect 29644 19916 29696 19922
rect 29644 19858 29696 19864
rect 28448 19848 28500 19854
rect 28448 19790 28500 19796
rect 27896 19780 27948 19786
rect 27896 19722 27948 19728
rect 27804 19712 27856 19718
rect 27724 19660 27804 19666
rect 27724 19654 27856 19660
rect 27724 19638 27844 19654
rect 27620 18896 27672 18902
rect 27620 18838 27672 18844
rect 27816 18766 27844 19638
rect 27908 18970 27936 19722
rect 29656 19514 29684 19858
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29656 19334 29684 19450
rect 30668 19378 30696 21830
rect 31852 19916 31904 19922
rect 31852 19858 31904 19864
rect 30748 19780 30800 19786
rect 30748 19722 30800 19728
rect 30760 19514 30788 19722
rect 31864 19514 31892 19858
rect 32128 19848 32180 19854
rect 32128 19790 32180 19796
rect 30748 19508 30800 19514
rect 30748 19450 30800 19456
rect 31852 19508 31904 19514
rect 31852 19450 31904 19456
rect 29564 19306 29684 19334
rect 30656 19372 30708 19378
rect 30656 19314 30708 19320
rect 31668 19372 31720 19378
rect 31668 19314 31720 19320
rect 27896 18964 27948 18970
rect 27896 18906 27948 18912
rect 29564 18766 29592 19306
rect 30196 19168 30248 19174
rect 30196 19110 30248 19116
rect 26792 18760 26844 18766
rect 26792 18702 26844 18708
rect 27804 18760 27856 18766
rect 27804 18702 27856 18708
rect 29552 18760 29604 18766
rect 29552 18702 29604 18708
rect 26608 17876 26660 17882
rect 26608 17818 26660 17824
rect 26516 17740 26568 17746
rect 26516 17682 26568 17688
rect 26424 17264 26476 17270
rect 26424 17206 26476 17212
rect 26332 17196 26384 17202
rect 26332 17138 26384 17144
rect 26056 17128 26108 17134
rect 26056 17070 26108 17076
rect 25964 16720 26016 16726
rect 25964 16662 26016 16668
rect 25976 16590 26004 16662
rect 26068 16658 26096 17070
rect 26240 16788 26292 16794
rect 26240 16730 26292 16736
rect 26056 16652 26108 16658
rect 26056 16594 26108 16600
rect 26252 16590 26280 16730
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 25228 16584 25280 16590
rect 25964 16584 26016 16590
rect 25228 16526 25280 16532
rect 25884 16532 25964 16538
rect 26240 16584 26292 16590
rect 25884 16526 26016 16532
rect 26160 16532 26240 16538
rect 26160 16526 26292 16532
rect 25148 15910 25176 16526
rect 25240 16250 25268 16526
rect 25884 16510 26004 16526
rect 26160 16510 26280 16526
rect 25884 16454 25912 16510
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25872 16448 25924 16454
rect 25872 16390 25924 16396
rect 25964 16448 26016 16454
rect 25964 16390 26016 16396
rect 25228 16244 25280 16250
rect 25228 16186 25280 16192
rect 25424 16114 25452 16390
rect 25884 16114 25912 16390
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 25136 15904 25188 15910
rect 25136 15846 25188 15852
rect 25228 15904 25280 15910
rect 25228 15846 25280 15852
rect 24308 15020 24360 15026
rect 24308 14962 24360 14968
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 23756 14952 23808 14958
rect 23756 14894 23808 14900
rect 24124 14884 24176 14890
rect 24124 14826 24176 14832
rect 23480 14408 23532 14414
rect 23480 14350 23532 14356
rect 23664 14408 23716 14414
rect 23664 14350 23716 14356
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 22928 13320 22980 13326
rect 22928 13262 22980 13268
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23388 13320 23440 13326
rect 23388 13262 23440 13268
rect 23020 13184 23072 13190
rect 23020 13126 23072 13132
rect 22848 12406 22968 12434
rect 22376 12096 22428 12102
rect 22376 12038 22428 12044
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 22282 11384 22338 11393
rect 21548 11348 21600 11354
rect 22282 11319 22338 11328
rect 21548 11290 21600 11296
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21376 10742 21404 11086
rect 22296 11082 22324 11319
rect 22560 11144 22612 11150
rect 22560 11086 22612 11092
rect 22284 11076 22336 11082
rect 22284 11018 22336 11024
rect 21732 11008 21784 11014
rect 21732 10950 21784 10956
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21364 10736 21416 10742
rect 21364 10678 21416 10684
rect 20812 10464 20864 10470
rect 20812 10406 20864 10412
rect 20824 10198 20852 10406
rect 20812 10192 20864 10198
rect 20812 10134 20864 10140
rect 21008 10130 21036 10678
rect 20444 10124 20496 10130
rect 20444 10066 20496 10072
rect 20996 10124 21048 10130
rect 20996 10066 21048 10072
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 18340 9654 18368 9998
rect 18432 9722 18460 9998
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 18420 9716 18472 9722
rect 18420 9658 18472 9664
rect 18328 9648 18380 9654
rect 18328 9590 18380 9596
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18616 9178 18644 9318
rect 16672 9172 16724 9178
rect 16672 9114 16724 9120
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 18604 9172 18656 9178
rect 18604 9114 18656 9120
rect 19444 9110 19472 9522
rect 19996 9178 20024 9998
rect 21008 9654 21036 10066
rect 21284 10062 21312 10678
rect 21744 10130 21772 10950
rect 22296 10674 22324 11018
rect 22572 10674 22600 11086
rect 22940 10742 22968 12406
rect 23032 11626 23060 13126
rect 23400 12850 23428 13262
rect 23676 12986 23704 14350
rect 23768 14074 23796 14350
rect 23756 14068 23808 14074
rect 23756 14010 23808 14016
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23756 13184 23808 13190
rect 23756 13126 23808 13132
rect 23664 12980 23716 12986
rect 23664 12922 23716 12928
rect 23388 12844 23440 12850
rect 23388 12786 23440 12792
rect 23768 12714 23796 13126
rect 23860 12782 23888 13262
rect 24136 12782 24164 14826
rect 24320 14618 24348 14962
rect 24308 14612 24360 14618
rect 24308 14554 24360 14560
rect 24596 14346 24624 14962
rect 24584 14340 24636 14346
rect 24584 14282 24636 14288
rect 25044 13456 25096 13462
rect 25044 13398 25096 13404
rect 24504 13110 24716 13138
rect 24504 12850 24532 13110
rect 24688 12986 24716 13110
rect 25056 12986 25084 13398
rect 24584 12980 24636 12986
rect 24584 12922 24636 12928
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 25044 12980 25096 12986
rect 25044 12922 25096 12928
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24308 12776 24360 12782
rect 24308 12718 24360 12724
rect 23756 12708 23808 12714
rect 23756 12650 23808 12656
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23112 11824 23164 11830
rect 23584 11778 23612 11834
rect 23112 11766 23164 11772
rect 23020 11620 23072 11626
rect 23020 11562 23072 11568
rect 23124 11150 23152 11766
rect 23492 11750 23612 11778
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 22928 10736 22980 10742
rect 22928 10678 22980 10684
rect 23124 10674 23152 11086
rect 23492 10674 23520 11750
rect 23664 11688 23716 11694
rect 23664 11630 23716 11636
rect 23676 11150 23704 11630
rect 23860 11286 23888 12718
rect 24320 12646 24348 12718
rect 24216 12640 24268 12646
rect 24214 12608 24216 12617
rect 24308 12640 24360 12646
rect 24268 12608 24270 12617
rect 24308 12582 24360 12588
rect 24214 12543 24270 12552
rect 24228 11898 24256 12543
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24122 11792 24178 11801
rect 24122 11727 24124 11736
rect 24176 11727 24178 11736
rect 24124 11698 24176 11704
rect 24136 11286 24164 11698
rect 24216 11552 24268 11558
rect 24216 11494 24268 11500
rect 23848 11280 23900 11286
rect 23848 11222 23900 11228
rect 24124 11280 24176 11286
rect 24124 11222 24176 11228
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 24228 11082 24256 11494
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24228 10674 24256 11018
rect 24320 10810 24348 12582
rect 24412 11762 24440 12786
rect 24504 11898 24532 12786
rect 24596 11898 24624 12922
rect 24950 12880 25006 12889
rect 24950 12815 24952 12824
rect 25004 12815 25006 12824
rect 24952 12786 25004 12792
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 24872 12238 24900 12650
rect 25056 12617 25084 12718
rect 25042 12608 25098 12617
rect 25042 12543 25098 12552
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 24860 12232 24912 12238
rect 24860 12174 24912 12180
rect 24492 11892 24544 11898
rect 24492 11834 24544 11840
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24400 11756 24452 11762
rect 24400 11698 24452 11704
rect 24308 10804 24360 10810
rect 24308 10746 24360 10752
rect 24412 10674 24440 11698
rect 25056 11558 25084 12310
rect 25148 11762 25176 15846
rect 25240 15366 25268 15846
rect 25884 15706 25912 16050
rect 25872 15700 25924 15706
rect 25872 15642 25924 15648
rect 25228 15360 25280 15366
rect 25228 15302 25280 15308
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25228 15020 25280 15026
rect 25228 14962 25280 14968
rect 25240 14006 25268 14962
rect 25504 14408 25556 14414
rect 25504 14350 25556 14356
rect 25516 14074 25544 14350
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25228 14000 25280 14006
rect 25228 13942 25280 13948
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25228 13864 25280 13870
rect 25226 13832 25228 13841
rect 25280 13832 25282 13841
rect 25226 13767 25282 13776
rect 25504 13796 25556 13802
rect 25504 13738 25556 13744
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25240 12986 25268 13262
rect 25412 13184 25464 13190
rect 25412 13126 25464 13132
rect 25228 12980 25280 12986
rect 25228 12922 25280 12928
rect 25320 12980 25372 12986
rect 25320 12922 25372 12928
rect 25226 12744 25282 12753
rect 25332 12714 25360 12922
rect 25226 12679 25282 12688
rect 25320 12708 25372 12714
rect 25240 12306 25268 12679
rect 25320 12650 25372 12656
rect 25228 12300 25280 12306
rect 25228 12242 25280 12248
rect 25424 12220 25452 13126
rect 25516 12782 25544 13738
rect 25608 13394 25636 13874
rect 25596 13388 25648 13394
rect 25596 13330 25648 13336
rect 25504 12776 25556 12782
rect 25504 12718 25556 12724
rect 25594 12744 25650 12753
rect 25594 12679 25596 12688
rect 25648 12679 25650 12688
rect 25596 12650 25648 12656
rect 25700 12594 25728 15302
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 25792 13734 25820 13874
rect 25780 13728 25832 13734
rect 25780 13670 25832 13676
rect 25778 12880 25834 12889
rect 25778 12815 25780 12824
rect 25832 12815 25834 12824
rect 25872 12844 25924 12850
rect 25780 12786 25832 12792
rect 25872 12786 25924 12792
rect 25780 12708 25832 12714
rect 25780 12650 25832 12656
rect 25516 12566 25728 12594
rect 25516 12434 25544 12566
rect 25516 12406 25636 12434
rect 25504 12232 25556 12238
rect 25424 12192 25504 12220
rect 25504 12174 25556 12180
rect 25608 11898 25636 12406
rect 25792 12102 25820 12650
rect 25884 12442 25912 12786
rect 25872 12436 25924 12442
rect 25976 12434 26004 16390
rect 26160 16250 26188 16510
rect 26528 16454 26556 17682
rect 26804 17678 26832 18702
rect 30208 18290 30236 19110
rect 31680 18834 31708 19314
rect 31944 19304 31996 19310
rect 31944 19246 31996 19252
rect 31956 18902 31984 19246
rect 32140 19174 32168 19790
rect 32508 19514 32536 21898
rect 32496 19508 32548 19514
rect 32496 19450 32548 19456
rect 32404 19372 32456 19378
rect 32404 19314 32456 19320
rect 32128 19168 32180 19174
rect 32128 19110 32180 19116
rect 31944 18896 31996 18902
rect 31944 18838 31996 18844
rect 31668 18828 31720 18834
rect 31668 18770 31720 18776
rect 32416 18766 32444 19314
rect 32600 18766 32628 22442
rect 32692 22438 32720 24006
rect 32968 22642 32996 24754
rect 33048 24744 33100 24750
rect 33048 24686 33100 24692
rect 33060 24070 33088 24686
rect 34164 24410 34192 24822
rect 34152 24404 34204 24410
rect 34152 24346 34204 24352
rect 34532 24206 34560 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34888 25288 34940 25294
rect 34888 25230 34940 25236
rect 34900 24954 34928 25230
rect 34888 24948 34940 24954
rect 34888 24890 34940 24896
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34520 24200 34572 24206
rect 34520 24142 34572 24148
rect 33048 24064 33100 24070
rect 33048 24006 33100 24012
rect 34060 24064 34112 24070
rect 34060 24006 34112 24012
rect 32956 22636 33008 22642
rect 32956 22578 33008 22584
rect 32680 22432 32732 22438
rect 32680 22374 32732 22380
rect 32692 21894 32720 22374
rect 34072 22030 34100 24006
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34612 23044 34664 23050
rect 34612 22986 34664 22992
rect 34152 22704 34204 22710
rect 34624 22681 34652 22986
rect 34152 22646 34204 22652
rect 34610 22672 34666 22681
rect 34164 22234 34192 22646
rect 34610 22607 34666 22616
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34152 22228 34204 22234
rect 34152 22170 34204 22176
rect 34060 22024 34112 22030
rect 34060 21966 34112 21972
rect 32680 21888 32732 21894
rect 32680 21830 32732 21836
rect 34428 21888 34480 21894
rect 34428 21830 34480 21836
rect 32692 19990 32720 21830
rect 34060 20868 34112 20874
rect 34060 20810 34112 20816
rect 34072 20505 34100 20810
rect 34058 20496 34114 20505
rect 34058 20431 34114 20440
rect 32680 19984 32732 19990
rect 32680 19926 32732 19932
rect 32692 18834 32720 19926
rect 34440 19836 34468 21830
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34520 20936 34572 20942
rect 34520 20878 34572 20884
rect 34532 20058 34560 20878
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34520 20052 34572 20058
rect 34520 19994 34572 20000
rect 34520 19848 34572 19854
rect 34440 19808 34520 19836
rect 34520 19790 34572 19796
rect 34532 19174 34560 19790
rect 34336 19168 34388 19174
rect 34336 19110 34388 19116
rect 34520 19168 34572 19174
rect 34520 19110 34572 19116
rect 32680 18828 32732 18834
rect 32680 18770 32732 18776
rect 33048 18828 33100 18834
rect 33048 18770 33100 18776
rect 32404 18760 32456 18766
rect 32404 18702 32456 18708
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 30288 18692 30340 18698
rect 30288 18634 30340 18640
rect 30300 18426 30328 18634
rect 30288 18420 30340 18426
rect 30288 18362 30340 18368
rect 30196 18284 30248 18290
rect 30196 18226 30248 18232
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26700 17264 26752 17270
rect 26700 17206 26752 17212
rect 26712 17066 26740 17206
rect 26700 17060 26752 17066
rect 26700 17002 26752 17008
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 27252 16992 27304 16998
rect 27252 16934 27304 16940
rect 26240 16448 26292 16454
rect 26240 16390 26292 16396
rect 26516 16448 26568 16454
rect 26516 16390 26568 16396
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 26252 16114 26280 16390
rect 26240 16108 26292 16114
rect 26240 16050 26292 16056
rect 26528 15366 26556 16390
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26332 14952 26384 14958
rect 26332 14894 26384 14900
rect 26240 14884 26292 14890
rect 26240 14826 26292 14832
rect 26252 14074 26280 14826
rect 26344 14074 26372 14894
rect 26528 14550 26556 15302
rect 26804 15026 26832 16934
rect 26976 16040 27028 16046
rect 26976 15982 27028 15988
rect 26988 15570 27016 15982
rect 26976 15564 27028 15570
rect 26976 15506 27028 15512
rect 27160 15428 27212 15434
rect 27160 15370 27212 15376
rect 27172 15162 27200 15370
rect 27160 15156 27212 15162
rect 27160 15098 27212 15104
rect 26792 15020 26844 15026
rect 26792 14962 26844 14968
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26620 14618 26648 14894
rect 26608 14612 26660 14618
rect 26608 14554 26660 14560
rect 26804 14550 26832 14962
rect 27068 14952 27120 14958
rect 27068 14894 27120 14900
rect 26516 14544 26568 14550
rect 26516 14486 26568 14492
rect 26792 14544 26844 14550
rect 26792 14486 26844 14492
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26436 14074 26464 14214
rect 26148 14068 26200 14074
rect 26148 14010 26200 14016
rect 26240 14068 26292 14074
rect 26240 14010 26292 14016
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26160 13954 26188 14010
rect 26056 13932 26108 13938
rect 26160 13926 26372 13954
rect 26056 13874 26108 13880
rect 26068 13784 26096 13874
rect 26240 13796 26292 13802
rect 26068 13756 26240 13784
rect 26068 12782 26096 13756
rect 26240 13738 26292 13744
rect 26344 13530 26372 13926
rect 26332 13524 26384 13530
rect 26332 13466 26384 13472
rect 26424 13184 26476 13190
rect 26424 13126 26476 13132
rect 26436 12850 26464 13126
rect 26148 12844 26200 12850
rect 26148 12786 26200 12792
rect 26424 12844 26476 12850
rect 26424 12786 26476 12792
rect 26056 12776 26108 12782
rect 26056 12718 26108 12724
rect 25976 12406 26096 12434
rect 25872 12378 25924 12384
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25596 11892 25648 11898
rect 25596 11834 25648 11840
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 25608 11354 25636 11834
rect 26068 11694 26096 12406
rect 26160 12238 26188 12786
rect 26436 12617 26464 12786
rect 26422 12608 26478 12617
rect 26422 12543 26478 12552
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26528 11762 26556 14486
rect 27080 14482 27108 14894
rect 27068 14476 27120 14482
rect 27068 14418 27120 14424
rect 27172 12850 27200 15098
rect 27264 15026 27292 16934
rect 30024 16658 30052 18022
rect 30012 16652 30064 16658
rect 30012 16594 30064 16600
rect 29644 16448 29696 16454
rect 29644 16390 29696 16396
rect 29656 16182 29684 16390
rect 29644 16176 29696 16182
rect 29644 16118 29696 16124
rect 29276 15904 29328 15910
rect 29276 15846 29328 15852
rect 29288 15706 29316 15846
rect 29276 15700 29328 15706
rect 29276 15642 29328 15648
rect 27528 15496 27580 15502
rect 27528 15438 27580 15444
rect 27540 15042 27568 15438
rect 29000 15428 29052 15434
rect 29000 15370 29052 15376
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27632 15162 27660 15302
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27540 15026 27844 15042
rect 27252 15020 27304 15026
rect 27540 15020 27856 15026
rect 27540 15014 27804 15020
rect 27252 14962 27304 14968
rect 27528 14952 27580 14958
rect 27528 14894 27580 14900
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 27264 13802 27292 14010
rect 27448 13802 27476 14214
rect 27540 13938 27568 14894
rect 27528 13932 27580 13938
rect 27528 13874 27580 13880
rect 27632 13802 27660 15014
rect 27804 14962 27856 14968
rect 29012 14958 29040 15370
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 28264 14816 28316 14822
rect 28264 14758 28316 14764
rect 28170 14648 28226 14657
rect 28170 14583 28226 14592
rect 28184 14414 28212 14583
rect 28276 14550 28304 14758
rect 29288 14550 29316 15642
rect 30024 15026 30052 16594
rect 32416 16250 32444 18702
rect 32404 16244 32456 16250
rect 32404 16186 32456 16192
rect 31944 16108 31996 16114
rect 31944 16050 31996 16056
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 31116 15904 31168 15910
rect 31116 15846 31168 15852
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 30380 15020 30432 15026
rect 30380 14962 30432 14968
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29920 14816 29972 14822
rect 29920 14758 29972 14764
rect 28264 14544 28316 14550
rect 28264 14486 28316 14492
rect 29276 14544 29328 14550
rect 29276 14486 29328 14492
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 28172 14408 28224 14414
rect 28172 14350 28224 14356
rect 28000 14074 28028 14350
rect 29288 14074 29316 14486
rect 29472 14414 29500 14758
rect 29460 14408 29512 14414
rect 29460 14350 29512 14356
rect 29932 14346 29960 14758
rect 29920 14340 29972 14346
rect 29920 14282 29972 14288
rect 27988 14068 28040 14074
rect 27988 14010 28040 14016
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 27710 13832 27766 13841
rect 27252 13796 27304 13802
rect 27252 13738 27304 13744
rect 27436 13796 27488 13802
rect 27436 13738 27488 13744
rect 27620 13796 27672 13802
rect 27710 13767 27766 13776
rect 27620 13738 27672 13744
rect 27264 13190 27292 13738
rect 27448 13394 27476 13738
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27632 12986 27660 13738
rect 27620 12980 27672 12986
rect 27620 12922 27672 12928
rect 27724 12850 27752 13767
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 28000 12986 28028 13262
rect 29288 12986 29316 14010
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29380 13530 29408 13670
rect 30392 13530 30420 14962
rect 30472 14000 30524 14006
rect 30472 13942 30524 13948
rect 30484 13530 30512 13942
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 30380 13524 30432 13530
rect 30380 13466 30432 13472
rect 30472 13524 30524 13530
rect 30472 13466 30524 13472
rect 27988 12980 28040 12986
rect 27988 12922 28040 12928
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29644 12912 29696 12918
rect 29644 12854 29696 12860
rect 27160 12844 27212 12850
rect 27160 12786 27212 12792
rect 27712 12844 27764 12850
rect 27712 12786 27764 12792
rect 28632 12844 28684 12850
rect 28632 12786 28684 12792
rect 28644 12102 28672 12786
rect 29656 12442 29684 12854
rect 29644 12436 29696 12442
rect 29644 12378 29696 12384
rect 30288 12436 30340 12442
rect 30392 12434 30420 13466
rect 30840 12640 30892 12646
rect 30840 12582 30892 12588
rect 30340 12406 30420 12434
rect 30288 12378 30340 12384
rect 29000 12232 29052 12238
rect 29000 12174 29052 12180
rect 29828 12232 29880 12238
rect 29828 12174 29880 12180
rect 27804 12096 27856 12102
rect 27804 12038 27856 12044
rect 28632 12096 28684 12102
rect 28632 12038 28684 12044
rect 26516 11756 26568 11762
rect 26516 11698 26568 11704
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 26792 11688 26844 11694
rect 26792 11630 26844 11636
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 26068 11286 26096 11630
rect 26148 11552 26200 11558
rect 26148 11494 26200 11500
rect 26160 11354 26188 11494
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 26056 11280 26108 11286
rect 26056 11222 26108 11228
rect 26804 11150 26832 11630
rect 26792 11144 26844 11150
rect 26792 11086 26844 11092
rect 27816 11082 27844 12038
rect 28080 11756 28132 11762
rect 28080 11698 28132 11704
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 28092 11014 28120 11698
rect 28644 11694 28672 12038
rect 29012 11898 29040 12174
rect 29000 11892 29052 11898
rect 29000 11834 29052 11840
rect 28632 11688 28684 11694
rect 28632 11630 28684 11636
rect 29840 11354 29868 12174
rect 30104 11824 30156 11830
rect 30104 11766 30156 11772
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 30116 11354 30144 11766
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30576 11354 30604 11630
rect 30668 11354 30696 11766
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 30564 11348 30616 11354
rect 30564 11290 30616 11296
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30668 11082 30696 11290
rect 30852 11218 30880 12582
rect 31128 12238 31156 15846
rect 31208 15496 31260 15502
rect 31208 15438 31260 15444
rect 31220 15026 31248 15438
rect 31956 15366 31984 16050
rect 32324 15638 32352 16050
rect 32600 15638 32628 18702
rect 33060 18086 33088 18770
rect 34348 18766 34376 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34336 18760 34388 18766
rect 34336 18702 34388 18708
rect 33048 18080 33100 18086
rect 33048 18022 33100 18028
rect 33060 16250 33088 18022
rect 33048 16244 33100 16250
rect 33048 16186 33100 16192
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 32588 15632 32640 15638
rect 32588 15574 32640 15580
rect 31944 15360 31996 15366
rect 31944 15302 31996 15308
rect 31208 15020 31260 15026
rect 31208 14962 31260 14968
rect 31852 15020 31904 15026
rect 31852 14962 31904 14968
rect 31864 14618 31892 14962
rect 31852 14612 31904 14618
rect 31852 14554 31904 14560
rect 31864 14482 31892 14554
rect 31852 14476 31904 14482
rect 31852 14418 31904 14424
rect 31300 14408 31352 14414
rect 31300 14350 31352 14356
rect 31312 13802 31340 14350
rect 31760 14272 31812 14278
rect 31760 14214 31812 14220
rect 31772 14006 31800 14214
rect 31760 14000 31812 14006
rect 31760 13942 31812 13948
rect 31300 13796 31352 13802
rect 31300 13738 31352 13744
rect 31312 13258 31340 13738
rect 31772 13326 31800 13942
rect 31956 13802 31984 15302
rect 32600 15162 32628 15574
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32680 15020 32732 15026
rect 32680 14962 32732 14968
rect 32220 14272 32272 14278
rect 32220 14214 32272 14220
rect 32232 13870 32260 14214
rect 32220 13864 32272 13870
rect 32220 13806 32272 13812
rect 31944 13796 31996 13802
rect 31944 13738 31996 13744
rect 32692 13326 32720 14962
rect 33060 14618 33088 16186
rect 34152 16176 34204 16182
rect 34152 16118 34204 16124
rect 33416 16040 33468 16046
rect 33416 15982 33468 15988
rect 33428 15706 33456 15982
rect 34164 15706 34192 16118
rect 33416 15700 33468 15706
rect 33416 15642 33468 15648
rect 34152 15700 34204 15706
rect 34152 15642 34204 15648
rect 34348 15502 34376 18702
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34532 18426 34560 18566
rect 34520 18420 34572 18426
rect 34520 18362 34572 18368
rect 34794 18320 34850 18329
rect 34794 18255 34796 18264
rect 34848 18255 34850 18264
rect 34796 18226 34848 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34612 16516 34664 16522
rect 34612 16458 34664 16464
rect 34624 16153 34652 16458
rect 34610 16144 34666 16153
rect 34610 16079 34666 16088
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34336 15496 34388 15502
rect 34336 15438 34388 15444
rect 33876 15360 33928 15366
rect 33876 15302 33928 15308
rect 33048 14612 33100 14618
rect 33048 14554 33100 14560
rect 33060 13938 33088 14554
rect 33048 13932 33100 13938
rect 33048 13874 33100 13880
rect 31760 13320 31812 13326
rect 31760 13262 31812 13268
rect 32680 13320 32732 13326
rect 32680 13262 32732 13268
rect 31300 13252 31352 13258
rect 31300 13194 31352 13200
rect 31116 12232 31168 12238
rect 31116 12174 31168 12180
rect 31208 12232 31260 12238
rect 31208 12174 31260 12180
rect 31128 11762 31156 12174
rect 31220 11830 31248 12174
rect 31208 11824 31260 11830
rect 31208 11766 31260 11772
rect 31116 11756 31168 11762
rect 31116 11698 31168 11704
rect 30840 11212 30892 11218
rect 30840 11154 30892 11160
rect 31128 11150 31156 11698
rect 31312 11354 31340 13194
rect 32404 13184 32456 13190
rect 32404 13126 32456 13132
rect 32416 12986 32444 13126
rect 32404 12980 32456 12986
rect 32404 12922 32456 12928
rect 32692 12442 32720 13262
rect 33060 12986 33088 13874
rect 33888 13258 33916 15302
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34612 14340 34664 14346
rect 34612 14282 34664 14288
rect 34060 14000 34112 14006
rect 34624 13977 34652 14282
rect 34060 13942 34112 13948
rect 34610 13968 34666 13977
rect 34072 13530 34100 13942
rect 34610 13903 34666 13912
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34060 13524 34112 13530
rect 34060 13466 34112 13472
rect 33876 13252 33928 13258
rect 33876 13194 33928 13200
rect 34428 13184 34480 13190
rect 34428 13126 34480 13132
rect 34520 13184 34572 13190
rect 34520 13126 34572 13132
rect 33048 12980 33100 12986
rect 33048 12922 33100 12928
rect 33060 12850 33088 12922
rect 34440 12850 34468 13126
rect 33048 12844 33100 12850
rect 33048 12786 33100 12792
rect 34428 12844 34480 12850
rect 34428 12786 34480 12792
rect 31760 12436 31812 12442
rect 31760 12378 31812 12384
rect 32680 12436 32732 12442
rect 32680 12378 32732 12384
rect 31392 12096 31444 12102
rect 31392 12038 31444 12044
rect 31404 11354 31432 12038
rect 31772 11762 31800 12378
rect 33060 11898 33088 12786
rect 34428 12640 34480 12646
rect 34428 12582 34480 12588
rect 34440 12238 34468 12582
rect 34428 12232 34480 12238
rect 34428 12174 34480 12180
rect 33048 11892 33100 11898
rect 33048 11834 33100 11840
rect 34532 11762 34560 13126
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 12164 34664 12170
rect 34612 12106 34664 12112
rect 34624 11801 34652 12106
rect 34610 11792 34666 11801
rect 31760 11756 31812 11762
rect 31760 11698 31812 11704
rect 32496 11756 32548 11762
rect 32496 11698 32548 11704
rect 34520 11756 34572 11762
rect 34610 11727 34666 11736
rect 34520 11698 34572 11704
rect 31668 11620 31720 11626
rect 31668 11562 31720 11568
rect 31300 11348 31352 11354
rect 31300 11290 31352 11296
rect 31392 11348 31444 11354
rect 31392 11290 31444 11296
rect 31680 11150 31708 11562
rect 31116 11144 31168 11150
rect 31116 11086 31168 11092
rect 31668 11144 31720 11150
rect 31668 11086 31720 11092
rect 30656 11076 30708 11082
rect 30656 11018 30708 11024
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 23480 10668 23532 10674
rect 23480 10610 23532 10616
rect 24216 10668 24268 10674
rect 24216 10610 24268 10616
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 22112 10266 22140 10610
rect 22100 10260 22152 10266
rect 22100 10202 22152 10208
rect 21732 10124 21784 10130
rect 21732 10066 21784 10072
rect 22664 10062 22692 10610
rect 23492 10266 23520 10610
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 28092 10062 28120 10950
rect 30668 10674 30696 11018
rect 31128 10810 31156 11086
rect 31772 10810 31800 11698
rect 32508 11286 32536 11698
rect 32772 11688 32824 11694
rect 34532 11665 34560 11698
rect 32772 11630 32824 11636
rect 34518 11656 34574 11665
rect 32784 11354 32812 11630
rect 34518 11591 34574 11600
rect 32864 11552 32916 11558
rect 32864 11494 32916 11500
rect 34244 11552 34296 11558
rect 34244 11494 34296 11500
rect 32876 11354 32904 11494
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 32864 11348 32916 11354
rect 32864 11290 32916 11296
rect 32496 11280 32548 11286
rect 32496 11222 32548 11228
rect 31116 10804 31168 10810
rect 31116 10746 31168 10752
rect 31760 10804 31812 10810
rect 31760 10746 31812 10752
rect 30656 10668 30708 10674
rect 30656 10610 30708 10616
rect 31128 10062 31156 10746
rect 32404 10532 32456 10538
rect 32404 10474 32456 10480
rect 21272 10056 21324 10062
rect 21272 9998 21324 10004
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 27528 10056 27580 10062
rect 27528 9998 27580 10004
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 31116 10056 31168 10062
rect 31116 9998 31168 10004
rect 20996 9648 21048 9654
rect 20996 9590 21048 9596
rect 27540 9586 27568 9998
rect 32312 9920 32364 9926
rect 32312 9862 32364 9868
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 27356 2650 27384 9522
rect 32036 9512 32088 9518
rect 32036 9454 32088 9460
rect 32048 9178 32076 9454
rect 32036 9172 32088 9178
rect 32036 9114 32088 9120
rect 32324 8906 32352 9862
rect 32416 9654 32444 10474
rect 32404 9648 32456 9654
rect 32404 9590 32456 9596
rect 32508 9518 32536 11222
rect 34060 9988 34112 9994
rect 34060 9930 34112 9936
rect 33140 9920 33192 9926
rect 33140 9862 33192 9868
rect 33152 9654 33180 9862
rect 33140 9648 33192 9654
rect 34072 9625 34100 9930
rect 34152 9920 34204 9926
rect 34152 9862 34204 9868
rect 33140 9590 33192 9596
rect 34058 9616 34114 9625
rect 34164 9586 34192 9862
rect 34058 9551 34114 9560
rect 34152 9580 34204 9586
rect 34152 9522 34204 9528
rect 32496 9512 32548 9518
rect 32496 9454 32548 9460
rect 33876 9376 33928 9382
rect 33876 9318 33928 9324
rect 34060 9376 34112 9382
rect 34060 9318 34112 9324
rect 32312 8900 32364 8906
rect 32312 8842 32364 8848
rect 33324 8832 33376 8838
rect 33324 8774 33376 8780
rect 33336 3534 33364 8774
rect 33888 5710 33916 9318
rect 34072 8974 34100 9318
rect 34060 8968 34112 8974
rect 34060 8910 34112 8916
rect 34256 7886 34284 11494
rect 34532 11354 34560 11591
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34520 11348 34572 11354
rect 34520 11290 34572 11296
rect 34428 11212 34480 11218
rect 34428 11154 34480 11160
rect 34440 10062 34468 11154
rect 34532 10810 34560 11290
rect 34520 10804 34572 10810
rect 34520 10746 34572 10752
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34428 10056 34480 10062
rect 34428 9998 34480 10004
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34244 7880 34296 7886
rect 34244 7822 34296 7828
rect 34612 7812 34664 7818
rect 34612 7754 34664 7760
rect 34624 7449 34652 7754
rect 34610 7440 34666 7449
rect 34610 7375 34666 7384
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 33876 5704 33928 5710
rect 33876 5646 33928 5652
rect 34336 5636 34388 5642
rect 34336 5578 34388 5584
rect 34348 5273 34376 5578
rect 34334 5264 34390 5273
rect 34334 5199 34390 5208
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 33324 3528 33376 3534
rect 33324 3470 33376 3476
rect 34888 3460 34940 3466
rect 34888 3402 34940 3408
rect 34900 3097 34928 3402
rect 34886 3088 34942 3097
rect 34886 3023 34942 3032
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 27344 2644 27396 2650
rect 27344 2586 27396 2592
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 27252 2440 27304 2446
rect 27252 2382 27304 2388
rect 952 2009 980 2382
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 9140 1306 9168 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 9048 1278 9168 1306
rect 9048 800 9076 1278
rect 27264 800 27292 2382
rect 9034 0 9090 800
rect 27250 0 27306 800
<< via2 >>
rect 938 36760 994 36816
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 938 34584 994 34640
rect 938 32408 994 32464
rect 1398 30232 1454 30288
rect 938 28056 994 28112
rect 1398 26152 1454 26208
rect 938 23704 994 23760
rect 938 21528 994 21584
rect 938 19352 994 19408
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 938 17196 994 17232
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4986 21564 4988 21584
rect 4988 21564 5040 21584
rect 5040 21564 5042 21584
rect 4986 21528 5042 21564
rect 5814 21564 5816 21584
rect 5816 21564 5868 21584
rect 5868 21564 5870 21584
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 938 17176 940 17196
rect 940 17176 992 17196
rect 992 17176 994 17196
rect 938 15020 994 15056
rect 938 15000 940 15020
rect 940 15000 992 15020
rect 992 15000 994 15020
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 938 12844 994 12880
rect 938 12824 940 12844
rect 940 12824 992 12844
rect 992 12824 994 12844
rect 938 10668 994 10704
rect 938 10648 940 10668
rect 940 10648 992 10668
rect 992 10648 994 10668
rect 938 8472 994 8528
rect 938 6296 994 6352
rect 938 4120 994 4176
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 5814 21528 5870 21564
rect 5446 20712 5502 20768
rect 11334 25900 11390 25936
rect 11334 25880 11336 25900
rect 11336 25880 11388 25900
rect 11388 25880 11390 25900
rect 14094 25900 14150 25936
rect 14094 25880 14096 25900
rect 14096 25880 14148 25900
rect 14148 25880 14150 25900
rect 14462 25764 14518 25800
rect 14462 25744 14464 25764
rect 14464 25744 14516 25764
rect 14516 25744 14518 25764
rect 5262 15136 5318 15192
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 8114 11636 8116 11656
rect 8116 11636 8168 11656
rect 8168 11636 8170 11656
rect 8114 11600 8170 11636
rect 13358 20052 13414 20088
rect 13358 20032 13360 20052
rect 13360 20032 13412 20052
rect 13412 20032 13414 20052
rect 17130 25744 17186 25800
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 21086 26444 21142 26480
rect 21086 26424 21088 26444
rect 21088 26424 21140 26444
rect 21140 26424 21142 26444
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 17958 20052 18014 20088
rect 17958 20032 17960 20052
rect 17960 20032 18012 20052
rect 18012 20032 18014 20052
rect 22926 26444 22982 26480
rect 22926 26424 22928 26444
rect 22928 26424 22980 26444
rect 22980 26424 22982 26444
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20994 23060 20996 23080
rect 20996 23060 21048 23080
rect 21048 23060 21050 23080
rect 20994 23024 21050 23060
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 23202 23024 23258 23080
rect 25134 26988 25190 27024
rect 25134 26968 25136 26988
rect 25136 26968 25188 26988
rect 25188 26968 25190 26988
rect 25686 26868 25688 26888
rect 25688 26868 25740 26888
rect 25740 26868 25742 26888
rect 25686 26832 25742 26868
rect 26330 26988 26386 27024
rect 26330 26968 26332 26988
rect 26332 26968 26384 26988
rect 26384 26968 26386 26988
rect 34334 35672 34390 35728
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34610 33496 34666 33552
rect 34058 31320 34114 31376
rect 26790 26832 26846 26888
rect 34058 29144 34114 29200
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 17406 18284 17462 18320
rect 17406 18264 17408 18284
rect 17408 18264 17460 18284
rect 17460 18264 17462 18284
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19338 18264 19394 18320
rect 34794 26988 34850 27024
rect 34794 26968 34796 26988
rect 34796 26968 34848 26988
rect 34848 26968 34850 26988
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34058 24792 34114 24848
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 17866 15408 17922 15464
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 16854 11756 16910 11792
rect 16854 11736 16856 11756
rect 16856 11736 16908 11756
rect 16908 11736 16910 11756
rect 16302 11328 16358 11384
rect 17590 11192 17646 11248
rect 18142 11192 18198 11248
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 20074 14456 20130 14512
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19338 12960 19394 13016
rect 19522 12824 19578 12880
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 18970 11464 19026 11520
rect 19890 11464 19946 11520
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20902 14492 20904 14512
rect 20904 14492 20956 14512
rect 20956 14492 20958 14512
rect 20902 14456 20958 14492
rect 22190 14592 22246 14648
rect 23202 15408 23258 15464
rect 22282 11328 22338 11384
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 24214 12588 24216 12608
rect 24216 12588 24268 12608
rect 24268 12588 24270 12608
rect 24214 12552 24270 12588
rect 24122 11756 24178 11792
rect 24122 11736 24124 11756
rect 24124 11736 24176 11756
rect 24176 11736 24178 11756
rect 24950 12844 25006 12880
rect 24950 12824 24952 12844
rect 24952 12824 25004 12844
rect 25004 12824 25006 12844
rect 25042 12552 25098 12608
rect 25226 13812 25228 13832
rect 25228 13812 25280 13832
rect 25280 13812 25282 13832
rect 25226 13776 25282 13812
rect 25226 12688 25282 12744
rect 25594 12708 25650 12744
rect 25594 12688 25596 12708
rect 25596 12688 25648 12708
rect 25648 12688 25650 12708
rect 25778 12844 25834 12880
rect 25778 12824 25780 12844
rect 25780 12824 25832 12844
rect 25832 12824 25834 12844
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34610 22616 34666 22672
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34058 20440 34114 20496
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 26422 12552 26478 12608
rect 28170 14592 28226 14648
rect 27710 13776 27766 13832
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34794 18284 34850 18320
rect 34794 18264 34796 18284
rect 34796 18264 34848 18284
rect 34848 18264 34850 18284
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34610 16088 34666 16144
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34610 13912 34666 13968
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34610 11736 34666 11792
rect 34518 11600 34574 11656
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34058 9560 34114 9616
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34610 7384 34666 7440
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34334 5208 34390 5264
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34886 3032 34942 3088
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 938 1944 994 2000
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 34329 35730 34395 35733
rect 35600 35730 36400 35760
rect 34329 35728 36400 35730
rect 34329 35672 34334 35728
rect 34390 35672 36400 35728
rect 34329 35670 36400 35672
rect 34329 35667 34395 35670
rect 35600 35640 36400 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 0 34642 800 34672
rect 933 34642 999 34645
rect 0 34640 999 34642
rect 0 34584 938 34640
rect 994 34584 999 34640
rect 0 34582 999 34584
rect 0 34552 800 34582
rect 933 34579 999 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 34605 33554 34671 33557
rect 35600 33554 36400 33584
rect 34605 33552 36400 33554
rect 34605 33496 34610 33552
rect 34666 33496 36400 33552
rect 34605 33494 36400 33496
rect 34605 33491 34671 33494
rect 35600 33464 36400 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 0 32466 800 32496
rect 933 32466 999 32469
rect 0 32464 999 32466
rect 0 32408 938 32464
rect 994 32408 999 32464
rect 0 32406 999 32408
rect 0 32376 800 32406
rect 933 32403 999 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 34053 31378 34119 31381
rect 35600 31378 36400 31408
rect 34053 31376 36400 31378
rect 34053 31320 34058 31376
rect 34114 31320 36400 31376
rect 34053 31318 36400 31320
rect 34053 31315 34119 31318
rect 35600 31288 36400 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 30290 800 30320
rect 1393 30290 1459 30293
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 800 30230
rect 1393 30227 1459 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 34053 29202 34119 29205
rect 35600 29202 36400 29232
rect 34053 29200 36400 29202
rect 34053 29144 34058 29200
rect 34114 29144 36400 29200
rect 34053 29142 36400 29144
rect 34053 29139 34119 29142
rect 35600 29112 36400 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 0 28114 800 28144
rect 933 28114 999 28117
rect 0 28112 999 28114
rect 0 28056 938 28112
rect 994 28056 999 28112
rect 0 28054 999 28056
rect 0 28024 800 28054
rect 933 28051 999 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 25129 27026 25195 27029
rect 26325 27026 26391 27029
rect 25129 27024 26391 27026
rect 25129 26968 25134 27024
rect 25190 26968 26330 27024
rect 26386 26968 26391 27024
rect 25129 26966 26391 26968
rect 25129 26963 25195 26966
rect 26325 26963 26391 26966
rect 34789 27026 34855 27029
rect 35600 27026 36400 27056
rect 34789 27024 36400 27026
rect 34789 26968 34794 27024
rect 34850 26968 36400 27024
rect 34789 26966 36400 26968
rect 34789 26963 34855 26966
rect 35600 26936 36400 26966
rect 25681 26890 25747 26893
rect 26785 26890 26851 26893
rect 25681 26888 26851 26890
rect 25681 26832 25686 26888
rect 25742 26832 26790 26888
rect 26846 26832 26851 26888
rect 25681 26830 26851 26832
rect 25681 26827 25747 26830
rect 26785 26827 26851 26830
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 21081 26482 21147 26485
rect 22921 26482 22987 26485
rect 21081 26480 22987 26482
rect 21081 26424 21086 26480
rect 21142 26424 22926 26480
rect 22982 26424 22987 26480
rect 21081 26422 22987 26424
rect 21081 26419 21147 26422
rect 22921 26419 22987 26422
rect 1393 26210 1459 26213
rect 798 26208 1459 26210
rect 798 26152 1398 26208
rect 1454 26152 1459 26208
rect 798 26150 1459 26152
rect 798 25968 858 26150
rect 1393 26147 1459 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25878 858 25968
rect 11329 25938 11395 25941
rect 14089 25938 14155 25941
rect 11329 25936 14155 25938
rect 11329 25880 11334 25936
rect 11390 25880 14094 25936
rect 14150 25880 14155 25936
rect 11329 25878 14155 25880
rect 0 25848 800 25878
rect 11329 25875 11395 25878
rect 14089 25875 14155 25878
rect 14457 25802 14523 25805
rect 17125 25802 17191 25805
rect 14457 25800 17191 25802
rect 14457 25744 14462 25800
rect 14518 25744 17130 25800
rect 17186 25744 17191 25800
rect 14457 25742 17191 25744
rect 14457 25739 14523 25742
rect 17125 25739 17191 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 34053 24850 34119 24853
rect 35600 24850 36400 24880
rect 34053 24848 36400 24850
rect 34053 24792 34058 24848
rect 34114 24792 36400 24848
rect 34053 24790 36400 24792
rect 34053 24787 34119 24790
rect 35600 24760 36400 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 20989 23082 21055 23085
rect 23197 23082 23263 23085
rect 20989 23080 23263 23082
rect 20989 23024 20994 23080
rect 21050 23024 23202 23080
rect 23258 23024 23263 23080
rect 20989 23022 23263 23024
rect 20989 23019 21055 23022
rect 23197 23019 23263 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 34605 22674 34671 22677
rect 35600 22674 36400 22704
rect 34605 22672 36400 22674
rect 34605 22616 34610 22672
rect 34666 22616 36400 22672
rect 34605 22614 36400 22616
rect 34605 22611 34671 22614
rect 35600 22584 36400 22614
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 4981 21586 5047 21589
rect 5809 21586 5875 21589
rect 4981 21584 5875 21586
rect 4981 21528 4986 21584
rect 5042 21528 5814 21584
rect 5870 21528 5875 21584
rect 4981 21526 5875 21528
rect 4981 21523 5047 21526
rect 5809 21523 5875 21526
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 5441 20772 5507 20773
rect 5390 20708 5396 20772
rect 5460 20770 5507 20772
rect 5460 20768 5552 20770
rect 5502 20712 5552 20768
rect 5460 20710 5552 20712
rect 5460 20708 5507 20710
rect 5441 20707 5507 20708
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 34053 20498 34119 20501
rect 35600 20498 36400 20528
rect 34053 20496 36400 20498
rect 34053 20440 34058 20496
rect 34114 20440 36400 20496
rect 34053 20438 36400 20440
rect 34053 20435 34119 20438
rect 35600 20408 36400 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 13353 20090 13419 20093
rect 17953 20090 18019 20093
rect 13353 20088 18019 20090
rect 13353 20032 13358 20088
rect 13414 20032 17958 20088
rect 18014 20032 18019 20088
rect 13353 20030 18019 20032
rect 13353 20027 13419 20030
rect 17953 20027 18019 20030
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 17401 18322 17467 18325
rect 19333 18322 19399 18325
rect 17401 18320 19399 18322
rect 17401 18264 17406 18320
rect 17462 18264 19338 18320
rect 19394 18264 19399 18320
rect 17401 18262 19399 18264
rect 17401 18259 17467 18262
rect 19333 18259 19399 18262
rect 34789 18322 34855 18325
rect 35600 18322 36400 18352
rect 34789 18320 36400 18322
rect 34789 18264 34794 18320
rect 34850 18264 36400 18320
rect 34789 18262 36400 18264
rect 34789 18259 34855 18262
rect 35600 18232 36400 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 0 17234 800 17264
rect 933 17234 999 17237
rect 0 17232 999 17234
rect 0 17176 938 17232
rect 994 17176 999 17232
rect 0 17174 999 17176
rect 0 17144 800 17174
rect 933 17171 999 17174
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 34605 16146 34671 16149
rect 35600 16146 36400 16176
rect 34605 16144 36400 16146
rect 34605 16088 34610 16144
rect 34666 16088 36400 16144
rect 34605 16086 36400 16088
rect 34605 16083 34671 16086
rect 35600 16056 36400 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 17861 15466 17927 15469
rect 23197 15466 23263 15469
rect 17861 15464 23263 15466
rect 17861 15408 17866 15464
rect 17922 15408 23202 15464
rect 23258 15408 23263 15464
rect 17861 15406 23263 15408
rect 17861 15403 17927 15406
rect 23197 15403 23263 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 5257 15194 5323 15197
rect 5390 15194 5396 15196
rect 5257 15192 5396 15194
rect 5257 15136 5262 15192
rect 5318 15136 5396 15192
rect 5257 15134 5396 15136
rect 5257 15131 5323 15134
rect 5390 15132 5396 15134
rect 5460 15132 5466 15196
rect 0 15058 800 15088
rect 933 15058 999 15061
rect 0 15056 999 15058
rect 0 15000 938 15056
rect 994 15000 999 15056
rect 0 14998 999 15000
rect 0 14968 800 14998
rect 933 14995 999 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 22185 14650 22251 14653
rect 28165 14650 28231 14653
rect 22185 14648 28231 14650
rect 22185 14592 22190 14648
rect 22246 14592 28170 14648
rect 28226 14592 28231 14648
rect 22185 14590 28231 14592
rect 22185 14587 22251 14590
rect 28165 14587 28231 14590
rect 20069 14514 20135 14517
rect 20897 14514 20963 14517
rect 20069 14512 20963 14514
rect 20069 14456 20074 14512
rect 20130 14456 20902 14512
rect 20958 14456 20963 14512
rect 20069 14454 20963 14456
rect 20069 14451 20135 14454
rect 20897 14451 20963 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 34605 13970 34671 13973
rect 35600 13970 36400 14000
rect 34605 13968 36400 13970
rect 34605 13912 34610 13968
rect 34666 13912 36400 13968
rect 34605 13910 36400 13912
rect 34605 13907 34671 13910
rect 35600 13880 36400 13910
rect 25221 13834 25287 13837
rect 27705 13834 27771 13837
rect 25221 13832 27771 13834
rect 25221 13776 25226 13832
rect 25282 13776 27710 13832
rect 27766 13776 27771 13832
rect 25221 13774 27771 13776
rect 25221 13771 25287 13774
rect 27705 13771 27771 13774
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 19333 13018 19399 13021
rect 19333 13016 19442 13018
rect 19333 12960 19338 13016
rect 19394 12960 19442 13016
rect 19333 12955 19442 12960
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 19382 12882 19442 12955
rect 19517 12882 19583 12885
rect 19382 12880 19583 12882
rect 19382 12824 19522 12880
rect 19578 12824 19583 12880
rect 19382 12822 19583 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 19517 12819 19583 12822
rect 24945 12882 25011 12885
rect 25773 12882 25839 12885
rect 24945 12880 25839 12882
rect 24945 12824 24950 12880
rect 25006 12824 25778 12880
rect 25834 12824 25839 12880
rect 24945 12822 25839 12824
rect 24945 12819 25011 12822
rect 25773 12819 25839 12822
rect 25221 12746 25287 12749
rect 25589 12746 25655 12749
rect 25221 12744 25655 12746
rect 25221 12688 25226 12744
rect 25282 12688 25594 12744
rect 25650 12688 25655 12744
rect 25221 12686 25655 12688
rect 25221 12683 25287 12686
rect 25589 12683 25655 12686
rect 24209 12610 24275 12613
rect 25037 12610 25103 12613
rect 26417 12610 26483 12613
rect 24209 12608 26483 12610
rect 24209 12552 24214 12608
rect 24270 12552 25042 12608
rect 25098 12552 26422 12608
rect 26478 12552 26483 12608
rect 24209 12550 26483 12552
rect 24209 12547 24275 12550
rect 25037 12547 25103 12550
rect 26417 12547 26483 12550
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 16849 11794 16915 11797
rect 24117 11794 24183 11797
rect 16849 11792 24183 11794
rect 16849 11736 16854 11792
rect 16910 11736 24122 11792
rect 24178 11736 24183 11792
rect 16849 11734 24183 11736
rect 16849 11731 16915 11734
rect 24117 11731 24183 11734
rect 34605 11794 34671 11797
rect 35600 11794 36400 11824
rect 34605 11792 36400 11794
rect 34605 11736 34610 11792
rect 34666 11736 36400 11792
rect 34605 11734 36400 11736
rect 34605 11731 34671 11734
rect 35600 11704 36400 11734
rect 8109 11658 8175 11661
rect 34513 11658 34579 11661
rect 8109 11656 34579 11658
rect 8109 11600 8114 11656
rect 8170 11600 34518 11656
rect 34574 11600 34579 11656
rect 8109 11598 34579 11600
rect 8109 11595 8175 11598
rect 34513 11595 34579 11598
rect 18965 11522 19031 11525
rect 19885 11522 19951 11525
rect 18965 11520 19951 11522
rect 18965 11464 18970 11520
rect 19026 11464 19890 11520
rect 19946 11464 19951 11520
rect 18965 11462 19951 11464
rect 18965 11459 19031 11462
rect 19885 11459 19951 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 16297 11386 16363 11389
rect 22277 11386 22343 11389
rect 16297 11384 22343 11386
rect 16297 11328 16302 11384
rect 16358 11328 22282 11384
rect 22338 11328 22343 11384
rect 16297 11326 22343 11328
rect 16297 11323 16363 11326
rect 22277 11323 22343 11326
rect 17585 11250 17651 11253
rect 18137 11250 18203 11253
rect 17585 11248 18203 11250
rect 17585 11192 17590 11248
rect 17646 11192 18142 11248
rect 18198 11192 18203 11248
rect 17585 11190 18203 11192
rect 17585 11187 17651 11190
rect 18137 11187 18203 11190
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 0 10706 800 10736
rect 933 10706 999 10709
rect 0 10704 999 10706
rect 0 10648 938 10704
rect 994 10648 999 10704
rect 0 10646 999 10648
rect 0 10616 800 10646
rect 933 10643 999 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 34053 9618 34119 9621
rect 35600 9618 36400 9648
rect 34053 9616 36400 9618
rect 34053 9560 34058 9616
rect 34114 9560 36400 9616
rect 34053 9558 36400 9560
rect 34053 9555 34119 9558
rect 35600 9528 36400 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 34605 7442 34671 7445
rect 35600 7442 36400 7472
rect 34605 7440 36400 7442
rect 34605 7384 34610 7440
rect 34666 7384 36400 7440
rect 34605 7382 36400 7384
rect 34605 7379 34671 7382
rect 35600 7352 36400 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 34329 5266 34395 5269
rect 35600 5266 36400 5296
rect 34329 5264 36400 5266
rect 34329 5208 34334 5264
rect 34390 5208 36400 5264
rect 34329 5206 36400 5208
rect 34329 5203 34395 5206
rect 35600 5176 36400 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 34881 3090 34947 3093
rect 35600 3090 36400 3120
rect 34881 3088 36400 3090
rect 34881 3032 34886 3088
rect 34942 3032 36400 3088
rect 34881 3030 36400 3032
rect 34881 3027 34947 3030
rect 35600 3000 36400 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
<< via3 >>
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 5396 20768 5460 20772
rect 5396 20712 5446 20768
rect 5446 20712 5460 20768
rect 5396 20708 5460 20712
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 5396 15132 5460 15196
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 36480 4528 36496
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 19568 35936 19888 36496
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 5395 20772 5461 20773
rect 5395 20708 5396 20772
rect 5460 20708 5461 20772
rect 5395 20707 5461 20708
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 5398 15197 5458 20707
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 5395 15196 5461 15197
rect 5395 15132 5396 15196
rect 5460 15132 5461 15196
rect 5395 15131 5461 15132
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 36480 35248 36496
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__and2_1  _0578_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3220 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0579_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0580_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0581_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0582_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0583_
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0584_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0585_
timestamp 1688980957
transform 1 0 5152 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0586_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0587_
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0588_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0589_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0590_
timestamp 1688980957
transform 1 0 4600 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0591_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0592_
timestamp 1688980957
transform 1 0 3220 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0594_
timestamp 1688980957
transform 1 0 4232 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4968 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0596_
timestamp 1688980957
transform 1 0 5060 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0597_
timestamp 1688980957
transform -1 0 5796 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0598_
timestamp 1688980957
transform -1 0 6256 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0599_
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0600_
timestamp 1688980957
transform 1 0 5060 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or4_2  _0601_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0602_
timestamp 1688980957
transform 1 0 5796 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0603_
timestamp 1688980957
transform -1 0 5336 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _0604_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _0605_
timestamp 1688980957
transform -1 0 6716 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0606_
timestamp 1688980957
transform -1 0 5796 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0607_
timestamp 1688980957
transform 1 0 5244 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0608_
timestamp 1688980957
transform 1 0 4968 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0609_
timestamp 1688980957
transform 1 0 4968 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0610_
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0611_
timestamp 1688980957
transform 1 0 5336 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0612_
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0613_
timestamp 1688980957
transform 1 0 4508 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0614_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _0615_
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0616_
timestamp 1688980957
transform 1 0 5428 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _0617_
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0618_
timestamp 1688980957
transform -1 0 6992 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0619_
timestamp 1688980957
transform -1 0 8464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0620_
timestamp 1688980957
transform 1 0 30728 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _0621_
timestamp 1688980957
transform 1 0 31464 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0622_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0623_
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0624_
timestamp 1688980957
transform -1 0 32292 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0625_
timestamp 1688980957
transform -1 0 32016 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _0626_
timestamp 1688980957
transform 1 0 31372 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0627_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__o31a_1  _0628_
timestamp 1688980957
transform 1 0 31372 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0629_
timestamp 1688980957
transform 1 0 30728 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0630_
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0631_
timestamp 1688980957
transform 1 0 32016 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0632_
timestamp 1688980957
transform 1 0 32660 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0633_
timestamp 1688980957
transform 1 0 31924 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0634_
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0635_
timestamp 1688980957
transform 1 0 31832 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0636_
timestamp 1688980957
transform 1 0 31832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0637_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0638_
timestamp 1688980957
transform 1 0 32752 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0639_
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0640_
timestamp 1688980957
transform 1 0 32752 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0641_
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0642_
timestamp 1688980957
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0643_
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0644_
timestamp 1688980957
transform 1 0 32384 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0645_
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0646_
timestamp 1688980957
transform 1 0 32384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0647_
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0648_
timestamp 1688980957
transform 1 0 31556 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0649_
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0650_
timestamp 1688980957
transform 1 0 32476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0651_
timestamp 1688980957
transform 1 0 31832 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _0652_
timestamp 1688980957
transform 1 0 31280 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _0653_
timestamp 1688980957
transform 1 0 30636 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _0654_
timestamp 1688980957
transform 1 0 31096 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0655_
timestamp 1688980957
transform 1 0 31372 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0656_
timestamp 1688980957
transform -1 0 31556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0657_
timestamp 1688980957
transform 1 0 30636 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _0658_
timestamp 1688980957
transform -1 0 31556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _0659_
timestamp 1688980957
transform -1 0 32292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0660_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  _0661_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  _0662_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _0663_
timestamp 1688980957
transform 1 0 22816 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0664_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  _0665_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_8  _0666_
timestamp 1688980957
transform 1 0 9016 0 1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  _0667_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0668_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22632 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0669_
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _0670_
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0671_
timestamp 1688980957
transform 1 0 21712 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0672_
timestamp 1688980957
transform 1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0673_
timestamp 1688980957
transform -1 0 23000 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0674_
timestamp 1688980957
transform -1 0 22816 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _0675_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0676_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22724 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0677_
timestamp 1688980957
transform -1 0 24288 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0678_
timestamp 1688980957
transform 1 0 23000 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0679_
timestamp 1688980957
transform -1 0 24196 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0680_
timestamp 1688980957
transform 1 0 23276 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _0681_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26036 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0682_
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0683_
timestamp 1688980957
transform -1 0 22816 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0684_
timestamp 1688980957
transform -1 0 23092 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0685_
timestamp 1688980957
transform 1 0 21896 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _0686_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23552 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0687_
timestamp 1688980957
transform -1 0 23736 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _0688_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0689_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _0690_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0691_
timestamp 1688980957
transform -1 0 24288 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0692_
timestamp 1688980957
transform 1 0 23184 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0693_
timestamp 1688980957
transform 1 0 23276 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0694_
timestamp 1688980957
transform 1 0 24380 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0695_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24748 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_1  _0696_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24288 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0697_
timestamp 1688980957
transform -1 0 24196 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _0698_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23920 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _0699_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23276 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _0700_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0701_
timestamp 1688980957
transform 1 0 22080 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0702_
timestamp 1688980957
transform -1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0703_
timestamp 1688980957
transform 1 0 22080 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0704_
timestamp 1688980957
transform 1 0 24932 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0705_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0706_
timestamp 1688980957
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0707_
timestamp 1688980957
transform -1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0708_
timestamp 1688980957
transform -1 0 24932 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0709_
timestamp 1688980957
transform -1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0710_
timestamp 1688980957
transform 1 0 25484 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0711_
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  _0712_
timestamp 1688980957
transform 1 0 8096 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0713_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _0714_
timestamp 1688980957
transform 1 0 9292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  _0715_
timestamp 1688980957
transform 1 0 8188 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0716_
timestamp 1688980957
transform 1 0 17204 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0717_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_6  _0718_
timestamp 1688980957
transform 1 0 10304 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0719_
timestamp 1688980957
transform 1 0 14168 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _0720_
timestamp 1688980957
transform 1 0 10580 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0721_
timestamp 1688980957
transform 1 0 14444 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0722_
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_8  _0723_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_2  _0724_
timestamp 1688980957
transform 1 0 12512 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _0725_
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_2  _0726_
timestamp 1688980957
transform -1 0 13156 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0727_
timestamp 1688980957
transform 1 0 11960 0 1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_2  _0728_
timestamp 1688980957
transform -1 0 19688 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _0729_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0730_
timestamp 1688980957
transform -1 0 17112 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0731_
timestamp 1688980957
transform -1 0 17756 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0732_
timestamp 1688980957
transform 1 0 16744 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0733_
timestamp 1688980957
transform 1 0 16652 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0734_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0735_
timestamp 1688980957
transform -1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _0736_
timestamp 1688980957
transform 1 0 17572 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0737_
timestamp 1688980957
transform -1 0 16376 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _0738_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _0739_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and4_1  _0740_
timestamp 1688980957
transform 1 0 16100 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0741_
timestamp 1688980957
transform -1 0 17480 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0742_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2ai_1  _0743_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _0744_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18124 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _0745_
timestamp 1688980957
transform 1 0 17572 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0746_
timestamp 1688980957
transform -1 0 21620 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _0747_
timestamp 1688980957
transform 1 0 21252 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _0748_
timestamp 1688980957
transform 1 0 20148 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0749_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0750_
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0751_
timestamp 1688980957
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _0752_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20056 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0753_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_4  _0754_
timestamp 1688980957
transform 1 0 18768 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_2  _0755_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21712 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0756_
timestamp 1688980957
transform -1 0 14536 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _0757_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_2  _0758_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16468 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0759_
timestamp 1688980957
transform -1 0 19136 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_4  _0760_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__a21o_1  _0761_
timestamp 1688980957
transform 1 0 18216 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0762_
timestamp 1688980957
transform -1 0 17572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o41ai_1  _0763_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18032 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _0764_
timestamp 1688980957
transform 1 0 16928 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _0765_
timestamp 1688980957
transform 1 0 16744 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a32oi_4  _0766_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24288 0 1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_1  _0767_
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1688980957
transform 1 0 21620 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _0769_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22356 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _0770_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23368 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _0771_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23460 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _0772_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25300 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _0773_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25392 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _0774_
timestamp 1688980957
transform -1 0 26772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _0775_
timestamp 1688980957
transform 1 0 23828 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _0776_
timestamp 1688980957
transform -1 0 24932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0777_
timestamp 1688980957
transform -1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0778_
timestamp 1688980957
transform 1 0 25392 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0779_
timestamp 1688980957
transform 1 0 24288 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _0780_
timestamp 1688980957
transform 1 0 24840 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0781_
timestamp 1688980957
transform 1 0 26128 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1688980957
transform -1 0 26220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0783_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26128 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _0784_
timestamp 1688980957
transform -1 0 27508 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0785_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0786_
timestamp 1688980957
transform 1 0 25392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0787_
timestamp 1688980957
transform -1 0 26496 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0788_
timestamp 1688980957
transform 1 0 25668 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _0789_
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0790_
timestamp 1688980957
transform 1 0 26864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _0791_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27692 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0792_
timestamp 1688980957
transform 1 0 27692 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0793_
timestamp 1688980957
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _0794_
timestamp 1688980957
transform 1 0 25852 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _0795_
timestamp 1688980957
transform -1 0 24932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0796_
timestamp 1688980957
transform -1 0 24564 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2111oi_1  _0797_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25392 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0798_
timestamp 1688980957
transform 1 0 26956 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _0799_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0800_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _0801_
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0802_
timestamp 1688980957
transform -1 0 18032 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0803_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _0804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18032 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0805_
timestamp 1688980957
transform -1 0 18676 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _0806_
timestamp 1688980957
transform -1 0 21344 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a22oi_2  _0807_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21252 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__o221a_1  _0808_
timestamp 1688980957
transform 1 0 18676 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand4b_2  _0809_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23276 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0810_
timestamp 1688980957
transform 1 0 17664 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0811_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23552 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _0812_
timestamp 1688980957
transform 1 0 22724 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0813_
timestamp 1688980957
transform -1 0 22632 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0814_
timestamp 1688980957
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0815_
timestamp 1688980957
transform -1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0816_
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0817_
timestamp 1688980957
transform -1 0 24840 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0818_
timestamp 1688980957
transform 1 0 23460 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _0819_
timestamp 1688980957
transform -1 0 24196 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0820_
timestamp 1688980957
transform -1 0 23000 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0821_
timestamp 1688980957
transform 1 0 21252 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0822_
timestamp 1688980957
transform 1 0 13892 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0823_
timestamp 1688980957
transform 1 0 11868 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a311o_1  _0824_
timestamp 1688980957
transform -1 0 14812 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2b_1  _0825_
timestamp 1688980957
transform -1 0 13248 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0826_
timestamp 1688980957
transform -1 0 12696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0827_
timestamp 1688980957
transform -1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0829_
timestamp 1688980957
transform -1 0 13984 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0830_
timestamp 1688980957
transform -1 0 14536 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _0831_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_2  _0832_
timestamp 1688980957
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 1688980957
transform -1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1688980957
transform -1 0 18768 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0835_
timestamp 1688980957
transform 1 0 20056 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _0836_
timestamp 1688980957
transform -1 0 18400 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2b_1  _0837_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _0838_
timestamp 1688980957
transform -1 0 13248 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _0839_
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _0840_
timestamp 1688980957
transform 1 0 11684 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _0841_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _0842_
timestamp 1688980957
transform 1 0 20516 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0843_
timestamp 1688980957
transform 1 0 21896 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0844_
timestamp 1688980957
transform -1 0 24012 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _0845_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22632 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _0846_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0847_
timestamp 1688980957
transform -1 0 23000 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _0848_
timestamp 1688980957
transform 1 0 22632 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_2  _0849_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24932 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0850_
timestamp 1688980957
transform -1 0 9660 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0851_
timestamp 1688980957
transform 1 0 9844 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _0852_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand4b_2  _0853_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _0854_
timestamp 1688980957
transform -1 0 12236 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _0855_
timestamp 1688980957
transform 1 0 11224 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _0856_
timestamp 1688980957
transform -1 0 12972 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _0857_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13892 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0858_
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _0859_
timestamp 1688980957
transform -1 0 8924 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _0860_
timestamp 1688980957
transform 1 0 9200 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _0861_
timestamp 1688980957
transform 1 0 8924 0 -1 25024
box -38 -48 2062 592
use sky130_fd_sc_hd__o311ai_4  _0862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__a211oi_1  _0863_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11224 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a2111o_1  _0864_
timestamp 1688980957
transform 1 0 10396 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _0865_
timestamp 1688980957
transform 1 0 13064 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _0866_
timestamp 1688980957
transform -1 0 15180 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _0867_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _0868_
timestamp 1688980957
transform 1 0 14904 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0869_
timestamp 1688980957
transform -1 0 17112 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0870_
timestamp 1688980957
transform 1 0 15364 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _0871_
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0872_
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _0873_
timestamp 1688980957
transform 1 0 14628 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0874_
timestamp 1688980957
transform 1 0 17940 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _0875_
timestamp 1688980957
transform 1 0 18768 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0876_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _0877_
timestamp 1688980957
transform 1 0 11316 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _0878_
timestamp 1688980957
transform 1 0 10948 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _0879_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _0880_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _0881_
timestamp 1688980957
transform 1 0 19228 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _0882_
timestamp 1688980957
transform -1 0 21344 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _0883_
timestamp 1688980957
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0884_
timestamp 1688980957
transform 1 0 20516 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0885_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0886_
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _0887_
timestamp 1688980957
transform -1 0 22632 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0888_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _0889_
timestamp 1688980957
transform 1 0 21896 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _0890_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _0891_
timestamp 1688980957
transform 1 0 20424 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a32oi_4  _0892_
timestamp 1688980957
transform -1 0 22356 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _0893_
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ba_1  _0894_
timestamp 1688980957
transform 1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0895_
timestamp 1688980957
transform 1 0 16560 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _0896_
timestamp 1688980957
transform 1 0 11224 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_2  _0897_
timestamp 1688980957
transform -1 0 14168 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _0898_
timestamp 1688980957
transform -1 0 13800 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o2111ai_4  _0899_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15272 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__a311o_1  _0900_
timestamp 1688980957
transform -1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0901_
timestamp 1688980957
transform 1 0 16008 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _0902_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17572 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a211o_1  _0903_
timestamp 1688980957
transform 1 0 15364 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _0904_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0905_
timestamp 1688980957
transform -1 0 15732 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0906_
timestamp 1688980957
transform -1 0 16560 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0907_
timestamp 1688980957
transform -1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0908_
timestamp 1688980957
transform -1 0 16008 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0909_
timestamp 1688980957
transform -1 0 16284 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0910_
timestamp 1688980957
transform -1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0911_
timestamp 1688980957
transform -1 0 17664 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _0912_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17664 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _0913_
timestamp 1688980957
transform -1 0 20240 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0914_
timestamp 1688980957
transform -1 0 15548 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0915_
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _0916_
timestamp 1688980957
transform 1 0 9568 0 1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_2  _0917_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0918_
timestamp 1688980957
transform -1 0 13800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0919_
timestamp 1688980957
transform -1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _0920_
timestamp 1688980957
transform 1 0 13156 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0921_
timestamp 1688980957
transform 1 0 10856 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0922_
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _0923_
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _0924_
timestamp 1688980957
transform 1 0 11316 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _0925_
timestamp 1688980957
transform 1 0 10672 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _0926_
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _0927_
timestamp 1688980957
transform 1 0 12052 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0928_
timestamp 1688980957
transform 1 0 12880 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _0929_
timestamp 1688980957
transform 1 0 11500 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_1  _0930_
timestamp 1688980957
transform -1 0 10856 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _0931_
timestamp 1688980957
transform -1 0 11500 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0932_
timestamp 1688980957
transform 1 0 15732 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0933_
timestamp 1688980957
transform 1 0 19136 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _0934_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20424 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__or3_1  _0935_
timestamp 1688980957
transform 1 0 20608 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _0936_
timestamp 1688980957
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _0937_
timestamp 1688980957
transform 1 0 26312 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0938_
timestamp 1688980957
transform 1 0 25668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0939_
timestamp 1688980957
transform 1 0 25392 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _0940_
timestamp 1688980957
transform 1 0 25944 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_2  _0941_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23092 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_1  _0942_
timestamp 1688980957
transform 1 0 27140 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0943_
timestamp 1688980957
transform -1 0 28428 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _0944_
timestamp 1688980957
transform 1 0 27600 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_2  _0945_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20608 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__o311a_1  _0946_
timestamp 1688980957
transform -1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _0947_
timestamp 1688980957
transform -1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0948_
timestamp 1688980957
transform -1 0 12972 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _0949_
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _0950_
timestamp 1688980957
transform 1 0 15088 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_1  _0951_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15732 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _0952_
timestamp 1688980957
transform 1 0 17664 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0953_
timestamp 1688980957
transform 1 0 17112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _0954_
timestamp 1688980957
transform -1 0 18584 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1688980957
transform 1 0 16468 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _0956_
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1688980957
transform -1 0 13064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0958_
timestamp 1688980957
transform -1 0 13340 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _0959_
timestamp 1688980957
transform -1 0 12052 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _0960_
timestamp 1688980957
transform -1 0 12788 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _0961_
timestamp 1688980957
transform 1 0 13156 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _0962_
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _0963_
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0964_
timestamp 1688980957
transform 1 0 17020 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _0965_
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _0966_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18400 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _0967_
timestamp 1688980957
transform -1 0 17296 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0968_
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _0969_
timestamp 1688980957
transform 1 0 17296 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0970_
timestamp 1688980957
transform -1 0 15732 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0971_
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _0972_
timestamp 1688980957
transform 1 0 15088 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0973_
timestamp 1688980957
transform -1 0 13340 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0974_
timestamp 1688980957
transform 1 0 12788 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0975_
timestamp 1688980957
transform -1 0 14628 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0976_
timestamp 1688980957
transform -1 0 13892 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1688980957
transform -1 0 12972 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _0978_
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _0979_
timestamp 1688980957
transform 1 0 13524 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1688980957
transform -1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _0981_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14812 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _0982_
timestamp 1688980957
transform -1 0 15364 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _0983_
timestamp 1688980957
transform 1 0 12972 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _0984_
timestamp 1688980957
transform -1 0 14076 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _0985_
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0986_
timestamp 1688980957
transform 1 0 17480 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _0987_
timestamp 1688980957
transform 1 0 18400 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _0988_
timestamp 1688980957
transform 1 0 19412 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_1  _0989_
timestamp 1688980957
transform 1 0 27508 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _0990_
timestamp 1688980957
transform -1 0 26312 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _0991_
timestamp 1688980957
transform -1 0 26864 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _0992_
timestamp 1688980957
transform -1 0 27600 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2111o_2  _0993_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25852 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _0994_
timestamp 1688980957
transform -1 0 22448 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _0995_
timestamp 1688980957
transform -1 0 20516 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _0996_
timestamp 1688980957
transform 1 0 20516 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0997_
timestamp 1688980957
transform -1 0 20976 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _0998_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _0999_
timestamp 1688980957
transform -1 0 22080 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _1000_
timestamp 1688980957
transform -1 0 22448 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1688980957
transform -1 0 27692 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1002_
timestamp 1688980957
transform 1 0 27232 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1003_
timestamp 1688980957
transform 1 0 25484 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1004_
timestamp 1688980957
transform 1 0 18676 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1005_
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _1006_
timestamp 1688980957
transform -1 0 19872 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1007_
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a41o_1  _1008_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _1009_
timestamp 1688980957
transform -1 0 18032 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1010_
timestamp 1688980957
transform 1 0 17204 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1011_
timestamp 1688980957
transform -1 0 17848 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_2  _1012_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18584 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1013_
timestamp 1688980957
transform -1 0 16376 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1014_
timestamp 1688980957
transform -1 0 15640 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1015_
timestamp 1688980957
transform -1 0 15088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1016_
timestamp 1688980957
transform 1 0 15272 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1017_
timestamp 1688980957
transform 1 0 15272 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1018_
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1019_
timestamp 1688980957
transform 1 0 12972 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1020_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1021_
timestamp 1688980957
transform 1 0 15640 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a31oi_1  _1022_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1023_
timestamp 1688980957
transform 1 0 15732 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_2  _1024_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14904 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1025_
timestamp 1688980957
transform 1 0 18952 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1026_
timestamp 1688980957
transform 1 0 19596 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ba_1  _1027_
timestamp 1688980957
transform -1 0 26312 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1028_
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1029_
timestamp 1688980957
transform -1 0 27416 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1030_
timestamp 1688980957
transform -1 0 19872 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1031_
timestamp 1688980957
transform 1 0 16744 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1032_
timestamp 1688980957
transform -1 0 16744 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1033_
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1034_
timestamp 1688980957
transform 1 0 16560 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1035_
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1036_
timestamp 1688980957
transform -1 0 16008 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _1037_
timestamp 1688980957
transform -1 0 16744 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1038_
timestamp 1688980957
transform 1 0 17112 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__a211oi_1  _1039_
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1040_
timestamp 1688980957
transform -1 0 19136 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_1  _1041_
timestamp 1688980957
transform 1 0 18032 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _1042_
timestamp 1688980957
transform -1 0 20056 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nor3b_1  _1043_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27324 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _1044_
timestamp 1688980957
transform -1 0 27232 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1045_
timestamp 1688980957
transform 1 0 27876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1046_
timestamp 1688980957
transform 1 0 29072 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1047_
timestamp 1688980957
transform 1 0 28152 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1048_
timestamp 1688980957
transform -1 0 27600 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1049_
timestamp 1688980957
transform -1 0 27232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _1050_
timestamp 1688980957
transform -1 0 26128 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1688980957
transform -1 0 24656 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1052_
timestamp 1688980957
transform 1 0 24656 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1053_
timestamp 1688980957
transform 1 0 24840 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _1054_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21620 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1055_
timestamp 1688980957
transform 1 0 17388 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1056_
timestamp 1688980957
transform -1 0 17940 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1057_
timestamp 1688980957
transform -1 0 19504 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1058_
timestamp 1688980957
transform -1 0 19872 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1059_
timestamp 1688980957
transform -1 0 20240 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1060_
timestamp 1688980957
transform -1 0 20516 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_4  _1061_
timestamp 1688980957
transform 1 0 20516 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1062_
timestamp 1688980957
transform 1 0 27508 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1063_
timestamp 1688980957
transform -1 0 24656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1064_
timestamp 1688980957
transform 1 0 23552 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1065_
timestamp 1688980957
transform -1 0 23552 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1066_
timestamp 1688980957
transform 1 0 23552 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1067_
timestamp 1688980957
transform -1 0 28060 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1068_
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _1069_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1688980957
transform 1 0 28336 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1071_
timestamp 1688980957
transform 1 0 25300 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1072_
timestamp 1688980957
transform 1 0 25668 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _1073_
timestamp 1688980957
transform 1 0 25760 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _1074_
timestamp 1688980957
transform 1 0 22080 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__a211o_1  _1075_
timestamp 1688980957
transform -1 0 26312 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1076_
timestamp 1688980957
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1077_
timestamp 1688980957
transform 1 0 26312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1078_
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1079_
timestamp 1688980957
transform 1 0 24196 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4bb_1  _1080_
timestamp 1688980957
transform 1 0 24656 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__o31ai_1  _1081_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26128 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1082_
timestamp 1688980957
transform -1 0 27692 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1083_
timestamp 1688980957
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 1688980957
transform 1 0 24932 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1085_
timestamp 1688980957
transform 1 0 24840 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1086_
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1087_
timestamp 1688980957
transform 1 0 27784 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1088_
timestamp 1688980957
transform 1 0 28520 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1089_
timestamp 1688980957
transform 1 0 27600 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1090_
timestamp 1688980957
transform 1 0 28520 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1091_
timestamp 1688980957
transform 1 0 28796 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1092_
timestamp 1688980957
transform 1 0 28336 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1093_
timestamp 1688980957
transform -1 0 29624 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1094_
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1095_
timestamp 1688980957
transform -1 0 27968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1096_
timestamp 1688980957
transform 1 0 28428 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1097_
timestamp 1688980957
transform 1 0 28244 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1098_
timestamp 1688980957
transform -1 0 29532 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1099_
timestamp 1688980957
transform 1 0 28704 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1100_
timestamp 1688980957
transform 1 0 29716 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1101_
timestamp 1688980957
transform -1 0 30452 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1102_
timestamp 1688980957
transform -1 0 27968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1103_
timestamp 1688980957
transform -1 0 28428 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1104_
timestamp 1688980957
transform 1 0 27784 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1105_
timestamp 1688980957
transform 1 0 27692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1106_
timestamp 1688980957
transform 1 0 28612 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1688980957
transform -1 0 21620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1108_
timestamp 1688980957
transform 1 0 20792 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1109_
timestamp 1688980957
transform 1 0 19320 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1110_
timestamp 1688980957
transform 1 0 20240 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _1111_
timestamp 1688980957
transform -1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1112_
timestamp 1688980957
transform 1 0 21712 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1113_
timestamp 1688980957
transform -1 0 26496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1114_
timestamp 1688980957
transform 1 0 25300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1115_
timestamp 1688980957
transform 1 0 25576 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1116_
timestamp 1688980957
transform -1 0 20516 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1117_
timestamp 1688980957
transform -1 0 21620 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1118_
timestamp 1688980957
transform 1 0 20792 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1119_
timestamp 1688980957
transform 1 0 19228 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1120_
timestamp 1688980957
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1121_
timestamp 1688980957
transform 1 0 20516 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1122_
timestamp 1688980957
transform 1 0 20148 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1123_
timestamp 1688980957
transform -1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1124_
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1125_
timestamp 1688980957
transform -1 0 23828 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1126_
timestamp 1688980957
transform 1 0 23644 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1127_
timestamp 1688980957
transform 1 0 24932 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1688980957
transform 1 0 26404 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1129_
timestamp 1688980957
transform -1 0 27508 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1130_
timestamp 1688980957
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1131_
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1132_
timestamp 1688980957
transform 1 0 27784 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_8  _1133_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  _1134_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1135_
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1688980957
transform -1 0 9936 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1137_
timestamp 1688980957
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1138_
timestamp 1688980957
transform 1 0 30176 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1139_
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1688980957
transform 1 0 31464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1141_
timestamp 1688980957
transform 1 0 30452 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1688980957
transform 1 0 30728 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1143_
timestamp 1688980957
transform 1 0 30820 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1688980957
transform 1 0 30636 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1145_
timestamp 1688980957
transform 1 0 30176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1146_
timestamp 1688980957
transform 1 0 31372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1147_
timestamp 1688980957
transform 1 0 30452 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1688980957
transform 1 0 29808 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1149_
timestamp 1688980957
transform -1 0 30268 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1150_
timestamp 1688980957
transform 1 0 29624 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1688980957
transform 1 0 27784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1152_
timestamp 1688980957
transform -1 0 29808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1153_
timestamp 1688980957
transform -1 0 10304 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1154_
timestamp 1688980957
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1155_
timestamp 1688980957
transform -1 0 8648 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1688980957
transform -1 0 10304 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1157_
timestamp 1688980957
transform -1 0 8648 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1158_
timestamp 1688980957
transform 1 0 7544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1159_
timestamp 1688980957
transform 1 0 9844 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1160_
timestamp 1688980957
transform 1 0 7360 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1161_
timestamp 1688980957
transform -1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1688980957
transform -1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1163_
timestamp 1688980957
transform -1 0 8648 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1164_
timestamp 1688980957
transform 1 0 8004 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1165_
timestamp 1688980957
transform -1 0 8464 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1688980957
transform -1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1167_
timestamp 1688980957
transform 1 0 7728 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1168_
timestamp 1688980957
transform -1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1169_
timestamp 1688980957
transform -1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1170_
timestamp 1688980957
transform 1 0 8004 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1171_
timestamp 1688980957
transform -1 0 10580 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1172_
timestamp 1688980957
transform -1 0 34224 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1173_
timestamp 1688980957
transform 1 0 32660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _1174_
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _1175_
timestamp 1688980957
transform -1 0 34592 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1176_
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1177_
timestamp 1688980957
transform -1 0 34592 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1178_
timestamp 1688980957
transform 1 0 34040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1179_
timestamp 1688980957
transform 1 0 34040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1180_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1181_
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1182_
timestamp 1688980957
transform 1 0 34132 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1183_
timestamp 1688980957
transform 1 0 34132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1185_
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1186_
timestamp 1688980957
transform -1 0 34408 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1187_
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1189_
timestamp 1688980957
transform -1 0 4232 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1190_
timestamp 1688980957
transform -1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1191_
timestamp 1688980957
transform -1 0 4876 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1192_
timestamp 1688980957
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1688980957
transform -1 0 4968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1194_
timestamp 1688980957
transform -1 0 3128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1195_
timestamp 1688980957
transform 1 0 4416 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1196_
timestamp 1688980957
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1197_
timestamp 1688980957
transform 1 0 2300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1198_
timestamp 1688980957
transform 1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1199_
timestamp 1688980957
transform -1 0 3680 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1200_
timestamp 1688980957
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1201_
timestamp 1688980957
transform -1 0 3128 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1202_
timestamp 1688980957
transform 1 0 2116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1203_
timestamp 1688980957
transform 1 0 2116 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1204_
timestamp 1688980957
transform 1 0 2208 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1205_
timestamp 1688980957
transform 1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _1206_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9568 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1207_
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1208_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28520 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1209_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1210_
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1211_
timestamp 1688980957
transform 1 0 29624 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1212_
timestamp 1688980957
transform 1 0 29532 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1213_
timestamp 1688980957
transform 1 0 29808 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1214_
timestamp 1688980957
transform 1 0 30084 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1215_
timestamp 1688980957
transform 1 0 29716 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1216_
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1217_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1218_
timestamp 1688980957
transform 1 0 29440 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1219_
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1220_
timestamp 1688980957
transform 1 0 28796 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1221_
timestamp 1688980957
transform 1 0 28612 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1222_
timestamp 1688980957
transform 1 0 26772 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1223_
timestamp 1688980957
transform 1 0 28336 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1224_
timestamp 1688980957
transform 1 0 8188 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1225_
timestamp 1688980957
transform 1 0 6532 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _1226_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1227_
timestamp 1688980957
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1228_
timestamp 1688980957
transform 1 0 6532 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1229_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1230_
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1231_
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1232_
timestamp 1688980957
transform 1 0 6440 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1233_
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1234_
timestamp 1688980957
transform 1 0 6992 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1235_
timestamp 1688980957
transform 1 0 6440 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1236_
timestamp 1688980957
transform 1 0 6348 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1237_
timestamp 1688980957
transform 1 0 6716 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1238_
timestamp 1688980957
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1239_
timestamp 1688980957
transform 1 0 6992 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1240_
timestamp 1688980957
transform 1 0 6992 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1241_
timestamp 1688980957
transform 1 0 8464 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1242_
timestamp 1688980957
transform 1 0 32108 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1243_
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1244_
timestamp 1688980957
transform 1 0 32476 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1245_
timestamp 1688980957
transform 1 0 32752 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1246_
timestamp 1688980957
transform 1 0 33028 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1247_
timestamp 1688980957
transform 1 0 33028 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1248_
timestamp 1688980957
transform 1 0 33120 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1249_
timestamp 1688980957
transform 1 0 32752 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1250_
timestamp 1688980957
transform 1 0 32752 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1251_
timestamp 1688980957
transform 1 0 33120 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1252_
timestamp 1688980957
transform 1 0 33120 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1253_
timestamp 1688980957
transform 1 0 32752 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1254_
timestamp 1688980957
transform 1 0 32752 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1255_
timestamp 1688980957
transform 1 0 32752 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1256_
timestamp 1688980957
transform 1 0 33120 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1257_
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1258_
timestamp 1688980957
transform 1 0 2852 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1259_
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1260_
timestamp 1688980957
transform 1 0 2760 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1261_
timestamp 1688980957
transform 1 0 2576 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1262_
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1263_
timestamp 1688980957
transform 1 0 1564 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1264_
timestamp 1688980957
transform 1 0 3404 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1265_
timestamp 1688980957
transform 1 0 2576 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1266_
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1267_
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1268_
timestamp 1688980957
transform 1 0 1564 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1269_
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1270_
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1271_
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1272_
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1273_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1274_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A
timestamp 1688980957
transform -1 0 33120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__B1
timestamp 1688980957
transform 1 0 31648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__B1
timestamp 1688980957
transform 1 0 30912 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__B
timestamp 1688980957
transform -1 0 31924 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1688980957
transform -1 0 23644 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__B
timestamp 1688980957
transform -1 0 24288 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1688980957
transform -1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__B
timestamp 1688980957
transform 1 0 22264 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__C
timestamp 1688980957
transform 1 0 22356 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__D
timestamp 1688980957
transform 1 0 21988 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B
timestamp 1688980957
transform 1 0 20884 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__C
timestamp 1688980957
transform -1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__D
timestamp 1688980957
transform 1 0 19964 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1688980957
transform 1 0 21252 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__B
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__C
timestamp 1688980957
transform -1 0 20884 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__D
timestamp 1688980957
transform -1 0 20516 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A
timestamp 1688980957
transform 1 0 20976 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B
timestamp 1688980957
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1688980957
transform 1 0 23368 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__B
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1688980957
transform 1 0 22356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1688980957
transform 1 0 23000 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A1
timestamp 1688980957
transform 1 0 22172 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B2
timestamp 1688980957
transform 1 0 23184 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1688980957
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__B
timestamp 1688980957
transform 1 0 22632 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1688980957
transform -1 0 24748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1688980957
transform 1 0 23552 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B
timestamp 1688980957
transform 1 0 25208 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B
timestamp 1688980957
transform 1 0 22540 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1688980957
transform -1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1688980957
transform 1 0 21712 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1688980957
transform -1 0 23276 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1688980957
transform 1 0 23000 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__B
timestamp 1688980957
transform 1 0 23552 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1688980957
transform -1 0 24104 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A1
timestamp 1688980957
transform -1 0 23920 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A2
timestamp 1688980957
transform -1 0 24012 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A1
timestamp 1688980957
transform 1 0 23000 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A2
timestamp 1688980957
transform 1 0 23368 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1688980957
transform 1 0 21344 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 1688980957
transform -1 0 21896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 1688980957
transform 1 0 20976 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__B
timestamp 1688980957
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1688980957
transform 1 0 17848 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B
timestamp 1688980957
transform 1 0 16100 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__B
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1688980957
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1688980957
transform 1 0 14260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1688980957
transform -1 0 12696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B
timestamp 1688980957
transform 1 0 12144 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1688980957
transform 1 0 14444 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1688980957
transform 1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A
timestamp 1688980957
transform 1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1688980957
transform 1 0 15732 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B
timestamp 1688980957
transform 1 0 15364 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1688980957
transform -1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1688980957
transform 1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1688980957
transform 1 0 14996 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1688980957
transform 1 0 15364 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 1688980957
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__C
timestamp 1688980957
transform -1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__D
timestamp 1688980957
transform -1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__C
timestamp 1688980957
transform 1 0 17388 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__D
timestamp 1688980957
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A
timestamp 1688980957
transform 1 0 21160 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B
timestamp 1688980957
transform 1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A
timestamp 1688980957
transform 1 0 14076 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1688980957
transform 1 0 18676 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__B
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B
timestamp 1688980957
transform 1 0 20056 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A1
timestamp 1688980957
transform -1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A2
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1688980957
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A1
timestamp 1688980957
transform 1 0 13432 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A2
timestamp 1688980957
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A_N
timestamp 1688980957
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B
timestamp 1688980957
transform 1 0 24748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__C
timestamp 1688980957
transform 1 0 25116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__D
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1688980957
transform 1 0 25852 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A2
timestamp 1688980957
transform 1 0 26128 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B1_N
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1_N
timestamp 1688980957
transform -1 0 27140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A
timestamp 1688980957
transform -1 0 23828 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B
timestamp 1688980957
transform 1 0 23644 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__C
timestamp 1688980957
transform 1 0 23276 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A1
timestamp 1688980957
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B1
timestamp 1688980957
transform 1 0 24196 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1
timestamp 1688980957
transform 1 0 26496 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A1
timestamp 1688980957
transform 1 0 26680 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A2
timestamp 1688980957
transform 1 0 25208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B1
timestamp 1688980957
transform 1 0 24840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1688980957
transform -1 0 24288 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__B
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1
timestamp 1688980957
transform 1 0 24656 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1688980957
transform -1 0 26772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B
timestamp 1688980957
transform -1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1688980957
transform -1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B
timestamp 1688980957
transform -1 0 27232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A
timestamp 1688980957
transform 1 0 25392 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B
timestamp 1688980957
transform 1 0 25024 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1688980957
transform -1 0 27968 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B
timestamp 1688980957
transform 1 0 25852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1688980957
transform 1 0 20700 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B
timestamp 1688980957
transform 1 0 20332 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B
timestamp 1688980957
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A
timestamp 1688980957
transform 1 0 20976 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__B
timestamp 1688980957
transform 1 0 20976 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A
timestamp 1688980957
transform 1 0 23184 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B
timestamp 1688980957
transform 1 0 22816 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1688980957
transform -1 0 23460 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2
timestamp 1688980957
transform 1 0 23276 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A
timestamp 1688980957
transform 1 0 21068 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__B
timestamp 1688980957
transform 1 0 14260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1688980957
transform -1 0 11408 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A1
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A3
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1688980957
transform 1 0 12328 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B_N
timestamp 1688980957
transform 1 0 12512 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B1
timestamp 1688980957
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1688980957
transform 1 0 14720 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__B
timestamp 1688980957
transform 1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1688980957
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A2
timestamp 1688980957
transform 1 0 12880 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B1
timestamp 1688980957
transform 1 0 13064 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A_N
timestamp 1688980957
transform 1 0 12788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C
timestamp 1688980957
transform 1 0 13064 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__D
timestamp 1688980957
transform 1 0 12512 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__B
timestamp 1688980957
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A1
timestamp 1688980957
transform -1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A2
timestamp 1688980957
transform 1 0 17940 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B1
timestamp 1688980957
transform 1 0 17572 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1688980957
transform 1 0 17204 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__C
timestamp 1688980957
transform 1 0 16836 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__D
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1688980957
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B_N
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1
timestamp 1688980957
transform -1 0 11408 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A2
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1_N
timestamp 1688980957
transform 1 0 12328 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__B
timestamp 1688980957
transform 1 0 10580 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__C
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__C1
timestamp 1688980957
transform -1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1688980957
transform -1 0 9476 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A2
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B1
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1688980957
transform 1 0 10856 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B
timestamp 1688980957
transform 1 0 8924 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1
timestamp 1688980957
transform -1 0 8832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A_N
timestamp 1688980957
transform 1 0 10120 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B
timestamp 1688980957
transform 1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__C
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__D
timestamp 1688980957
transform 1 0 10488 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A1
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2
timestamp 1688980957
transform 1 0 11132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B1_N
timestamp 1688980957
transform 1 0 10948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1688980957
transform 1 0 10488 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A
timestamp 1688980957
transform 1 0 12328 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B
timestamp 1688980957
transform 1 0 11960 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A1
timestamp 1688980957
transform 1 0 13064 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A2
timestamp 1688980957
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1688980957
transform -1 0 8096 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B
timestamp 1688980957
transform 1 0 8648 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1688980957
transform 1 0 10120 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A1
timestamp 1688980957
transform 1 0 10488 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1688980957
transform 1 0 14720 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B
timestamp 1688980957
transform 1 0 14536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1688980957
transform -1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A
timestamp 1688980957
transform 1 0 14536 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1688980957
transform 1 0 11960 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B
timestamp 1688980957
transform -1 0 10580 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1688980957
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1688980957
transform 1 0 13248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A
timestamp 1688980957
transform 1 0 13156 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1688980957
transform 1 0 12788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__C1
timestamp 1688980957
transform 1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1688980957
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1688980957
transform -1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1688980957
transform 1 0 15088 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B
timestamp 1688980957
transform 1 0 15732 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1688980957
transform 1 0 10304 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B
timestamp 1688980957
transform 1 0 10672 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1688980957
transform 1 0 9292 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B
timestamp 1688980957
transform -1 0 9660 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__C
timestamp 1688980957
transform 1 0 8924 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__D
timestamp 1688980957
transform -1 0 8464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1688980957
transform 1 0 13340 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A
timestamp 1688980957
transform 1 0 14352 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B
timestamp 1688980957
transform 1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A
timestamp 1688980957
transform 1 0 10672 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1688980957
transform 1 0 10304 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1688980957
transform 1 0 11960 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1688980957
transform 1 0 11132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1688980957
transform 1 0 11684 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B
timestamp 1688980957
transform 1 0 26128 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1688980957
transform 1 0 25208 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B
timestamp 1688980957
transform 1 0 25024 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1688980957
transform 1 0 17480 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__B
timestamp 1688980957
transform 1 0 18124 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1688980957
transform 1 0 16928 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1688980957
transform 1 0 14996 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__B
timestamp 1688980957
transform -1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1688980957
transform 1 0 14996 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B_N
timestamp 1688980957
transform -1 0 13156 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1688980957
transform -1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A
timestamp 1688980957
transform -1 0 13984 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A1
timestamp 1688980957
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1688980957
transform 1 0 20056 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__B
timestamp 1688980957
transform 1 0 19872 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1688980957
transform 1 0 20516 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B2
timestamp 1688980957
transform 1 0 20148 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1688980957
transform 1 0 20516 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A1_N
timestamp 1688980957
transform 1 0 21712 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2_N
timestamp 1688980957
transform 1 0 21436 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A1
timestamp 1688980957
transform 1 0 21620 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A1
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A2
timestamp 1688980957
transform 1 0 17664 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A3
timestamp 1688980957
transform 1 0 17296 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A4
timestamp 1688980957
transform 1 0 16928 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1688980957
transform 1 0 17480 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A
timestamp 1688980957
transform -1 0 16100 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B
timestamp 1688980957
transform -1 0 15456 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A1
timestamp 1688980957
transform 1 0 16008 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B1
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A1
timestamp 1688980957
transform 1 0 16008 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1688980957
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A1
timestamp 1688980957
transform 1 0 17480 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__B1
timestamp 1688980957
transform 1 0 16928 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B1
timestamp 1688980957
transform -1 0 15456 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__A
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A1
timestamp 1688980957
transform 1 0 20792 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__S
timestamp 1688980957
transform -1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1688980957
transform -1 0 19596 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B2
timestamp 1688980957
transform 1 0 19872 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1688980957
transform -1 0 26220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__B
timestamp 1688980957
transform -1 0 26864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1688980957
transform -1 0 25300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__B
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__A
timestamp 1688980957
transform -1 0 22264 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__C
timestamp 1688980957
transform 1 0 21344 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A1
timestamp 1688980957
transform 1 0 19412 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A2
timestamp 1688980957
transform 1 0 18676 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__B2
timestamp 1688980957
transform 1 0 18860 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1688980957
transform -1 0 22172 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A3
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A1
timestamp 1688980957
transform -1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1688980957
transform -1 0 28980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A
timestamp 1688980957
transform 1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__A
timestamp 1688980957
transform 1 0 10120 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1688980957
transform -1 0 29164 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__A
timestamp 1688980957
transform 1 0 29992 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A
timestamp 1688980957
transform 1 0 30084 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A
timestamp 1688980957
transform 1 0 31280 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__A
timestamp 1688980957
transform 1 0 30268 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1688980957
transform 1 0 30544 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__A
timestamp 1688980957
transform 1 0 30452 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1688980957
transform 1 0 29992 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1688980957
transform 1 0 31188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A
timestamp 1688980957
transform 1 0 30268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__A
timestamp 1688980957
transform 1 0 29624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A
timestamp 1688980957
transform 1 0 29808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1688980957
transform 1 0 30084 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__A
timestamp 1688980957
transform 1 0 28244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__A
timestamp 1688980957
transform 1 0 29992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1688980957
transform 1 0 10212 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A
timestamp 1688980957
transform 1 0 28060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1688980957
transform 1 0 8648 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__A
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A
timestamp 1688980957
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__A
timestamp 1688980957
transform 1 0 8004 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1688980957
transform 1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A
timestamp 1688980957
transform 1 0 7820 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__A
timestamp 1688980957
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A
timestamp 1688980957
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1688980957
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__A
timestamp 1688980957
transform 1 0 7544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__A
timestamp 1688980957
transform -1 0 8832 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__A
timestamp 1688980957
transform -1 0 7452 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__A
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__A
timestamp 1688980957
transform 1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__A
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__A
timestamp 1688980957
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1688980957
transform 1 0 10580 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__A
timestamp 1688980957
transform -1 0 34592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__A
timestamp 1688980957
transform 1 0 32476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1688980957
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A
timestamp 1688980957
transform -1 0 34960 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__A
timestamp 1688980957
transform -1 0 34684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1688980957
transform 1 0 33488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A
timestamp 1688980957
transform 1 0 33856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A
timestamp 1688980957
transform 1 0 33856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A
timestamp 1688980957
transform 1 0 34132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__A
timestamp 1688980957
transform 1 0 34500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__A
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A
timestamp 1688980957
transform 1 0 34500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1688980957
transform 1 0 34500 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A
timestamp 1688980957
transform 1 0 34592 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__A
timestamp 1688980957
transform 1 0 34132 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A
timestamp 1688980957
transform -1 0 32844 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1688980957
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A
timestamp 1688980957
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A
timestamp 1688980957
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1688980957
transform 1 0 4232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A
timestamp 1688980957
transform 1 0 4968 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A
timestamp 1688980957
transform -1 0 4140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A
timestamp 1688980957
transform 1 0 4232 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A
timestamp 1688980957
transform 1 0 4232 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A
timestamp 1688980957
transform -1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__A
timestamp 1688980957
transform 1 0 2024 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1688980957
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__A
timestamp 1688980957
transform 1 0 2668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A
timestamp 1688980957
transform 1 0 3312 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A
timestamp 1688980957
transform -1 0 2116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1688980957
transform 1 0 2576 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1688980957
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1688980957
transform 1 0 11500 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1688980957
transform 1 0 11040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1688980957
transform 1 0 28336 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1688980957
transform 1 0 29256 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1688980957
transform 1 0 29348 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1688980957
transform 1 0 29440 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1688980957
transform 1 0 29348 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1688980957
transform 1 0 29624 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1688980957
transform 1 0 29900 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1688980957
transform 1 0 29532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1688980957
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1688980957
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1688980957
transform 1 0 29256 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1688980957
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1688980957
transform 1 0 28612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1688980957
transform 1 0 28428 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__CLK
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__CLK
timestamp 1688980957
transform 1 0 28152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1688980957
transform 1 0 9016 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1688980957
transform 1 0 10212 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1688980957
transform 1 0 8372 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1688980957
transform 1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__CLK
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__CLK
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__CLK
timestamp 1688980957
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__CLK
timestamp 1688980957
transform 1 0 9108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__CLK
timestamp 1688980957
transform 1 0 9016 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1234__CLK
timestamp 1688980957
transform 1 0 9108 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__CLK
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__CLK
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1237__CLK
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__CLK
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__CLK
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1240__CLK
timestamp 1688980957
transform 1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__CLK
timestamp 1688980957
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__CLK
timestamp 1688980957
transform 1 0 31924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__CLK
timestamp 1688980957
transform 1 0 31832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__CLK
timestamp 1688980957
transform 1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1245__CLK
timestamp 1688980957
transform 1 0 32568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__CLK
timestamp 1688980957
transform 1 0 32844 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__CLK
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__CLK
timestamp 1688980957
transform 1 0 32936 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__CLK
timestamp 1688980957
transform 1 0 32568 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__CLK
timestamp 1688980957
transform 1 0 32568 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__CLK
timestamp 1688980957
transform 1 0 32936 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__CLK
timestamp 1688980957
transform 1 0 32936 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__CLK
timestamp 1688980957
transform 1 0 32568 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__CLK
timestamp 1688980957
transform 1 0 32568 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__CLK
timestamp 1688980957
transform 1 0 32568 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__CLK
timestamp 1688980957
transform 1 0 32936 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__CLK
timestamp 1688980957
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__CLK
timestamp 1688980957
transform 1 0 4876 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__CLK
timestamp 1688980957
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__CLK
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__CLK
timestamp 1688980957
transform 1 0 4600 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__CLK
timestamp 1688980957
transform 1 0 4692 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__CLK
timestamp 1688980957
transform 1 0 3404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__CLK
timestamp 1688980957
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__CLK
timestamp 1688980957
transform 1 0 4600 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__CLK
timestamp 1688980957
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__CLK
timestamp 1688980957
transform 1 0 3404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__CLK
timestamp 1688980957
transform 1 0 3404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__CLK
timestamp 1688980957
transform 1 0 3404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__CLK
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__CLK
timestamp 1688980957
transform 1 0 3404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__CLK
timestamp 1688980957
transform 1 0 3404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__CLK
timestamp 1688980957
transform 1 0 3036 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__CLK
timestamp 1688980957
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_max_cap49_A
timestamp 1688980957
transform 1 0 32660 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_103
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_281 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_288
timestamp 1688980957
transform 1 0 27600 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_300
timestamp 1688980957
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_367
timestamp 1688980957
transform 1 0 34868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_367
timestamp 1688980957
transform 1 0 34868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_367
timestamp 1688980957
transform 1 0 34868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_367
timestamp 1688980957
transform 1 0 34868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 1688980957
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1688980957
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_367
timestamp 1688980957
transform 1 0 34868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_367
timestamp 1688980957
transform 1 0 34868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_181
timestamp 1688980957
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_202
timestamp 1688980957
transform 1 0 19688 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_214
timestamp 1688980957
transform 1 0 20792 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_226
timestamp 1688980957
transform 1 0 21896 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_238
timestamp 1688980957
transform 1 0 23000 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_11
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_16
timestamp 1688980957
transform 1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_20
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_32
timestamp 1688980957
transform 1 0 4048 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_44
timestamp 1688980957
transform 1 0 5152 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_214
timestamp 1688980957
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_333
timestamp 1688980957
transform 1 0 31740 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_360
timestamp 1688980957
transform 1 0 34224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_364
timestamp 1688980957
transform 1 0 34592 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_24
timestamp 1688980957
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_178
timestamp 1688980957
transform 1 0 17480 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_182
timestamp 1688980957
transform 1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_193
timestamp 1688980957
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_205
timestamp 1688980957
transform 1 0 19964 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_214
timestamp 1688980957
transform 1 0 20792 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_231
timestamp 1688980957
transform 1 0 22356 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_243
timestamp 1688980957
transform 1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_291
timestamp 1688980957
transform 1 0 27876 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_295
timestamp 1688980957
transform 1 0 28244 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_327
timestamp 1688980957
transform 1 0 31188 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_331
timestamp 1688980957
transform 1 0 31556 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_335
timestamp 1688980957
transform 1 0 31924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_339
timestamp 1688980957
transform 1 0 32292 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_346
timestamp 1688980957
transform 1 0 32936 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_6
timestamp 1688980957
transform 1 0 1656 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_18
timestamp 1688980957
transform 1 0 2760 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_43
timestamp 1688980957
transform 1 0 5060 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_47
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_79
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_84
timestamp 1688980957
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_88
timestamp 1688980957
transform 1 0 9200 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_100
timestamp 1688980957
transform 1 0 10304 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_184
timestamp 1688980957
transform 1 0 18032 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_196
timestamp 1688980957
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_208
timestamp 1688980957
transform 1 0 20240 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_214
timestamp 1688980957
transform 1 0 20792 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_241
timestamp 1688980957
transform 1 0 23276 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_255
timestamp 1688980957
transform 1 0 24564 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_267
timestamp 1688980957
transform 1 0 25668 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_331
timestamp 1688980957
transform 1 0 31556 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_365
timestamp 1688980957
transform 1 0 34684 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_24
timestamp 1688980957
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_34
timestamp 1688980957
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_38
timestamp 1688980957
transform 1 0 4600 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_50
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_58
timestamp 1688980957
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_105
timestamp 1688980957
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_161
timestamp 1688980957
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_171
timestamp 1688980957
transform 1 0 16836 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_220
timestamp 1688980957
transform 1 0 21344 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_226
timestamp 1688980957
transform 1 0 21896 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_263
timestamp 1688980957
transform 1 0 25300 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_273
timestamp 1688980957
transform 1 0 26220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_299
timestamp 1688980957
transform 1 0 28612 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_303
timestamp 1688980957
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_317
timestamp 1688980957
transform 1 0 30268 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_328
timestamp 1688980957
transform 1 0 31280 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_336
timestamp 1688980957
transform 1 0 32016 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_14
timestamp 1688980957
transform 1 0 2392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_18
timestamp 1688980957
transform 1 0 2760 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_42
timestamp 1688980957
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_46
timestamp 1688980957
transform 1 0 5336 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_50
timestamp 1688980957
transform 1 0 5704 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_119
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_122
timestamp 1688980957
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_131
timestamp 1688980957
transform 1 0 13156 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_136
timestamp 1688980957
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_140
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_150
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_155
timestamp 1688980957
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_178
timestamp 1688980957
transform 1 0 17480 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_208
timestamp 1688980957
transform 1 0 20240 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_259
timestamp 1688980957
transform 1 0 24932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_276
timestamp 1688980957
transform 1 0 26496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_364
timestamp 1688980957
transform 1 0 34592 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_37
timestamp 1688980957
transform 1 0 4508 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_40
timestamp 1688980957
transform 1 0 4784 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_48
timestamp 1688980957
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_57
timestamp 1688980957
transform 1 0 6348 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_89
timestamp 1688980957
transform 1 0 9292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_117
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_179
timestamp 1688980957
transform 1 0 17572 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_192
timestamp 1688980957
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_201
timestamp 1688980957
transform 1 0 19596 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_214
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_223
timestamp 1688980957
transform 1 0 21620 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_231
timestamp 1688980957
transform 1 0 22356 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_243
timestamp 1688980957
transform 1 0 23460 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_266
timestamp 1688980957
transform 1 0 25576 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_278
timestamp 1688980957
transform 1 0 26680 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_293
timestamp 1688980957
transform 1 0 28060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_297
timestamp 1688980957
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_313
timestamp 1688980957
transform 1 0 29900 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_317
timestamp 1688980957
transform 1 0 30268 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_323
timestamp 1688980957
transform 1 0 30820 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_330
timestamp 1688980957
transform 1 0 31464 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_334
timestamp 1688980957
transform 1 0 31832 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_346
timestamp 1688980957
transform 1 0 32936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_6
timestamp 1688980957
transform 1 0 1656 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_41
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_52
timestamp 1688980957
transform 1 0 5888 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_78
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_82
timestamp 1688980957
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_86
timestamp 1688980957
transform 1 0 9016 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_90
timestamp 1688980957
transform 1 0 9384 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_98
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_101
timestamp 1688980957
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_109
timestamp 1688980957
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_121
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_129
timestamp 1688980957
transform 1 0 12972 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_133
timestamp 1688980957
transform 1 0 13340 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_136
timestamp 1688980957
transform 1 0 13616 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_155
timestamp 1688980957
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_159
timestamp 1688980957
transform 1 0 15732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_174
timestamp 1688980957
transform 1 0 17112 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_179
timestamp 1688980957
transform 1 0 17572 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_183
timestamp 1688980957
transform 1 0 17940 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_189
timestamp 1688980957
transform 1 0 18492 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_197
timestamp 1688980957
transform 1 0 19228 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_203
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_207
timestamp 1688980957
transform 1 0 20148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_212
timestamp 1688980957
transform 1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_216
timestamp 1688980957
transform 1 0 20976 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_220
timestamp 1688980957
transform 1 0 21344 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_291
timestamp 1688980957
transform 1 0 27876 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_319
timestamp 1688980957
transform 1 0 30452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_331
timestamp 1688980957
transform 1 0 31556 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_367
timestamp 1688980957
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_23
timestamp 1688980957
transform 1 0 3220 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_44
timestamp 1688980957
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_56
timestamp 1688980957
transform 1 0 6256 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_88
timestamp 1688980957
transform 1 0 9200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_124
timestamp 1688980957
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_128
timestamp 1688980957
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_132
timestamp 1688980957
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_136
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_147
timestamp 1688980957
transform 1 0 14628 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_157
timestamp 1688980957
transform 1 0 15548 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_161
timestamp 1688980957
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_174
timestamp 1688980957
transform 1 0 17112 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_186
timestamp 1688980957
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_190
timestamp 1688980957
transform 1 0 18584 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_206
timestamp 1688980957
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_223
timestamp 1688980957
transform 1 0 21620 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_227
timestamp 1688980957
transform 1 0 21988 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_243
timestamp 1688980957
transform 1 0 23460 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_288
timestamp 1688980957
transform 1 0 27600 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_297
timestamp 1688980957
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_305
timestamp 1688980957
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_322
timestamp 1688980957
transform 1 0 30728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_344
timestamp 1688980957
transform 1 0 32752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_348
timestamp 1688980957
transform 1 0 33120 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_354
timestamp 1688980957
transform 1 0 33672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_63
timestamp 1688980957
transform 1 0 6900 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_75
timestamp 1688980957
transform 1 0 8004 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_84
timestamp 1688980957
transform 1 0 8832 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_88
timestamp 1688980957
transform 1 0 9200 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_92
timestamp 1688980957
transform 1 0 9568 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_96
timestamp 1688980957
transform 1 0 9936 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_100
timestamp 1688980957
transform 1 0 10304 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_121
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_131
timestamp 1688980957
transform 1 0 13156 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_135
timestamp 1688980957
transform 1 0 13524 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_138
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_143
timestamp 1688980957
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_150
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_155
timestamp 1688980957
transform 1 0 15364 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_165
timestamp 1688980957
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_196
timestamp 1688980957
transform 1 0 19136 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_206
timestamp 1688980957
transform 1 0 20056 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_229
timestamp 1688980957
transform 1 0 22172 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_240
timestamp 1688980957
transform 1 0 23184 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_252
timestamp 1688980957
transform 1 0 24288 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_258
timestamp 1688980957
transform 1 0 24840 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_292
timestamp 1688980957
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_304
timestamp 1688980957
transform 1 0 29072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_328
timestamp 1688980957
transform 1 0 31280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_344
timestamp 1688980957
transform 1 0 32752 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_367
timestamp 1688980957
transform 1 0 34868 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_32
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_36
timestamp 1688980957
transform 1 0 4416 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_47
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_106
timestamp 1688980957
transform 1 0 10856 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_110
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_123
timestamp 1688980957
transform 1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_127
timestamp 1688980957
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_131
timestamp 1688980957
transform 1 0 13156 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_135
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_145
timestamp 1688980957
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_148
timestamp 1688980957
transform 1 0 14720 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_154
timestamp 1688980957
transform 1 0 15272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_157
timestamp 1688980957
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_161
timestamp 1688980957
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_174
timestamp 1688980957
transform 1 0 17112 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_180
timestamp 1688980957
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_184
timestamp 1688980957
transform 1 0 18032 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_192
timestamp 1688980957
transform 1 0 18768 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_201
timestamp 1688980957
transform 1 0 19596 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_226
timestamp 1688980957
transform 1 0 21896 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_249
timestamp 1688980957
transform 1 0 24012 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_271
timestamp 1688980957
transform 1 0 26036 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_279
timestamp 1688980957
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_286
timestamp 1688980957
transform 1 0 27416 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_297
timestamp 1688980957
transform 1 0 28428 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_305
timestamp 1688980957
transform 1 0 29164 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_329
timestamp 1688980957
transform 1 0 31372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_335
timestamp 1688980957
transform 1 0 31924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_339
timestamp 1688980957
transform 1 0 32292 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_347
timestamp 1688980957
transform 1 0 33028 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_6
timestamp 1688980957
transform 1 0 1656 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_18
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_75
timestamp 1688980957
transform 1 0 8004 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_88
timestamp 1688980957
transform 1 0 9200 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_100
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_106
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_145
timestamp 1688980957
transform 1 0 14444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_174
timestamp 1688980957
transform 1 0 17112 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_180
timestamp 1688980957
transform 1 0 17664 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_192
timestamp 1688980957
transform 1 0 18768 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_198
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_211
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_215
timestamp 1688980957
transform 1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_244
timestamp 1688980957
transform 1 0 23552 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_266
timestamp 1688980957
transform 1 0 25576 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_297
timestamp 1688980957
transform 1 0 28428 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_309
timestamp 1688980957
transform 1 0 29532 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_315
timestamp 1688980957
transform 1 0 30084 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_341
timestamp 1688980957
transform 1 0 32476 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_345
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_357
timestamp 1688980957
transform 1 0 33948 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_365
timestamp 1688980957
transform 1 0 34684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_33
timestamp 1688980957
transform 1 0 4140 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_37
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_47
timestamp 1688980957
transform 1 0 5428 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_76
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_80
timestamp 1688980957
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_91
timestamp 1688980957
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_113
timestamp 1688980957
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_122
timestamp 1688980957
transform 1 0 12328 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_168
timestamp 1688980957
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_172
timestamp 1688980957
transform 1 0 16928 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_175
timestamp 1688980957
transform 1 0 17204 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_179
timestamp 1688980957
transform 1 0 17572 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_183
timestamp 1688980957
transform 1 0 17940 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_188
timestamp 1688980957
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_192
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_204
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_208
timestamp 1688980957
transform 1 0 20240 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_218
timestamp 1688980957
transform 1 0 21160 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_222
timestamp 1688980957
transform 1 0 21528 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_234
timestamp 1688980957
transform 1 0 22632 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_240
timestamp 1688980957
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_259
timestamp 1688980957
transform 1 0 24932 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_262
timestamp 1688980957
transform 1 0 25208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_266
timestamp 1688980957
transform 1 0 25576 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_271
timestamp 1688980957
transform 1 0 26036 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_279
timestamp 1688980957
transform 1 0 26772 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_283
timestamp 1688980957
transform 1 0 27140 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_295
timestamp 1688980957
transform 1 0 28244 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_303
timestamp 1688980957
transform 1 0 28980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_332
timestamp 1688980957
transform 1 0 31648 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_343
timestamp 1688980957
transform 1 0 32660 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_355
timestamp 1688980957
transform 1 0 33764 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_361
timestamp 1688980957
transform 1 0 34316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_47
timestamp 1688980957
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_100
timestamp 1688980957
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_108
timestamp 1688980957
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_132
timestamp 1688980957
transform 1 0 13248 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_142
timestamp 1688980957
transform 1 0 14168 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_150
timestamp 1688980957
transform 1 0 14904 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_156
timestamp 1688980957
transform 1 0 15456 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_177
timestamp 1688980957
transform 1 0 17388 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_214
timestamp 1688980957
transform 1 0 20792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_221
timestamp 1688980957
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_232
timestamp 1688980957
transform 1 0 22448 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_240
timestamp 1688980957
transform 1 0 23184 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_243
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_255
timestamp 1688980957
transform 1 0 24564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_260
timestamp 1688980957
transform 1 0 25024 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_316
timestamp 1688980957
transform 1 0 30176 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_328
timestamp 1688980957
transform 1 0 31280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_342
timestamp 1688980957
transform 1 0 32568 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_36
timestamp 1688980957
transform 1 0 4416 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_48
timestamp 1688980957
transform 1 0 5520 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_60
timestamp 1688980957
transform 1 0 6624 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_71
timestamp 1688980957
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_75
timestamp 1688980957
transform 1 0 8004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1688980957
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_101
timestamp 1688980957
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_105
timestamp 1688980957
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_116
timestamp 1688980957
transform 1 0 11776 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_120
timestamp 1688980957
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_124
timestamp 1688980957
transform 1 0 12512 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_134
timestamp 1688980957
transform 1 0 13432 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_149
timestamp 1688980957
transform 1 0 14812 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_161
timestamp 1688980957
transform 1 0 15916 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_167
timestamp 1688980957
transform 1 0 16468 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_181
timestamp 1688980957
transform 1 0 17756 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_185
timestamp 1688980957
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_201
timestamp 1688980957
transform 1 0 19596 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_213
timestamp 1688980957
transform 1 0 20700 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_225
timestamp 1688980957
transform 1 0 21804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_239
timestamp 1688980957
transform 1 0 23092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_243
timestamp 1688980957
transform 1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_276
timestamp 1688980957
transform 1 0 26496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_280
timestamp 1688980957
transform 1 0 26864 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_284
timestamp 1688980957
transform 1 0 27232 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_288
timestamp 1688980957
transform 1 0 27600 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_292
timestamp 1688980957
transform 1 0 27968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_304
timestamp 1688980957
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_312
timestamp 1688980957
transform 1 0 29808 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_316
timestamp 1688980957
transform 1 0 30176 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_328
timestamp 1688980957
transform 1 0 31280 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_340
timestamp 1688980957
transform 1 0 32384 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_6
timestamp 1688980957
transform 1 0 1656 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_19
timestamp 1688980957
transform 1 0 2852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_36
timestamp 1688980957
transform 1 0 4416 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_50
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_94
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_98
timestamp 1688980957
transform 1 0 10120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_102
timestamp 1688980957
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_122
timestamp 1688980957
transform 1 0 12328 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_130
timestamp 1688980957
transform 1 0 13064 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_154
timestamp 1688980957
transform 1 0 15272 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_188
timestamp 1688980957
transform 1 0 18400 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_200
timestamp 1688980957
transform 1 0 19504 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_208
timestamp 1688980957
transform 1 0 20240 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_238
timestamp 1688980957
transform 1 0 23000 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_258
timestamp 1688980957
transform 1 0 24840 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_275
timestamp 1688980957
transform 1 0 26404 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_287
timestamp 1688980957
transform 1 0 27508 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_299
timestamp 1688980957
transform 1 0 28612 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_311
timestamp 1688980957
transform 1 0 29716 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_323
timestamp 1688980957
transform 1 0 30820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_47
timestamp 1688980957
transform 1 0 5428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_55
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_81
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_105
timestamp 1688980957
transform 1 0 10764 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_123
timestamp 1688980957
transform 1 0 12420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_127
timestamp 1688980957
transform 1 0 12788 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_144
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_148
timestamp 1688980957
transform 1 0 14720 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_168
timestamp 1688980957
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_175
timestamp 1688980957
transform 1 0 17204 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_210
timestamp 1688980957
transform 1 0 20424 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_214
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_226
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_234
timestamp 1688980957
transform 1 0 22632 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_238
timestamp 1688980957
transform 1 0 23000 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_242
timestamp 1688980957
transform 1 0 23368 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_247
timestamp 1688980957
transform 1 0 23828 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_263
timestamp 1688980957
transform 1 0 25300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_267
timestamp 1688980957
transform 1 0 25668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_271
timestamp 1688980957
transform 1 0 26036 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_275
timestamp 1688980957
transform 1 0 26404 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_279
timestamp 1688980957
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_291
timestamp 1688980957
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_303
timestamp 1688980957
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_35
timestamp 1688980957
transform 1 0 4324 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_77
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_85
timestamp 1688980957
transform 1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_89
timestamp 1688980957
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_103
timestamp 1688980957
transform 1 0 10580 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_126
timestamp 1688980957
transform 1 0 12696 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1688980957
transform 1 0 15088 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_187
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_243
timestamp 1688980957
transform 1 0 23460 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_255
timestamp 1688980957
transform 1 0 24564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_259
timestamp 1688980957
transform 1 0 24932 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_263
timestamp 1688980957
transform 1 0 25300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_270
timestamp 1688980957
transform 1 0 25944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_274
timestamp 1688980957
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_313
timestamp 1688980957
transform 1 0 29900 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_319
timestamp 1688980957
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_331
timestamp 1688980957
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_341
timestamp 1688980957
transform 1 0 32476 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_344
timestamp 1688980957
transform 1 0 32752 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_35
timestamp 1688980957
transform 1 0 4324 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_43
timestamp 1688980957
transform 1 0 5060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_49
timestamp 1688980957
transform 1 0 5612 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_57
timestamp 1688980957
transform 1 0 6348 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_79
timestamp 1688980957
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_101
timestamp 1688980957
transform 1 0 10396 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_105
timestamp 1688980957
transform 1 0 10764 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_116
timestamp 1688980957
transform 1 0 11776 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_120
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_124
timestamp 1688980957
transform 1 0 12512 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_129
timestamp 1688980957
transform 1 0 12972 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_138
timestamp 1688980957
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_190
timestamp 1688980957
transform 1 0 18584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_194
timestamp 1688980957
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_248
timestamp 1688980957
transform 1 0 23920 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_259
timestamp 1688980957
transform 1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_279
timestamp 1688980957
transform 1 0 26772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_283
timestamp 1688980957
transform 1 0 27140 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_302
timestamp 1688980957
transform 1 0 28888 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_329
timestamp 1688980957
transform 1 0 31372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_343
timestamp 1688980957
transform 1 0 32660 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_29
timestamp 1688980957
transform 1 0 3772 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_40
timestamp 1688980957
transform 1 0 4784 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_82
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_124
timestamp 1688980957
transform 1 0 12512 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_129
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_133
timestamp 1688980957
transform 1 0 13340 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_145
timestamp 1688980957
transform 1 0 14444 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_153
timestamp 1688980957
transform 1 0 15180 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_164
timestamp 1688980957
transform 1 0 16192 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_174
timestamp 1688980957
transform 1 0 17112 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_178
timestamp 1688980957
transform 1 0 17480 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_182
timestamp 1688980957
transform 1 0 17848 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_197
timestamp 1688980957
transform 1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_208
timestamp 1688980957
transform 1 0 20240 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_234
timestamp 1688980957
transform 1 0 22632 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_238
timestamp 1688980957
transform 1 0 23000 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_246
timestamp 1688980957
transform 1 0 23736 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_250
timestamp 1688980957
transform 1 0 24104 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_253
timestamp 1688980957
transform 1 0 24380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_259
timestamp 1688980957
transform 1 0 24932 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_264
timestamp 1688980957
transform 1 0 25392 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_270
timestamp 1688980957
transform 1 0 25944 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_274
timestamp 1688980957
transform 1 0 26312 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_278
timestamp 1688980957
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_311
timestamp 1688980957
transform 1 0 29716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_324
timestamp 1688980957
transform 1 0 30912 0 -1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_342
timestamp 1688980957
transform 1 0 32568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_354
timestamp 1688980957
transform 1 0 33672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_358
timestamp 1688980957
transform 1 0 34040 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_365
timestamp 1688980957
transform 1 0 34684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_6
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_38
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_46
timestamp 1688980957
transform 1 0 5336 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_58
timestamp 1688980957
transform 1 0 6440 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_73
timestamp 1688980957
transform 1 0 7820 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_100
timestamp 1688980957
transform 1 0 10304 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_126
timestamp 1688980957
transform 1 0 12696 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_145
timestamp 1688980957
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_149
timestamp 1688980957
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_159
timestamp 1688980957
transform 1 0 15732 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_176
timestamp 1688980957
transform 1 0 17296 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_184
timestamp 1688980957
transform 1 0 18032 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_192
timestamp 1688980957
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_214
timestamp 1688980957
transform 1 0 20792 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_226
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_236
timestamp 1688980957
transform 1 0 22816 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_257
timestamp 1688980957
transform 1 0 24748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_262
timestamp 1688980957
transform 1 0 25208 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_283
timestamp 1688980957
transform 1 0 27140 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_287
timestamp 1688980957
transform 1 0 27508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_292
timestamp 1688980957
transform 1 0 27968 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_298
timestamp 1688980957
transform 1 0 28520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_306
timestamp 1688980957
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_331
timestamp 1688980957
transform 1 0 31556 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_340
timestamp 1688980957
transform 1 0 32384 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_11
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_22
timestamp 1688980957
transform 1 0 3128 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_26
timestamp 1688980957
transform 1 0 3496 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_38
timestamp 1688980957
transform 1 0 4600 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 1688980957
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_83
timestamp 1688980957
transform 1 0 8740 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_91
timestamp 1688980957
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_96
timestamp 1688980957
transform 1 0 9936 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_100
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_104
timestamp 1688980957
transform 1 0 10672 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_108
timestamp 1688980957
transform 1 0 11040 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_132
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_146
timestamp 1688980957
transform 1 0 14536 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_150
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_159
timestamp 1688980957
transform 1 0 15732 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_165
timestamp 1688980957
transform 1 0 16284 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_180
timestamp 1688980957
transform 1 0 17664 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_192
timestamp 1688980957
transform 1 0 18768 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_204
timestamp 1688980957
transform 1 0 19872 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_211
timestamp 1688980957
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_233
timestamp 1688980957
transform 1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_241
timestamp 1688980957
transform 1 0 23276 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_248
timestamp 1688980957
transform 1 0 23920 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_255
timestamp 1688980957
transform 1 0 24564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_264
timestamp 1688980957
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_271
timestamp 1688980957
transform 1 0 26036 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_275
timestamp 1688980957
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_296
timestamp 1688980957
transform 1 0 28336 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_303
timestamp 1688980957
transform 1 0 28980 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_315
timestamp 1688980957
transform 1 0 30084 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_327
timestamp 1688980957
transform 1 0 31188 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_367
timestamp 1688980957
transform 1 0 34868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_23
timestamp 1688980957
transform 1 0 3220 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_56
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_81
timestamp 1688980957
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_89
timestamp 1688980957
transform 1 0 9292 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_100
timestamp 1688980957
transform 1 0 10304 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_120
timestamp 1688980957
transform 1 0 12144 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_126
timestamp 1688980957
transform 1 0 12696 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_146
timestamp 1688980957
transform 1 0 14536 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_158
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_166
timestamp 1688980957
transform 1 0 16376 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_190
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_217
timestamp 1688980957
transform 1 0 21068 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_223
timestamp 1688980957
transform 1 0 21620 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_239
timestamp 1688980957
transform 1 0 23092 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_260
timestamp 1688980957
transform 1 0 25024 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_264
timestamp 1688980957
transform 1 0 25392 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_280
timestamp 1688980957
transform 1 0 26864 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_292
timestamp 1688980957
transform 1 0 27968 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_304
timestamp 1688980957
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_14
timestamp 1688980957
transform 1 0 2392 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_18
timestamp 1688980957
transform 1 0 2760 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_62
timestamp 1688980957
transform 1 0 6808 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_102
timestamp 1688980957
transform 1 0 10488 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_108
timestamp 1688980957
transform 1 0 11040 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_126
timestamp 1688980957
transform 1 0 12696 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_132
timestamp 1688980957
transform 1 0 13248 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_136
timestamp 1688980957
transform 1 0 13616 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_144
timestamp 1688980957
transform 1 0 14352 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_176
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_188
timestamp 1688980957
transform 1 0 18400 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_203
timestamp 1688980957
transform 1 0 19780 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_215
timestamp 1688980957
transform 1 0 20884 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_235
timestamp 1688980957
transform 1 0 22724 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_240
timestamp 1688980957
transform 1 0 23184 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_244
timestamp 1688980957
transform 1 0 23552 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_256
timestamp 1688980957
transform 1 0 24656 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_268
timestamp 1688980957
transform 1 0 25760 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_272
timestamp 1688980957
transform 1 0 26128 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_297
timestamp 1688980957
transform 1 0 28428 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_309
timestamp 1688980957
transform 1 0 29532 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_321
timestamp 1688980957
transform 1 0 30636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_6
timestamp 1688980957
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_18
timestamp 1688980957
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_32
timestamp 1688980957
transform 1 0 4048 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_36
timestamp 1688980957
transform 1 0 4416 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_56
timestamp 1688980957
transform 1 0 6256 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_68
timestamp 1688980957
transform 1 0 7360 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_78
timestamp 1688980957
transform 1 0 8280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_100
timestamp 1688980957
transform 1 0 10304 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_131
timestamp 1688980957
transform 1 0 13156 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_136
timestamp 1688980957
transform 1 0 13616 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_149
timestamp 1688980957
transform 1 0 14812 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_156
timestamp 1688980957
transform 1 0 15456 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_168
timestamp 1688980957
transform 1 0 16560 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_176
timestamp 1688980957
transform 1 0 17296 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_185
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_212
timestamp 1688980957
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_216
timestamp 1688980957
transform 1 0 20976 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_222
timestamp 1688980957
transform 1 0 21528 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_226
timestamp 1688980957
transform 1 0 21896 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_230
timestamp 1688980957
transform 1 0 22264 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_239
timestamp 1688980957
transform 1 0 23092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_279
timestamp 1688980957
transform 1 0 26772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_302
timestamp 1688980957
transform 1 0 28888 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_319
timestamp 1688980957
transform 1 0 30452 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_326
timestamp 1688980957
transform 1 0 31096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_339
timestamp 1688980957
transform 1 0 32292 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_348
timestamp 1688980957
transform 1 0 33120 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_356
timestamp 1688980957
transform 1 0 33856 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_362
timestamp 1688980957
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_14
timestamp 1688980957
transform 1 0 2392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_36
timestamp 1688980957
transform 1 0 4416 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_40
timestamp 1688980957
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_52
timestamp 1688980957
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_65
timestamp 1688980957
transform 1 0 7084 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_72
timestamp 1688980957
transform 1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_77
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_83
timestamp 1688980957
transform 1 0 8740 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_87
timestamp 1688980957
transform 1 0 9108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_91
timestamp 1688980957
transform 1 0 9476 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_100
timestamp 1688980957
transform 1 0 10304 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_104
timestamp 1688980957
transform 1 0 10672 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_108
timestamp 1688980957
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_117
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_120
timestamp 1688980957
transform 1 0 12144 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_129
timestamp 1688980957
transform 1 0 12972 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_144
timestamp 1688980957
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_148
timestamp 1688980957
transform 1 0 14720 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_157
timestamp 1688980957
transform 1 0 15548 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_187
timestamp 1688980957
transform 1 0 18308 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_195
timestamp 1688980957
transform 1 0 19044 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_207
timestamp 1688980957
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_211
timestamp 1688980957
transform 1 0 20516 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_214
timestamp 1688980957
transform 1 0 20792 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_218
timestamp 1688980957
transform 1 0 21160 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_236
timestamp 1688980957
transform 1 0 22816 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_240
timestamp 1688980957
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_246
timestamp 1688980957
transform 1 0 23736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_250
timestamp 1688980957
transform 1 0 24104 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_260
timestamp 1688980957
transform 1 0 25024 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_272
timestamp 1688980957
transform 1 0 26128 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_347
timestamp 1688980957
transform 1 0 33028 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_23
timestamp 1688980957
transform 1 0 3220 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_33
timestamp 1688980957
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_39
timestamp 1688980957
transform 1 0 4692 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_49
timestamp 1688980957
transform 1 0 5612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_80
timestamp 1688980957
transform 1 0 8464 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_91
timestamp 1688980957
transform 1 0 9476 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_114
timestamp 1688980957
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_126
timestamp 1688980957
transform 1 0 12696 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_132
timestamp 1688980957
transform 1 0 13248 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_136
timestamp 1688980957
transform 1 0 13616 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_145
timestamp 1688980957
transform 1 0 14444 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_166
timestamp 1688980957
transform 1 0 16376 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_172
timestamp 1688980957
transform 1 0 16928 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_180
timestamp 1688980957
transform 1 0 17664 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_204
timestamp 1688980957
transform 1 0 19872 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_208
timestamp 1688980957
transform 1 0 20240 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_232
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_270
timestamp 1688980957
transform 1 0 25944 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_282
timestamp 1688980957
transform 1 0 27048 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_294
timestamp 1688980957
transform 1 0 28152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1688980957
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_52
timestamp 1688980957
transform 1 0 5888 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_78
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_92
timestamp 1688980957
transform 1 0 9568 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_98
timestamp 1688980957
transform 1 0 10120 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_102
timestamp 1688980957
transform 1 0 10488 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_106
timestamp 1688980957
transform 1 0 10856 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_116
timestamp 1688980957
transform 1 0 11776 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_120
timestamp 1688980957
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_124
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_129
timestamp 1688980957
transform 1 0 12972 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_141
timestamp 1688980957
transform 1 0 14076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_153
timestamp 1688980957
transform 1 0 15180 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_176
timestamp 1688980957
transform 1 0 17296 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_183
timestamp 1688980957
transform 1 0 17940 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_187
timestamp 1688980957
transform 1 0 18308 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_199
timestamp 1688980957
transform 1 0 19412 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_203
timestamp 1688980957
transform 1 0 19780 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_206
timestamp 1688980957
transform 1 0 20056 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_218
timestamp 1688980957
transform 1 0 21160 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_238
timestamp 1688980957
transform 1 0 23000 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_242
timestamp 1688980957
transform 1 0 23368 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_246
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_252
timestamp 1688980957
transform 1 0 24288 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_264
timestamp 1688980957
transform 1 0 25392 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_276
timestamp 1688980957
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_289
timestamp 1688980957
transform 1 0 27692 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_295
timestamp 1688980957
transform 1 0 28244 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_310
timestamp 1688980957
transform 1 0 29624 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_318
timestamp 1688980957
transform 1 0 30360 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_325
timestamp 1688980957
transform 1 0 31004 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_333
timestamp 1688980957
transform 1 0 31740 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_367
timestamp 1688980957
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_6
timestamp 1688980957
transform 1 0 1656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_18
timestamp 1688980957
transform 1 0 2760 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_22
timestamp 1688980957
transform 1 0 3128 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_33
timestamp 1688980957
transform 1 0 4140 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_45
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_57
timestamp 1688980957
transform 1 0 6348 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_69
timestamp 1688980957
transform 1 0 7452 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_79
timestamp 1688980957
transform 1 0 8372 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_98
timestamp 1688980957
transform 1 0 10120 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_122
timestamp 1688980957
transform 1 0 12328 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_148
timestamp 1688980957
transform 1 0 14720 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_160
timestamp 1688980957
transform 1 0 15824 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_164
timestamp 1688980957
transform 1 0 16192 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_170
timestamp 1688980957
transform 1 0 16744 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_190
timestamp 1688980957
transform 1 0 18584 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_205
timestamp 1688980957
transform 1 0 19964 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_213
timestamp 1688980957
transform 1 0 20700 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_217
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_225
timestamp 1688980957
transform 1 0 21804 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_231
timestamp 1688980957
transform 1 0 22356 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_235
timestamp 1688980957
transform 1 0 22724 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_240
timestamp 1688980957
transform 1 0 23184 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_244
timestamp 1688980957
transform 1 0 23552 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_290
timestamp 1688980957
transform 1 0 27784 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_332
timestamp 1688980957
transform 1 0 31648 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_344
timestamp 1688980957
transform 1 0 32752 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_348
timestamp 1688980957
transform 1 0 33120 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_356
timestamp 1688980957
transform 1 0 33856 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_362
timestamp 1688980957
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_73
timestamp 1688980957
transform 1 0 7820 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_117
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_121
timestamp 1688980957
transform 1 0 12236 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_135
timestamp 1688980957
transform 1 0 13524 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_139
timestamp 1688980957
transform 1 0 13892 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_151
timestamp 1688980957
transform 1 0 14996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_157
timestamp 1688980957
transform 1 0 15548 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_163
timestamp 1688980957
transform 1 0 16100 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_214
timestamp 1688980957
transform 1 0 20792 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_229
timestamp 1688980957
transform 1 0 22172 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_233
timestamp 1688980957
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_259
timestamp 1688980957
transform 1 0 24932 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_270
timestamp 1688980957
transform 1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_278
timestamp 1688980957
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_309
timestamp 1688980957
transform 1 0 29532 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_312
timestamp 1688980957
transform 1 0 29808 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_324
timestamp 1688980957
transform 1 0 30912 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_347
timestamp 1688980957
transform 1 0 33028 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_80
timestamp 1688980957
transform 1 0 8464 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_93
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_103
timestamp 1688980957
transform 1 0 10580 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_126
timestamp 1688980957
transform 1 0 12696 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1688980957
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_145
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_149
timestamp 1688980957
transform 1 0 14812 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_171
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_183
timestamp 1688980957
transform 1 0 17940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_207
timestamp 1688980957
transform 1 0 20148 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_211
timestamp 1688980957
transform 1 0 20516 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_215
timestamp 1688980957
transform 1 0 20884 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_231
timestamp 1688980957
transform 1 0 22356 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_235
timestamp 1688980957
transform 1 0 22724 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_272
timestamp 1688980957
transform 1 0 26128 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_284
timestamp 1688980957
transform 1 0 27232 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_291
timestamp 1688980957
transform 1 0 27876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_303
timestamp 1688980957
transform 1 0 28980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_322
timestamp 1688980957
transform 1 0 30728 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_338
timestamp 1688980957
transform 1 0 32200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_346
timestamp 1688980957
transform 1 0 32936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_83
timestamp 1688980957
transform 1 0 8740 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_87
timestamp 1688980957
transform 1 0 9108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_91
timestamp 1688980957
transform 1 0 9476 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_95
timestamp 1688980957
transform 1 0 9844 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_99
timestamp 1688980957
transform 1 0 10212 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_102
timestamp 1688980957
transform 1 0 10488 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_130
timestamp 1688980957
transform 1 0 13064 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_142
timestamp 1688980957
transform 1 0 14168 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_146
timestamp 1688980957
transform 1 0 14536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_176
timestamp 1688980957
transform 1 0 17296 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_180
timestamp 1688980957
transform 1 0 17664 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_188
timestamp 1688980957
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_192
timestamp 1688980957
transform 1 0 18768 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_204
timestamp 1688980957
transform 1 0 19872 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_210
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_213
timestamp 1688980957
transform 1 0 20700 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_229
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_232
timestamp 1688980957
transform 1 0 22448 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_236
timestamp 1688980957
transform 1 0 22816 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_240
timestamp 1688980957
transform 1 0 23184 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_244
timestamp 1688980957
transform 1 0 23552 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_248
timestamp 1688980957
transform 1 0 23920 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_260
timestamp 1688980957
transform 1 0 25024 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_272
timestamp 1688980957
transform 1 0 26128 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_295
timestamp 1688980957
transform 1 0 28244 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_344
timestamp 1688980957
transform 1 0 32752 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_356
timestamp 1688980957
transform 1 0 33856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_362
timestamp 1688980957
transform 1 0 34408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_365
timestamp 1688980957
transform 1 0 34684 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_6
timestamp 1688980957
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_18
timestamp 1688980957
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_105
timestamp 1688980957
transform 1 0 10764 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_117
timestamp 1688980957
transform 1 0 11868 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_125
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_170
timestamp 1688980957
transform 1 0 16744 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_187
timestamp 1688980957
transform 1 0 18308 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_206
timestamp 1688980957
transform 1 0 20056 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_214
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_218
timestamp 1688980957
transform 1 0 21160 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_222
timestamp 1688980957
transform 1 0 21528 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_226
timestamp 1688980957
transform 1 0 21896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_234
timestamp 1688980957
transform 1 0 22632 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_248
timestamp 1688980957
transform 1 0 23920 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_274
timestamp 1688980957
transform 1 0 26312 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_286
timestamp 1688980957
transform 1 0 27416 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_298
timestamp 1688980957
transform 1 0 28520 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_306
timestamp 1688980957
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_327
timestamp 1688980957
transform 1 0 31188 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_330
timestamp 1688980957
transform 1 0 31464 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_136
timestamp 1688980957
transform 1 0 13616 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_148
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_156
timestamp 1688980957
transform 1 0 15456 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_160
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_163
timestamp 1688980957
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_183
timestamp 1688980957
transform 1 0 17940 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_191
timestamp 1688980957
transform 1 0 18676 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_208
timestamp 1688980957
transform 1 0 20240 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_241
timestamp 1688980957
transform 1 0 23276 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_245
timestamp 1688980957
transform 1 0 23644 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_284
timestamp 1688980957
transform 1 0 27232 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_296
timestamp 1688980957
transform 1 0 28336 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_333
timestamp 1688980957
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_340
timestamp 1688980957
transform 1 0 32384 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_344
timestamp 1688980957
transform 1 0 32752 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_211
timestamp 1688980957
transform 1 0 20516 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_223
timestamp 1688980957
transform 1 0 21620 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_227
timestamp 1688980957
transform 1 0 21988 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_235
timestamp 1688980957
transform 1 0 22724 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_247
timestamp 1688980957
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_263
timestamp 1688980957
transform 1 0 25300 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_278
timestamp 1688980957
transform 1 0 26680 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_297
timestamp 1688980957
transform 1 0 28428 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_341
timestamp 1688980957
transform 1 0 32476 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_313
timestamp 1688980957
transform 1 0 29900 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_319
timestamp 1688980957
transform 1 0 30452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_331
timestamp 1688980957
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_341
timestamp 1688980957
transform 1 0 32476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_353
timestamp 1688980957
transform 1 0 33580 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_365
timestamp 1688980957
transform 1 0 34684 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_6
timestamp 1688980957
transform 1 0 1656 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_18
timestamp 1688980957
transform 1 0 2760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_241
timestamp 1688980957
transform 1 0 23276 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_272
timestamp 1688980957
transform 1 0 26128 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_300
timestamp 1688980957
transform 1 0 28704 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_346
timestamp 1688980957
transform 1 0 32936 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_262
timestamp 1688980957
transform 1 0 25208 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_268
timestamp 1688980957
transform 1 0 25760 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_309
timestamp 1688980957
transform 1 0 29532 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_320
timestamp 1688980957
transform 1 0 30544 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_332
timestamp 1688980957
transform 1 0 31648 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_341
timestamp 1688980957
transform 1 0 32476 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_344
timestamp 1688980957
transform 1 0 32752 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_257
timestamp 1688980957
transform 1 0 24748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_296
timestamp 1688980957
transform 1 0 28336 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_302
timestamp 1688980957
transform 1 0 28888 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_329
timestamp 1688980957
transform 1 0 31372 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_342
timestamp 1688980957
transform 1 0 32568 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_318
timestamp 1688980957
transform 1 0 30360 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_333
timestamp 1688980957
transform 1 0 31740 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_357
timestamp 1688980957
transform 1 0 33948 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_362
timestamp 1688980957
transform 1 0 34408 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_366
timestamp 1688980957
transform 1 0 34776 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_6
timestamp 1688980957
transform 1 0 1656 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_18
timestamp 1688980957
transform 1 0 2760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_341
timestamp 1688980957
transform 1 0 32476 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_348
timestamp 1688980957
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_360
timestamp 1688980957
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_367
timestamp 1688980957
transform 1 0 34868 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_367
timestamp 1688980957
transform 1 0 34868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_6
timestamp 1688980957
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_18
timestamp 1688980957
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_26
timestamp 1688980957
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_367
timestamp 1688980957
transform 1 0 34868 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_367
timestamp 1688980957
transform 1 0 34868 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_6
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_18
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_367
timestamp 1688980957
transform 1 0 34868 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_6
timestamp 1688980957
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1688980957
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_69
timestamp 1688980957
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_81
timestamp 1688980957
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_113
timestamp 1688980957
transform 1 0 11500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_125
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_169
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_181
timestamp 1688980957
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_237
timestamp 1688980957
transform 1 0 22908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_249
timestamp 1688980957
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_281
timestamp 1688980957
transform 1 0 26956 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_293
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_305
timestamp 1688980957
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_337
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1688980957
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 1656 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap8
timestamp 1688980957
transform 1 0 17940 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  max_cap48
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  max_cap49
timestamp 1688980957
transform -1 0 32476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output20
timestamp 1688980957
transform 1 0 33120 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 1688980957
transform -1 0 34592 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 1688980957
transform -1 0 34960 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 1688980957
transform -1 0 34592 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 1688980957
transform -1 0 34592 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 1688980957
transform -1 0 34592 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 1688980957
transform 1 0 33120 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 1688980957
transform 1 0 33120 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 1688980957
transform -1 0 34592 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 1688980957
transform -1 0 34592 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 1688980957
transform -1 0 34592 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 1688980957
transform -1 0 34592 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 1688980957
transform -1 0 34592 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 1688980957
transform -1 0 34960 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 1688980957
transform -1 0 34592 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output35
timestamp 1688980957
transform -1 0 34592 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 35236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 35236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 35236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 35236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 35236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 35236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 35236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 35236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 35236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 35236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 35236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 35236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 35236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 35236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 35236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 35236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 35236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 35236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 35236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 35236 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 35236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 35236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 35236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 35236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 35236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 35236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 35236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 35236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 35236 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 35236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 35236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 35236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 35236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 35236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 35236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 35236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 35236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 35236 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 35236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 35236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 35236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 35236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 35236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 35236 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 35236 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 35236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 35236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 35236 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 11408 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 21712 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 32016 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire1
timestamp 1688980957
transform -1 0 24288 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire2
timestamp 1688980957
transform 1 0 25392 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire3
timestamp 1688980957
transform -1 0 25024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire4
timestamp 1688980957
transform 1 0 25668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire5
timestamp 1688980957
transform -1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire6
timestamp 1688980957
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire7
timestamp 1688980957
transform -1 0 25484 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire9
timestamp 1688980957
transform -1 0 18492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire36
timestamp 1688980957
transform 1 0 26496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire37
timestamp 1688980957
transform -1 0 26036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire38
timestamp 1688980957
transform -1 0 25760 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire39
timestamp 1688980957
transform -1 0 25208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire40
timestamp 1688980957
transform 1 0 26312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire41
timestamp 1688980957
transform -1 0 26312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire42
timestamp 1688980957
transform -1 0 26036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire43
timestamp 1688980957
transform -1 0 25760 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire44
timestamp 1688980957
transform -1 0 25208 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire45
timestamp 1688980957
transform -1 0 24932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire46
timestamp 1688980957
transform 1 0 25944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  wire47
timestamp 1688980957
transform -1 0 24748 0 1 11968
box -38 -48 314 592
<< labels >>
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 a[0]
port 0 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 a[1]
port 1 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 a[2]
port 2 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 a[3]
port 3 nsew signal input
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 a[4]
port 4 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 a[5]
port 5 nsew signal input
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 a[6]
port 6 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 a[7]
port 7 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 b[0]
port 8 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 b[1]
port 9 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 b[2]
port 10 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 b[3]
port 11 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 b[4]
port 12 nsew signal input
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 b[5]
port 13 nsew signal input
flabel metal3 s 0 32376 800 32496 0 FreeSans 480 0 0 0 b[6]
port 14 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 b[7]
port 15 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 control
port 17 nsew signal input
flabel metal3 s 35600 3000 36400 3120 0 FreeSans 480 0 0 0 p[0]
port 18 nsew signal tristate
flabel metal3 s 35600 24760 36400 24880 0 FreeSans 480 0 0 0 p[10]
port 19 nsew signal tristate
flabel metal3 s 35600 26936 36400 27056 0 FreeSans 480 0 0 0 p[11]
port 20 nsew signal tristate
flabel metal3 s 35600 29112 36400 29232 0 FreeSans 480 0 0 0 p[12]
port 21 nsew signal tristate
flabel metal3 s 35600 31288 36400 31408 0 FreeSans 480 0 0 0 p[13]
port 22 nsew signal tristate
flabel metal3 s 35600 33464 36400 33584 0 FreeSans 480 0 0 0 p[14]
port 23 nsew signal tristate
flabel metal3 s 35600 35640 36400 35760 0 FreeSans 480 0 0 0 p[15]
port 24 nsew signal tristate
flabel metal3 s 35600 5176 36400 5296 0 FreeSans 480 0 0 0 p[1]
port 25 nsew signal tristate
flabel metal3 s 35600 7352 36400 7472 0 FreeSans 480 0 0 0 p[2]
port 26 nsew signal tristate
flabel metal3 s 35600 9528 36400 9648 0 FreeSans 480 0 0 0 p[3]
port 27 nsew signal tristate
flabel metal3 s 35600 11704 36400 11824 0 FreeSans 480 0 0 0 p[4]
port 28 nsew signal tristate
flabel metal3 s 35600 13880 36400 14000 0 FreeSans 480 0 0 0 p[5]
port 29 nsew signal tristate
flabel metal3 s 35600 16056 36400 16176 0 FreeSans 480 0 0 0 p[6]
port 30 nsew signal tristate
flabel metal3 s 35600 18232 36400 18352 0 FreeSans 480 0 0 0 p[7]
port 31 nsew signal tristate
flabel metal3 s 35600 20408 36400 20528 0 FreeSans 480 0 0 0 p[8]
port 32 nsew signal tristate
flabel metal3 s 35600 22584 36400 22704 0 FreeSans 480 0 0 0 p[9]
port 33 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 rst
port 34 nsew signal input
flabel metal4 s 4208 2128 4528 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 34928 2128 35248 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 19568 2128 19888 36496 0 FreeSans 1920 90 0 0 vssd1
port 36 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36400 38800
<< end >>
