VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vmsu_8bit_top
  CLASS BLOCK ;
  FOREIGN vmsu_8bit_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 182.000 BY 194.000 ;
  PIN a[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END a[0]
  PIN a[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.200 4.000 42.800 ;
    END
  END a[1]
  PIN a[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END a[2]
  PIN a[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END a[3]
  PIN a[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END a[4]
  PIN a[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END a[5]
  PIN a[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END a[6]
  PIN a[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END a[7]
  PIN b[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END b[0]
  PIN b[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.080 4.000 53.680 ;
    END
  END b[1]
  PIN b[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END b[2]
  PIN b[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END b[3]
  PIN b[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 118.360 4.000 118.960 ;
    END
  END b[4]
  PIN b[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END b[5]
  PIN b[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END b[6]
  PIN b[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END b[7]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END clk
  PIN control
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END control
  PIN p[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 15.000 182.000 15.600 ;
    END
  END p[0]
  PIN p[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 123.800 182.000 124.400 ;
    END
  END p[10]
  PIN p[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 134.680 182.000 135.280 ;
    END
  END p[11]
  PIN p[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 145.560 182.000 146.160 ;
    END
  END p[12]
  PIN p[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 156.440 182.000 157.040 ;
    END
  END p[13]
  PIN p[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 167.320 182.000 167.920 ;
    END
  END p[14]
  PIN p[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 178.200 182.000 178.800 ;
    END
  END p[15]
  PIN p[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 25.880 182.000 26.480 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 36.760 182.000 37.360 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 47.640 182.000 48.240 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 58.520 182.000 59.120 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 69.400 182.000 70.000 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 80.280 182.000 80.880 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 91.160 182.000 91.760 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 102.040 182.000 102.640 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 178.000 112.920 182.000 113.520 ;
    END
  END p[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 182.480 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 182.480 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 182.480 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 176.180 182.325 ;
      LAYER met1 ;
        RECT 4.670 10.640 176.480 182.480 ;
      LAYER met2 ;
        RECT 4.690 4.280 176.210 184.125 ;
        RECT 4.690 4.000 44.890 4.280 ;
        RECT 45.730 4.000 135.970 4.280 ;
        RECT 136.810 4.000 176.210 4.280 ;
      LAYER met3 ;
        RECT 4.400 183.240 178.000 184.105 ;
        RECT 3.990 179.200 178.000 183.240 ;
        RECT 3.990 177.800 177.600 179.200 ;
        RECT 3.990 173.760 178.000 177.800 ;
        RECT 4.400 172.360 178.000 173.760 ;
        RECT 3.990 168.320 178.000 172.360 ;
        RECT 3.990 166.920 177.600 168.320 ;
        RECT 3.990 162.880 178.000 166.920 ;
        RECT 4.400 161.480 178.000 162.880 ;
        RECT 3.990 157.440 178.000 161.480 ;
        RECT 3.990 156.040 177.600 157.440 ;
        RECT 3.990 152.000 178.000 156.040 ;
        RECT 4.400 150.600 178.000 152.000 ;
        RECT 3.990 146.560 178.000 150.600 ;
        RECT 3.990 145.160 177.600 146.560 ;
        RECT 3.990 141.120 178.000 145.160 ;
        RECT 4.400 139.720 178.000 141.120 ;
        RECT 3.990 135.680 178.000 139.720 ;
        RECT 3.990 134.280 177.600 135.680 ;
        RECT 3.990 130.240 178.000 134.280 ;
        RECT 4.400 128.840 178.000 130.240 ;
        RECT 3.990 124.800 178.000 128.840 ;
        RECT 3.990 123.400 177.600 124.800 ;
        RECT 3.990 119.360 178.000 123.400 ;
        RECT 4.400 117.960 178.000 119.360 ;
        RECT 3.990 113.920 178.000 117.960 ;
        RECT 3.990 112.520 177.600 113.920 ;
        RECT 3.990 108.480 178.000 112.520 ;
        RECT 4.400 107.080 178.000 108.480 ;
        RECT 3.990 103.040 178.000 107.080 ;
        RECT 3.990 101.640 177.600 103.040 ;
        RECT 3.990 97.600 178.000 101.640 ;
        RECT 4.400 96.200 178.000 97.600 ;
        RECT 3.990 92.160 178.000 96.200 ;
        RECT 3.990 90.760 177.600 92.160 ;
        RECT 3.990 86.720 178.000 90.760 ;
        RECT 4.400 85.320 178.000 86.720 ;
        RECT 3.990 81.280 178.000 85.320 ;
        RECT 3.990 79.880 177.600 81.280 ;
        RECT 3.990 75.840 178.000 79.880 ;
        RECT 4.400 74.440 178.000 75.840 ;
        RECT 3.990 70.400 178.000 74.440 ;
        RECT 3.990 69.000 177.600 70.400 ;
        RECT 3.990 64.960 178.000 69.000 ;
        RECT 4.400 63.560 178.000 64.960 ;
        RECT 3.990 59.520 178.000 63.560 ;
        RECT 3.990 58.120 177.600 59.520 ;
        RECT 3.990 54.080 178.000 58.120 ;
        RECT 4.400 52.680 178.000 54.080 ;
        RECT 3.990 48.640 178.000 52.680 ;
        RECT 3.990 47.240 177.600 48.640 ;
        RECT 3.990 43.200 178.000 47.240 ;
        RECT 4.400 41.800 178.000 43.200 ;
        RECT 3.990 37.760 178.000 41.800 ;
        RECT 3.990 36.360 177.600 37.760 ;
        RECT 3.990 32.320 178.000 36.360 ;
        RECT 4.400 30.920 178.000 32.320 ;
        RECT 3.990 26.880 178.000 30.920 ;
        RECT 3.990 25.480 177.600 26.880 ;
        RECT 3.990 21.440 178.000 25.480 ;
        RECT 4.400 20.040 178.000 21.440 ;
        RECT 3.990 16.000 178.000 20.040 ;
        RECT 3.990 14.600 177.600 16.000 ;
        RECT 3.990 10.560 178.000 14.600 ;
        RECT 4.400 9.695 178.000 10.560 ;
  END
END vmsu_8bit_top
END LIBRARY

