magic
tech sky130A
magscale 1 2
timestamp 1726899427
<< viali >>
rect 18245 19329 18279 19363
rect 18153 19261 18187 19295
rect 18521 19125 18555 19159
rect 13277 18785 13311 18819
rect 16405 18785 16439 18819
rect 18061 18785 18095 18819
rect 19901 18785 19935 18819
rect 12633 18717 12667 18751
rect 12725 18717 12759 18751
rect 16497 18717 16531 18751
rect 18245 18717 18279 18751
rect 19993 18717 20027 18751
rect 20637 18717 20671 18751
rect 20913 18717 20947 18751
rect 21373 18717 21407 18751
rect 20453 18649 20487 18683
rect 21005 18649 21039 18683
rect 21189 18649 21223 18683
rect 16865 18581 16899 18615
rect 18429 18581 18463 18615
rect 20361 18581 20395 18615
rect 20821 18581 20855 18615
rect 20361 18377 20395 18411
rect 12633 18309 12667 18343
rect 15577 18309 15611 18343
rect 18429 18309 18463 18343
rect 12909 18241 12943 18275
rect 14565 18241 14599 18275
rect 15669 18241 15703 18275
rect 15761 18241 15795 18275
rect 15945 18241 15979 18275
rect 18613 18241 18647 18275
rect 18705 18241 18739 18275
rect 19993 18241 20027 18275
rect 20177 18241 20211 18275
rect 20637 18241 20671 18275
rect 20913 18241 20947 18275
rect 11805 18173 11839 18207
rect 12725 18173 12759 18207
rect 21649 18173 21683 18207
rect 13093 18037 13127 18071
rect 15945 18037 15979 18071
rect 18429 18037 18463 18071
rect 14841 17833 14875 17867
rect 15945 17833 15979 17867
rect 16313 17833 16347 17867
rect 19809 17833 19843 17867
rect 10793 17697 10827 17731
rect 13093 17697 13127 17731
rect 15025 17697 15059 17731
rect 15485 17697 15519 17731
rect 16681 17697 16715 17731
rect 16773 17697 16807 17731
rect 16957 17697 16991 17731
rect 17693 17697 17727 17731
rect 18061 17697 18095 17731
rect 18889 17697 18923 17731
rect 10333 17629 10367 17663
rect 10609 17629 10643 17663
rect 10885 17629 10919 17663
rect 11345 17629 11379 17663
rect 11529 17629 11563 17663
rect 12081 17629 12115 17663
rect 12357 17629 12391 17663
rect 12541 17629 12575 17663
rect 13185 17629 13219 17663
rect 13461 17629 13495 17663
rect 13737 17629 13771 17663
rect 15117 17629 15151 17663
rect 15761 17629 15795 17663
rect 16037 17629 16071 17663
rect 16497 17629 16531 17663
rect 16589 17629 16623 17663
rect 17049 17629 17083 17663
rect 17325 17629 17359 17663
rect 17509 17629 17543 17663
rect 18153 17629 18187 17663
rect 18429 17629 18463 17663
rect 18797 17629 18831 17663
rect 19349 17629 19383 17663
rect 19441 17629 19475 17663
rect 19809 17629 19843 17663
rect 11437 17561 11471 17595
rect 12173 17561 12207 17595
rect 12725 17561 12759 17595
rect 13553 17561 13587 17595
rect 13921 17561 13955 17595
rect 18521 17561 18555 17595
rect 10425 17493 10459 17527
rect 13369 17493 13403 17527
rect 17141 17493 17175 17527
rect 18337 17493 18371 17527
rect 19073 17493 19107 17527
rect 19993 17493 20027 17527
rect 10517 17289 10551 17323
rect 15593 17289 15627 17323
rect 15761 17289 15795 17323
rect 18721 17289 18755 17323
rect 18889 17289 18923 17323
rect 10701 17221 10735 17255
rect 12265 17221 12299 17255
rect 15393 17221 15427 17255
rect 17141 17221 17175 17255
rect 17233 17221 17267 17255
rect 18521 17221 18555 17255
rect 20637 17221 20671 17255
rect 21833 17221 21867 17255
rect 9873 17153 9907 17187
rect 10609 17153 10643 17187
rect 10793 17153 10827 17187
rect 12449 17153 12483 17187
rect 12541 17153 12575 17187
rect 13001 17153 13035 17187
rect 13185 17153 13219 17187
rect 13277 17153 13311 17187
rect 16221 17153 16255 17187
rect 16405 17153 16439 17187
rect 16773 17153 16807 17187
rect 16865 17153 16899 17187
rect 16957 17153 16991 17187
rect 17417 17153 17451 17187
rect 17509 17153 17543 17187
rect 20821 17153 20855 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 21097 17153 21131 17187
rect 21281 17153 21315 17187
rect 22385 17153 22419 17187
rect 9689 17085 9723 17119
rect 22477 17085 22511 17119
rect 12541 17017 12575 17051
rect 13277 17017 13311 17051
rect 22109 17017 22143 17051
rect 15577 16949 15611 16983
rect 16405 16949 16439 16983
rect 17509 16949 17543 16983
rect 18705 16949 18739 16983
rect 20913 16949 20947 16983
rect 21465 16949 21499 16983
rect 9689 16745 9723 16779
rect 14841 16745 14875 16779
rect 9505 16677 9539 16711
rect 9229 16609 9263 16643
rect 9597 16609 9631 16643
rect 9781 16609 9815 16643
rect 10057 16609 10091 16643
rect 16865 16609 16899 16643
rect 17785 16609 17819 16643
rect 22661 16609 22695 16643
rect 9137 16541 9171 16575
rect 9873 16541 9907 16575
rect 9965 16541 9999 16575
rect 10149 16541 10183 16575
rect 14565 16541 14599 16575
rect 14933 16541 14967 16575
rect 15117 16541 15151 16575
rect 15301 16541 15335 16575
rect 16957 16541 16991 16575
rect 21005 16541 21039 16575
rect 22109 16541 22143 16575
rect 22477 16541 22511 16575
rect 22017 16473 22051 16507
rect 14657 16405 14691 16439
rect 14749 16405 14783 16439
rect 15301 16405 15335 16439
rect 22477 16405 22511 16439
rect 11345 16201 11379 16235
rect 14289 16201 14323 16235
rect 14657 16201 14691 16235
rect 19349 16201 19383 16235
rect 21373 16201 21407 16235
rect 24133 16201 24167 16235
rect 10793 16133 10827 16167
rect 11161 16133 11195 16167
rect 13737 16133 13771 16167
rect 15025 16133 15059 16167
rect 15301 16133 15335 16167
rect 15393 16133 15427 16167
rect 15761 16133 15795 16167
rect 21097 16133 21131 16167
rect 26065 16133 26099 16167
rect 10425 16065 10459 16099
rect 10977 16065 11011 16099
rect 15117 16065 15151 16099
rect 15485 16065 15519 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 17969 16065 18003 16099
rect 18521 16065 18555 16099
rect 19809 16065 19843 16099
rect 20269 16065 20303 16099
rect 20545 16065 20579 16099
rect 20637 16065 20671 16099
rect 20729 16065 20763 16099
rect 20913 16065 20947 16099
rect 21005 16065 21039 16099
rect 21189 16065 21223 16099
rect 21281 16065 21315 16099
rect 21465 16065 21499 16099
rect 22201 16065 22235 16099
rect 23305 16065 23339 16099
rect 23765 16065 23799 16099
rect 23858 16065 23892 16099
rect 24685 16065 24719 16099
rect 27077 16065 27111 16099
rect 28181 16065 28215 16099
rect 28365 16065 28399 16099
rect 10241 15997 10275 16031
rect 12909 15997 12943 16031
rect 13829 15997 13863 16031
rect 14381 15997 14415 16031
rect 14473 15997 14507 16031
rect 14749 15997 14783 16031
rect 14841 15997 14875 16031
rect 17417 15997 17451 16031
rect 18061 15997 18095 16031
rect 18429 15997 18463 16031
rect 19717 15997 19751 16031
rect 20085 15997 20119 16031
rect 20821 15997 20855 16031
rect 22109 15997 22143 16031
rect 23397 15997 23431 16031
rect 25697 15997 25731 16031
rect 28089 15997 28123 16031
rect 14197 15929 14231 15963
rect 15669 15929 15703 15963
rect 17693 15929 17727 15963
rect 23673 15929 23707 15963
rect 26341 15929 26375 15963
rect 10701 15861 10735 15895
rect 19441 15861 19475 15895
rect 22569 15861 22603 15895
rect 26525 15861 26559 15895
rect 28181 15861 28215 15895
rect 9689 15657 9723 15691
rect 10885 15657 10919 15691
rect 11437 15657 11471 15691
rect 15301 15657 15335 15691
rect 21557 15657 21591 15691
rect 27721 15657 27755 15691
rect 10701 15589 10735 15623
rect 13369 15589 13403 15623
rect 27169 15589 27203 15623
rect 27261 15589 27295 15623
rect 12173 15521 12207 15555
rect 12817 15521 12851 15555
rect 13737 15521 13771 15555
rect 16405 15521 16439 15555
rect 17785 15521 17819 15555
rect 25697 15521 25731 15555
rect 26525 15521 26559 15555
rect 27629 15521 27663 15555
rect 9413 15453 9447 15487
rect 9689 15453 9723 15487
rect 11161 15453 11195 15487
rect 11989 15453 12023 15487
rect 14749 15453 14783 15487
rect 15117 15453 15151 15487
rect 15945 15453 15979 15487
rect 16037 15453 16071 15487
rect 16221 15453 16255 15487
rect 16773 15453 16807 15487
rect 16957 15453 16991 15487
rect 21097 15453 21131 15487
rect 21189 15453 21223 15487
rect 21373 15453 21407 15487
rect 24961 15453 24995 15487
rect 25145 15453 25179 15487
rect 27077 15453 27111 15487
rect 27353 15453 27387 15487
rect 27905 15453 27939 15487
rect 11069 15385 11103 15419
rect 11253 15385 11287 15419
rect 11437 15385 11471 15419
rect 14933 15385 14967 15419
rect 15025 15385 15059 15419
rect 27537 15385 27571 15419
rect 9505 15317 9539 15351
rect 10885 15317 10919 15351
rect 13093 15317 13127 15351
rect 13277 15317 13311 15351
rect 25053 15317 25087 15351
rect 26893 15317 26927 15351
rect 27813 15317 27847 15351
rect 9321 15113 9355 15147
rect 9689 15113 9723 15147
rect 10241 15113 10275 15147
rect 10609 15113 10643 15147
rect 17141 15113 17175 15147
rect 17233 15113 17267 15147
rect 9413 15045 9447 15079
rect 9873 15045 9907 15079
rect 10333 15045 10367 15079
rect 10517 15045 10551 15079
rect 12633 15045 12667 15079
rect 21373 15045 21407 15079
rect 9505 14977 9539 15011
rect 9784 14999 9818 15033
rect 10057 14977 10091 15011
rect 10609 14977 10643 15011
rect 11989 14977 12023 15011
rect 12173 14977 12207 15011
rect 12265 14977 12299 15011
rect 12357 14977 12391 15011
rect 13093 14977 13127 15011
rect 13277 14977 13311 15011
rect 16957 14977 16991 15011
rect 17509 14977 17543 15011
rect 17601 14977 17635 15011
rect 17969 14977 18003 15011
rect 19625 14977 19659 15011
rect 21189 14977 21223 15011
rect 21465 14977 21499 15011
rect 9137 14909 9171 14943
rect 16773 14909 16807 14943
rect 17693 14909 17727 14943
rect 19533 14909 19567 14943
rect 13093 14841 13127 14875
rect 19993 14841 20027 14875
rect 17785 14773 17819 14807
rect 21465 14773 21499 14807
rect 9689 14569 9723 14603
rect 10057 14569 10091 14603
rect 12173 14569 12207 14603
rect 15117 14569 15151 14603
rect 15577 14569 15611 14603
rect 16313 14569 16347 14603
rect 17509 14569 17543 14603
rect 17877 14569 17911 14603
rect 18245 14569 18279 14603
rect 22109 14569 22143 14603
rect 23673 14569 23707 14603
rect 24409 14569 24443 14603
rect 12357 14501 12391 14535
rect 21833 14501 21867 14535
rect 24041 14501 24075 14535
rect 24777 14501 24811 14535
rect 10149 14433 10183 14467
rect 13001 14433 13035 14467
rect 13185 14433 13219 14467
rect 17785 14433 17819 14467
rect 23765 14433 23799 14467
rect 25789 14433 25823 14467
rect 9137 14365 9171 14399
rect 9505 14365 9539 14399
rect 9781 14365 9815 14399
rect 9873 14365 9907 14399
rect 11529 14365 11563 14399
rect 11713 14365 11747 14399
rect 11805 14365 11839 14399
rect 11897 14365 11931 14399
rect 12357 14365 12391 14399
rect 12541 14365 12575 14399
rect 12909 14365 12943 14399
rect 13277 14365 13311 14399
rect 13553 14365 13587 14399
rect 14105 14365 14139 14399
rect 14289 14365 14323 14399
rect 14381 14365 14415 14399
rect 14473 14365 14507 14399
rect 15301 14365 15335 14399
rect 15393 14365 15427 14399
rect 15669 14365 15703 14399
rect 15853 14365 15887 14399
rect 15945 14365 15979 14399
rect 16037 14365 16071 14399
rect 17693 14365 17727 14399
rect 18061 14365 18095 14399
rect 18245 14365 18279 14399
rect 21373 14365 21407 14399
rect 21649 14365 21683 14399
rect 23489 14365 23523 14399
rect 24409 14365 24443 14399
rect 24501 14365 24535 14399
rect 24961 14365 24995 14399
rect 25145 14365 25179 14399
rect 25605 14365 25639 14399
rect 25881 14365 25915 14399
rect 26065 14365 26099 14399
rect 9321 14297 9355 14331
rect 9413 14297 9447 14331
rect 15577 14297 15611 14331
rect 17969 14297 18003 14331
rect 21465 14297 21499 14331
rect 21951 14297 21985 14331
rect 22125 14297 22159 14331
rect 25329 14297 25363 14331
rect 9965 14229 9999 14263
rect 11069 14229 11103 14263
rect 11345 14229 11379 14263
rect 13829 14229 13863 14263
rect 14749 14229 14783 14263
rect 22293 14229 22327 14263
rect 23305 14229 23339 14263
rect 25421 14229 25455 14263
rect 25881 14229 25915 14263
rect 9413 14025 9447 14059
rect 10241 14025 10275 14059
rect 12173 14025 12207 14059
rect 12725 14025 12759 14059
rect 13277 14025 13311 14059
rect 14473 14025 14507 14059
rect 15853 14025 15887 14059
rect 18705 14025 18739 14059
rect 19073 14025 19107 14059
rect 19717 14025 19751 14059
rect 20821 14025 20855 14059
rect 21925 14025 21959 14059
rect 22753 14025 22787 14059
rect 9965 13957 9999 13991
rect 12817 13957 12851 13991
rect 13829 13957 13863 13991
rect 15209 13957 15243 13991
rect 18429 13957 18463 13991
rect 22201 13957 22235 13991
rect 22385 13957 22419 13991
rect 24225 13957 24259 13991
rect 9689 13889 9723 13923
rect 10885 13889 10919 13923
rect 12541 13889 12575 13923
rect 14197 13889 14231 13923
rect 14841 13889 14875 13923
rect 14933 13889 14967 13923
rect 15025 13889 15059 13923
rect 15577 13889 15611 13923
rect 18705 13889 18739 13923
rect 18797 13889 18831 13923
rect 19349 13889 19383 13923
rect 19533 13889 19567 13923
rect 20729 13889 20763 13923
rect 21097 13889 21131 13923
rect 21373 13889 21407 13923
rect 21463 13889 21497 13923
rect 21649 13889 21683 13923
rect 21833 13889 21867 13923
rect 22017 13889 22051 13923
rect 22937 13889 22971 13923
rect 23029 13889 23063 13923
rect 23213 13889 23247 13923
rect 23305 13889 23339 13923
rect 23397 13889 23431 13923
rect 23581 13889 23615 13923
rect 23673 13889 23707 13923
rect 23765 13889 23799 13923
rect 24133 13889 24167 13923
rect 24317 13889 24351 13923
rect 24409 13889 24443 13923
rect 24593 13889 24627 13923
rect 24869 13889 24903 13923
rect 25145 13889 25179 13923
rect 25237 13889 25271 13923
rect 25421 13889 25455 13923
rect 25697 13889 25731 13923
rect 9597 13821 9631 13855
rect 10057 13821 10091 13855
rect 10517 13821 10551 13855
rect 12357 13821 12391 13855
rect 12909 13821 12943 13855
rect 13645 13821 13679 13855
rect 13921 13821 13955 13855
rect 14289 13821 14323 13855
rect 14565 13821 14599 13855
rect 14749 13821 14783 13855
rect 15301 13821 15335 13855
rect 15669 13821 15703 13855
rect 19073 13821 19107 13855
rect 19257 13821 19291 13855
rect 22569 13821 22603 13855
rect 25789 13821 25823 13855
rect 10609 13753 10643 13787
rect 18613 13753 18647 13787
rect 18889 13753 18923 13787
rect 26065 13753 26099 13787
rect 10747 13685 10781 13719
rect 21189 13685 21223 13719
rect 24041 13685 24075 13719
rect 24501 13685 24535 13719
rect 24777 13685 24811 13719
rect 25421 13685 25455 13719
rect 14933 13481 14967 13515
rect 15025 13481 15059 13515
rect 23213 13481 23247 13515
rect 23489 13481 23523 13515
rect 24593 13481 24627 13515
rect 25973 13481 26007 13515
rect 26985 13481 27019 13515
rect 14197 13413 14231 13447
rect 17049 13413 17083 13447
rect 17233 13413 17267 13447
rect 24961 13413 24995 13447
rect 27353 13413 27387 13447
rect 15577 13345 15611 13379
rect 16313 13345 16347 13379
rect 18613 13345 18647 13379
rect 19993 13345 20027 13379
rect 25513 13345 25547 13379
rect 26341 13345 26375 13379
rect 27077 13345 27111 13379
rect 9873 13277 9907 13311
rect 10057 13277 10091 13311
rect 15209 13277 15243 13311
rect 15301 13277 15335 13311
rect 16405 13277 16439 13311
rect 16681 13277 16715 13311
rect 17601 13277 17635 13311
rect 17785 13277 17819 13311
rect 18061 13277 18095 13311
rect 18521 13277 18555 13311
rect 19901 13277 19935 13311
rect 23029 13277 23063 13311
rect 23213 13277 23247 13311
rect 23305 13277 23339 13311
rect 23489 13277 23523 13311
rect 24869 13277 24903 13311
rect 25053 13277 25087 13311
rect 25605 13277 25639 13311
rect 25789 13277 25823 13311
rect 26249 13277 26283 13311
rect 26985 13277 27019 13311
rect 27445 13277 27479 13311
rect 27629 13277 27663 13311
rect 9689 13209 9723 13243
rect 14197 13209 14231 13243
rect 15393 13209 15427 13243
rect 16773 13209 16807 13243
rect 18245 13209 18279 13243
rect 18429 13209 18463 13243
rect 24409 13209 24443 13243
rect 24625 13209 24659 13243
rect 10333 13141 10367 13175
rect 10701 13141 10735 13175
rect 14657 13141 14691 13175
rect 14749 13141 14783 13175
rect 17693 13141 17727 13175
rect 20269 13141 20303 13175
rect 24041 13141 24075 13175
rect 24777 13141 24811 13175
rect 26617 13141 26651 13175
rect 27813 13141 27847 13175
rect 11161 12937 11195 12971
rect 15485 12937 15519 12971
rect 16681 12937 16715 12971
rect 19901 12937 19935 12971
rect 26801 12937 26835 12971
rect 9045 12869 9079 12903
rect 9245 12869 9279 12903
rect 9873 12869 9907 12903
rect 10977 12869 11011 12903
rect 15669 12869 15703 12903
rect 19441 12869 19475 12903
rect 21925 12869 21959 12903
rect 8769 12801 8803 12835
rect 8953 12801 8987 12835
rect 9689 12801 9723 12835
rect 10333 12801 10367 12835
rect 10885 12801 10919 12835
rect 11069 12801 11103 12835
rect 11161 12801 11195 12835
rect 11345 12801 11379 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 11989 12801 12023 12835
rect 12265 12801 12299 12835
rect 14657 12801 14691 12835
rect 15853 12801 15887 12835
rect 16037 12801 16071 12835
rect 17233 12801 17267 12835
rect 17417 12801 17451 12835
rect 18981 12801 19015 12835
rect 26525 12801 26559 12835
rect 27905 12801 27939 12835
rect 9505 12733 9539 12767
rect 9965 12733 9999 12767
rect 10425 12733 10459 12767
rect 12173 12733 12207 12767
rect 12541 12733 12575 12767
rect 15209 12733 15243 12767
rect 17049 12733 17083 12767
rect 26801 12733 26835 12767
rect 27813 12733 27847 12767
rect 11805 12665 11839 12699
rect 11897 12665 11931 12699
rect 15025 12665 15059 12699
rect 15117 12665 15151 12699
rect 17141 12665 17175 12699
rect 19717 12665 19751 12699
rect 22201 12665 22235 12699
rect 8953 12597 8987 12631
rect 9229 12597 9263 12631
rect 9413 12597 9447 12631
rect 12357 12597 12391 12631
rect 12817 12597 12851 12631
rect 16957 12597 16991 12631
rect 19073 12597 19107 12631
rect 22385 12597 22419 12631
rect 26617 12597 26651 12631
rect 28273 12597 28307 12631
rect 9321 12393 9355 12427
rect 11253 12393 11287 12427
rect 11713 12393 11747 12427
rect 12081 12393 12115 12427
rect 15025 12393 15059 12427
rect 15945 12393 15979 12427
rect 16405 12393 16439 12427
rect 16497 12393 16531 12427
rect 19257 12393 19291 12427
rect 22293 12393 22327 12427
rect 25789 12393 25823 12427
rect 26525 12393 26559 12427
rect 9689 12325 9723 12359
rect 9781 12325 9815 12359
rect 16865 12325 16899 12359
rect 28733 12325 28767 12359
rect 9597 12257 9631 12291
rect 16037 12257 16071 12291
rect 17233 12257 17267 12291
rect 18337 12257 18371 12291
rect 18981 12257 19015 12291
rect 22385 12257 22419 12291
rect 23857 12257 23891 12291
rect 25237 12257 25271 12291
rect 29101 12257 29135 12291
rect 10149 12189 10183 12223
rect 11069 12189 11103 12223
rect 11345 12189 11379 12223
rect 11529 12189 11563 12223
rect 11621 12189 11655 12223
rect 11805 12189 11839 12223
rect 13277 12189 13311 12223
rect 13461 12189 13495 12223
rect 14749 12189 14783 12223
rect 14841 12189 14875 12223
rect 16221 12189 16255 12223
rect 16681 12189 16715 12223
rect 16773 12189 16807 12223
rect 16957 12189 16991 12223
rect 17141 12189 17175 12223
rect 17417 12189 17451 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 18797 12189 18831 12223
rect 18889 12189 18923 12223
rect 19073 12189 19107 12223
rect 19533 12189 19567 12223
rect 22109 12189 22143 12223
rect 22661 12189 22695 12223
rect 23029 12189 23063 12223
rect 23765 12189 23799 12223
rect 23949 12189 23983 12223
rect 24593 12189 24627 12223
rect 24777 12189 24811 12223
rect 25053 12189 25087 12223
rect 25605 12189 25639 12223
rect 25789 12189 25823 12223
rect 26157 12189 26191 12223
rect 26341 12189 26375 12223
rect 27905 12189 27939 12223
rect 28181 12189 28215 12223
rect 28273 12189 28307 12223
rect 28457 12189 28491 12223
rect 28917 12189 28951 12223
rect 10885 12121 10919 12155
rect 14381 12121 14415 12155
rect 14473 12121 14507 12155
rect 15945 12121 15979 12155
rect 18429 12121 18463 12155
rect 18613 12121 18647 12155
rect 19257 12121 19291 12155
rect 28641 12121 28675 12155
rect 10701 12053 10735 12087
rect 13369 12053 13403 12087
rect 17601 12053 17635 12087
rect 19441 12053 19475 12087
rect 21925 12053 21959 12087
rect 23673 12053 23707 12087
rect 24409 12053 24443 12087
rect 24869 12053 24903 12087
rect 27721 12053 27755 12087
rect 28089 12053 28123 12087
rect 9321 11849 9355 11883
rect 11989 11849 12023 11883
rect 14473 11849 14507 11883
rect 18429 11849 18463 11883
rect 22385 11849 22419 11883
rect 26525 11849 26559 11883
rect 9597 11713 9631 11747
rect 9689 11713 9723 11747
rect 9781 11713 9815 11747
rect 9965 11713 9999 11747
rect 10425 11713 10459 11747
rect 11529 11713 11563 11747
rect 11805 11713 11839 11747
rect 12081 11713 12115 11747
rect 12265 11713 12299 11747
rect 12449 11713 12483 11747
rect 14197 11713 14231 11747
rect 15025 11713 15059 11747
rect 16681 11713 16715 11747
rect 16865 11713 16899 11747
rect 18337 11713 18371 11747
rect 18521 11713 18555 11747
rect 19257 11713 19291 11747
rect 19441 11713 19475 11747
rect 19993 11713 20027 11747
rect 20453 11713 20487 11747
rect 22017 11713 22051 11747
rect 22569 11713 22603 11747
rect 22661 11713 22695 11747
rect 22845 11713 22879 11747
rect 23029 11713 23063 11747
rect 23213 11713 23247 11747
rect 24409 11713 24443 11747
rect 24501 11713 24535 11747
rect 24685 11713 24719 11747
rect 25237 11713 25271 11747
rect 26157 11713 26191 11747
rect 26341 11713 26375 11747
rect 27813 11713 27847 11747
rect 27905 11713 27939 11747
rect 28089 11713 28123 11747
rect 28181 11713 28215 11747
rect 28641 11713 28675 11747
rect 9229 11645 9263 11679
rect 10517 11645 10551 11679
rect 11621 11645 11655 11679
rect 13829 11645 13863 11679
rect 13921 11645 13955 11679
rect 14289 11645 14323 11679
rect 19901 11645 19935 11679
rect 20361 11645 20395 11679
rect 21925 11645 21959 11679
rect 25329 11645 25363 11679
rect 26065 11645 26099 11679
rect 28549 11645 28583 11679
rect 10977 11577 11011 11611
rect 11345 11577 11379 11611
rect 24869 11577 24903 11611
rect 28273 11577 28307 11611
rect 10149 11509 10183 11543
rect 11529 11509 11563 11543
rect 15117 11509 15151 11543
rect 16865 11509 16899 11543
rect 19349 11509 19383 11543
rect 19717 11509 19751 11543
rect 20821 11509 20855 11543
rect 23397 11509 23431 11543
rect 27629 11509 27663 11543
rect 9137 11305 9171 11339
rect 11253 11305 11287 11339
rect 11713 11305 11747 11339
rect 12081 11305 12115 11339
rect 14933 11305 14967 11339
rect 15485 11305 15519 11339
rect 16405 11305 16439 11339
rect 19625 11305 19659 11339
rect 25329 11305 25363 11339
rect 25513 11305 25547 11339
rect 27445 11305 27479 11339
rect 25237 11237 25271 11271
rect 9689 11169 9723 11203
rect 12265 11169 12299 11203
rect 12725 11169 12759 11203
rect 15393 11169 15427 11203
rect 15577 11169 15611 11203
rect 24869 11169 24903 11203
rect 27629 11169 27663 11203
rect 9321 11101 9355 11135
rect 9413 11101 9447 11135
rect 9781 11101 9815 11135
rect 10057 11101 10091 11135
rect 11161 11101 11195 11135
rect 12357 11101 12391 11135
rect 14841 11101 14875 11135
rect 15117 11101 15151 11135
rect 15209 11101 15243 11135
rect 15761 11101 15795 11135
rect 16405 11101 16439 11135
rect 16497 11101 16531 11135
rect 19533 11101 19567 11135
rect 19717 11101 19751 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 27721 11101 27755 11135
rect 28365 11101 28399 11135
rect 11069 11033 11103 11067
rect 12633 11033 12667 11067
rect 15485 11033 15519 11067
rect 16681 11033 16715 11067
rect 27997 11033 28031 11067
rect 28181 11033 28215 11067
rect 15945 10965 15979 10999
rect 16221 10965 16255 10999
rect 12725 10761 12759 10795
rect 21649 10761 21683 10795
rect 21833 10761 21867 10795
rect 24777 10761 24811 10795
rect 15025 10693 15059 10727
rect 16037 10693 16071 10727
rect 16129 10693 16163 10727
rect 10425 10625 10459 10659
rect 10885 10625 10919 10659
rect 12357 10625 12391 10659
rect 13001 10625 13035 10659
rect 13737 10625 13771 10659
rect 14841 10625 14875 10659
rect 15117 10625 15151 10659
rect 15209 10625 15243 10659
rect 15853 10625 15887 10659
rect 16221 10625 16255 10659
rect 17233 10625 17267 10659
rect 21373 10625 21407 10659
rect 21465 10625 21499 10659
rect 22017 10625 22051 10659
rect 22109 10625 22143 10659
rect 22201 10625 22235 10659
rect 22385 10625 22419 10659
rect 22477 10625 22511 10659
rect 23305 10625 23339 10659
rect 23603 10625 23637 10659
rect 24593 10625 24627 10659
rect 26525 10625 26559 10659
rect 26709 10625 26743 10659
rect 12449 10557 12483 10591
rect 17325 10557 17359 10591
rect 21189 10557 21223 10591
rect 21281 10557 21315 10591
rect 23489 10557 23523 10591
rect 24409 10557 24443 10591
rect 17601 10489 17635 10523
rect 23673 10489 23707 10523
rect 9321 10421 9355 10455
rect 15393 10421 15427 10455
rect 16405 10421 16439 10455
rect 23397 10421 23431 10455
rect 26525 10421 26559 10455
rect 10885 10217 10919 10251
rect 17601 10217 17635 10251
rect 18337 10217 18371 10251
rect 20821 10217 20855 10251
rect 22477 10217 22511 10251
rect 23397 10217 23431 10251
rect 23857 10217 23891 10251
rect 24133 10217 24167 10251
rect 24777 10217 24811 10251
rect 13921 10149 13955 10183
rect 18153 10149 18187 10183
rect 20177 10149 20211 10183
rect 12725 10081 12759 10115
rect 17509 10081 17543 10115
rect 18337 10081 18371 10115
rect 19809 10081 19843 10115
rect 20269 10081 20303 10115
rect 22661 10081 22695 10115
rect 22753 10081 22787 10115
rect 23581 10081 23615 10115
rect 26801 10081 26835 10115
rect 7297 10013 7331 10047
rect 7757 10013 7791 10047
rect 9045 10013 9079 10047
rect 9413 10013 9447 10047
rect 11713 10013 11747 10047
rect 13369 10013 13403 10047
rect 13645 10013 13679 10047
rect 13737 10013 13771 10047
rect 14105 10013 14139 10047
rect 14473 10013 14507 10047
rect 15761 10013 15795 10047
rect 15945 10013 15979 10047
rect 16129 10013 16163 10047
rect 16313 10013 16347 10047
rect 16497 10013 16531 10047
rect 17972 10013 18006 10047
rect 18521 10013 18555 10047
rect 18797 10013 18831 10047
rect 18981 10013 19015 10047
rect 19717 10013 19751 10047
rect 19901 10013 19935 10047
rect 19993 10013 20027 10047
rect 20545 10013 20579 10047
rect 21465 10013 21499 10047
rect 21741 10013 21775 10047
rect 21833 10013 21867 10047
rect 21944 10013 21978 10047
rect 22106 10013 22140 10047
rect 22385 10013 22419 10047
rect 23673 10013 23707 10047
rect 24501 10013 24535 10047
rect 24593 10013 24627 10047
rect 24961 10013 24995 10047
rect 25145 10013 25179 10047
rect 26985 10013 27019 10047
rect 27169 10013 27203 10047
rect 27261 10013 27295 10047
rect 27445 10013 27479 10047
rect 13553 9945 13587 9979
rect 14289 9945 14323 9979
rect 14381 9945 14415 9979
rect 18245 9945 18279 9979
rect 20637 9945 20671 9979
rect 21557 9945 21591 9979
rect 23397 9945 23431 9979
rect 14657 9877 14691 9911
rect 17969 9877 18003 9911
rect 18705 9877 18739 9911
rect 18889 9877 18923 9911
rect 20453 9877 20487 9911
rect 22293 9877 22327 9911
rect 22753 9877 22787 9911
rect 25053 9877 25087 9911
rect 27353 9877 27387 9911
rect 20545 9673 20579 9707
rect 21557 9673 21591 9707
rect 24041 9673 24075 9707
rect 24777 9673 24811 9707
rect 13553 9605 13587 9639
rect 17509 9605 17543 9639
rect 21189 9605 21223 9639
rect 23029 9605 23063 9639
rect 26065 9605 26099 9639
rect 8769 9537 8803 9571
rect 9229 9537 9263 9571
rect 11897 9537 11931 9571
rect 12081 9537 12115 9571
rect 17785 9537 17819 9571
rect 17969 9537 18003 9571
rect 18061 9537 18095 9571
rect 18245 9537 18279 9571
rect 19717 9537 19751 9571
rect 20177 9537 20211 9571
rect 20361 9537 20395 9571
rect 21373 9537 21407 9571
rect 22109 9537 22143 9571
rect 22293 9537 22327 9571
rect 23765 9537 23799 9571
rect 23857 9537 23891 9571
rect 24133 9537 24167 9571
rect 24593 9537 24627 9571
rect 24869 9537 24903 9571
rect 25053 9537 25087 9571
rect 25421 9537 25455 9571
rect 25789 9537 25823 9571
rect 27169 9537 27203 9571
rect 17601 9469 17635 9503
rect 19809 9469 19843 9503
rect 20085 9469 20119 9503
rect 23397 9469 23431 9503
rect 23489 9469 23523 9503
rect 24409 9469 24443 9503
rect 25697 9469 25731 9503
rect 25881 9469 25915 9503
rect 27261 9469 27295 9503
rect 27537 9469 27571 9503
rect 25605 9401 25639 9435
rect 17693 9333 17727 9367
rect 18061 9333 18095 9367
rect 22201 9333 22235 9367
rect 24225 9333 24259 9367
rect 25053 9333 25087 9367
rect 25237 9333 25271 9367
rect 25789 9333 25823 9367
rect 11897 9129 11931 9163
rect 14841 9129 14875 9163
rect 15853 9129 15887 9163
rect 16589 9129 16623 9163
rect 21649 9129 21683 9163
rect 23765 9129 23799 9163
rect 24961 9129 24995 9163
rect 27537 9129 27571 9163
rect 14381 9061 14415 9095
rect 16221 9061 16255 9095
rect 23305 9061 23339 9095
rect 27169 9061 27203 9095
rect 15025 8993 15059 9027
rect 15235 8993 15269 9027
rect 20913 8993 20947 9027
rect 21833 8993 21867 9027
rect 24593 8993 24627 9027
rect 10241 8925 10275 8959
rect 10425 8925 10459 8959
rect 14289 8925 14323 8959
rect 14473 8925 14507 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 15393 8925 15427 8959
rect 15485 8925 15519 8959
rect 15853 8925 15887 8959
rect 16129 8925 16163 8959
rect 16405 8925 16439 8959
rect 16773 8925 16807 8959
rect 16865 8925 16899 8959
rect 17049 8925 17083 8959
rect 17141 8925 17175 8959
rect 17325 8925 17359 8959
rect 17693 8925 17727 8959
rect 20821 8925 20855 8959
rect 21005 8925 21039 8959
rect 21097 8925 21131 8959
rect 21465 8925 21499 8959
rect 22017 8925 22051 8959
rect 23857 8925 23891 8959
rect 24777 8925 24811 8959
rect 25237 8925 25271 8959
rect 25421 8925 25455 8959
rect 27905 8925 27939 8959
rect 28089 8925 28123 8959
rect 17601 8857 17635 8891
rect 21281 8857 21315 8891
rect 21373 8857 21407 8891
rect 27537 8857 27571 8891
rect 14657 8789 14691 8823
rect 15669 8789 15703 8823
rect 22201 8789 22235 8823
rect 24225 8789 24259 8823
rect 25329 8789 25363 8823
rect 27721 8789 27755 8823
rect 28917 8789 28951 8823
rect 10517 8585 10551 8619
rect 14749 8585 14783 8619
rect 15393 8585 15427 8619
rect 19901 8585 19935 8619
rect 23673 8585 23707 8619
rect 27185 8585 27219 8619
rect 27353 8585 27387 8619
rect 27537 8585 27571 8619
rect 28089 8585 28123 8619
rect 6837 8517 6871 8551
rect 12173 8517 12207 8551
rect 17509 8517 17543 8551
rect 26525 8517 26559 8551
rect 26709 8517 26743 8551
rect 26985 8517 27019 8551
rect 7297 8449 7331 8483
rect 7573 8449 7607 8483
rect 7849 8449 7883 8483
rect 8033 8449 8067 8483
rect 8217 8449 8251 8483
rect 8769 8449 8803 8483
rect 9413 8449 9447 8483
rect 10701 8449 10735 8483
rect 10977 8449 11011 8483
rect 11161 8449 11195 8483
rect 11529 8449 11563 8483
rect 11713 8449 11747 8483
rect 11805 8449 11839 8483
rect 11898 8449 11932 8483
rect 12725 8449 12759 8483
rect 13093 8449 13127 8483
rect 14657 8449 14691 8483
rect 15025 8449 15059 8483
rect 16773 8449 16807 8483
rect 18705 8449 18739 8483
rect 18889 8449 18923 8483
rect 18981 8449 19015 8483
rect 19349 8449 19383 8483
rect 20545 8449 20579 8483
rect 23857 8449 23891 8483
rect 24041 8449 24075 8483
rect 25053 8449 25087 8483
rect 25237 8449 25271 8483
rect 26801 8449 26835 8483
rect 27445 8449 27479 8483
rect 27629 8449 27663 8483
rect 27721 8449 27755 8483
rect 27814 8449 27848 8483
rect 10149 8381 10183 8415
rect 10885 8381 10919 8415
rect 14565 8381 14599 8415
rect 15117 8381 15151 8415
rect 20085 8381 20119 8415
rect 20177 8381 20211 8415
rect 24225 8381 24259 8415
rect 10793 8313 10827 8347
rect 14933 8313 14967 8347
rect 25513 8313 25547 8347
rect 26525 8313 26559 8347
rect 24501 8245 24535 8279
rect 25237 8245 25271 8279
rect 27169 8245 27203 8279
rect 12265 8041 12299 8075
rect 12449 8041 12483 8075
rect 19073 8041 19107 8075
rect 23305 8041 23339 8075
rect 25421 8041 25455 8075
rect 25881 8041 25915 8075
rect 26525 8041 26559 8075
rect 23397 7973 23431 8007
rect 24777 7973 24811 8007
rect 24869 7973 24903 8007
rect 26433 7973 26467 8007
rect 9229 7905 9263 7939
rect 9505 7905 9539 7939
rect 12909 7905 12943 7939
rect 13737 7905 13771 7939
rect 18337 7905 18371 7939
rect 18889 7905 18923 7939
rect 20545 7905 20579 7939
rect 23489 7905 23523 7939
rect 23581 7905 23615 7939
rect 25145 7905 25179 7939
rect 9597 7837 9631 7871
rect 9965 7837 9999 7871
rect 10149 7837 10183 7871
rect 10425 7837 10459 7871
rect 10609 7837 10643 7871
rect 15025 7837 15059 7871
rect 15209 7837 15243 7871
rect 15301 7837 15335 7871
rect 15485 7837 15519 7871
rect 17877 7837 17911 7871
rect 18153 7837 18187 7871
rect 18429 7837 18463 7871
rect 18797 7837 18831 7871
rect 19809 7837 19843 7871
rect 20085 7837 20119 7871
rect 20177 7837 20211 7871
rect 20269 7837 20303 7871
rect 20637 7837 20671 7871
rect 20913 7837 20947 7871
rect 21189 7837 21223 7871
rect 21373 7837 21407 7871
rect 21649 7837 21683 7871
rect 21833 7837 21867 7871
rect 23121 7837 23155 7871
rect 23213 7837 23247 7871
rect 23856 7837 23890 7871
rect 23949 7837 23983 7871
rect 24501 7837 24535 7871
rect 24685 7837 24719 7871
rect 24961 7837 24995 7871
rect 25237 7837 25271 7871
rect 25513 7837 25547 7871
rect 26157 7837 26191 7871
rect 26525 7837 26559 7871
rect 26709 7837 26743 7871
rect 10701 7769 10735 7803
rect 12081 7769 12115 7803
rect 12265 7769 12299 7803
rect 25329 7769 25363 7803
rect 25697 7769 25731 7803
rect 26249 7769 26283 7803
rect 26433 7769 26467 7803
rect 15025 7701 15059 7735
rect 15393 7701 15427 7735
rect 17969 7701 18003 7735
rect 19901 7701 19935 7735
rect 20729 7701 20763 7735
rect 21097 7701 21131 7735
rect 21281 7701 21315 7735
rect 21833 7701 21867 7735
rect 25897 7701 25931 7735
rect 26065 7701 26099 7735
rect 16129 7497 16163 7531
rect 18521 7497 18555 7531
rect 20269 7497 20303 7531
rect 21465 7497 21499 7531
rect 23029 7497 23063 7531
rect 23397 7497 23431 7531
rect 25421 7497 25455 7531
rect 26801 7497 26835 7531
rect 18245 7429 18279 7463
rect 20637 7429 20671 7463
rect 8861 7361 8895 7395
rect 8953 7361 8987 7395
rect 10333 7361 10367 7395
rect 10701 7361 10735 7395
rect 12633 7361 12667 7395
rect 12909 7361 12943 7395
rect 13553 7361 13587 7395
rect 14841 7361 14875 7395
rect 15117 7361 15151 7395
rect 16037 7361 16071 7395
rect 16313 7361 16347 7395
rect 16773 7361 16807 7395
rect 17141 7361 17175 7395
rect 18429 7361 18463 7395
rect 18521 7361 18555 7395
rect 20269 7361 20303 7395
rect 20453 7361 20487 7395
rect 20821 7361 20855 7395
rect 20911 7383 20945 7417
rect 21005 7361 21039 7395
rect 21097 7361 21131 7395
rect 21281 7361 21315 7395
rect 22187 7361 22221 7395
rect 23673 7361 23707 7395
rect 23857 7361 23891 7395
rect 23949 7361 23983 7395
rect 24041 7361 24075 7395
rect 25053 7361 25087 7395
rect 26801 7361 26835 7395
rect 27261 7361 27295 7395
rect 27721 7361 27755 7395
rect 27813 7361 27847 7395
rect 27997 7361 28031 7395
rect 28089 7361 28123 7395
rect 28365 7361 28399 7395
rect 28549 7361 28583 7395
rect 10425 7293 10459 7327
rect 11069 7293 11103 7327
rect 12725 7293 12759 7327
rect 13277 7293 13311 7327
rect 14473 7293 14507 7327
rect 14933 7293 14967 7327
rect 15025 7293 15059 7327
rect 16497 7293 16531 7327
rect 17785 7293 17819 7327
rect 22109 7293 22143 7327
rect 24317 7293 24351 7327
rect 24961 7293 24995 7327
rect 26525 7293 26559 7327
rect 26985 7293 27019 7327
rect 27077 7293 27111 7327
rect 28457 7293 28491 7327
rect 9321 7225 9355 7259
rect 13093 7225 13127 7259
rect 14197 7225 14231 7259
rect 20913 7225 20947 7259
rect 26709 7225 26743 7259
rect 27445 7225 27479 7259
rect 12725 7157 12759 7191
rect 15301 7157 15335 7191
rect 22385 7157 22419 7191
rect 28273 7157 28307 7191
rect 8309 6953 8343 6987
rect 9275 6953 9309 6987
rect 16037 6953 16071 6987
rect 17785 6953 17819 6987
rect 21189 6953 21223 6987
rect 23581 6953 23615 6987
rect 9413 6885 9447 6919
rect 7849 6817 7883 6851
rect 9505 6817 9539 6851
rect 18521 6817 18555 6851
rect 18981 6817 19015 6851
rect 28181 6817 28215 6851
rect 28457 6817 28491 6851
rect 8125 6749 8159 6783
rect 10425 6749 10459 6783
rect 10701 6749 10735 6783
rect 12633 6749 12667 6783
rect 13185 6749 13219 6783
rect 14197 6749 14231 6783
rect 14565 6749 14599 6783
rect 16129 6749 16163 6783
rect 16221 6749 16255 6783
rect 16405 6749 16439 6783
rect 17509 6749 17543 6783
rect 17785 6749 17819 6783
rect 18613 6749 18647 6783
rect 19441 6749 19475 6783
rect 19625 6749 19659 6783
rect 19809 6749 19843 6783
rect 20177 6749 20211 6783
rect 20361 6749 20395 6783
rect 21281 6749 21315 6783
rect 21373 6749 21407 6783
rect 28089 6749 28123 6783
rect 8033 6681 8067 6715
rect 9137 6681 9171 6715
rect 17693 6681 17727 6715
rect 21097 6681 21131 6715
rect 9781 6613 9815 6647
rect 16589 6613 16623 6647
rect 19993 6613 20027 6647
rect 14841 6409 14875 6443
rect 14933 6409 14967 6443
rect 16329 6409 16363 6443
rect 17233 6409 17267 6443
rect 17877 6409 17911 6443
rect 19533 6409 19567 6443
rect 11345 6341 11379 6375
rect 14013 6341 14047 6375
rect 14749 6341 14783 6375
rect 16129 6341 16163 6375
rect 17693 6341 17727 6375
rect 8309 6273 8343 6307
rect 8585 6273 8619 6307
rect 9689 6273 9723 6307
rect 10241 6273 10275 6307
rect 12081 6273 12115 6307
rect 13277 6273 13311 6307
rect 13737 6273 13771 6307
rect 15301 6273 15335 6307
rect 15485 6273 15519 6307
rect 17969 6273 18003 6307
rect 18153 6273 18187 6307
rect 18245 6273 18279 6307
rect 19441 6273 19475 6307
rect 19625 6273 19659 6307
rect 11621 6205 11655 6239
rect 12817 6205 12851 6239
rect 13001 6205 13035 6239
rect 16773 6205 16807 6239
rect 17325 6205 17359 6239
rect 12541 6137 12575 6171
rect 14565 6137 14599 6171
rect 15117 6137 15151 6171
rect 16497 6137 16531 6171
rect 17049 6137 17083 6171
rect 18337 6137 18371 6171
rect 15393 6069 15427 6103
rect 16313 6069 16347 6103
rect 17693 6069 17727 6103
rect 18153 6069 18187 6103
rect 9091 5865 9125 5899
rect 10149 5865 10183 5899
rect 10793 5865 10827 5899
rect 11253 5865 11287 5899
rect 13185 5865 13219 5899
rect 14841 5865 14875 5899
rect 15301 5865 15335 5899
rect 17417 5865 17451 5899
rect 22937 5865 22971 5899
rect 23765 5865 23799 5899
rect 9229 5797 9263 5831
rect 9597 5797 9631 5831
rect 12817 5797 12851 5831
rect 23121 5797 23155 5831
rect 26709 5797 26743 5831
rect 27169 5797 27203 5831
rect 7205 5729 7239 5763
rect 9321 5729 9355 5763
rect 10885 5729 10919 5763
rect 12541 5729 12575 5763
rect 20361 5729 20395 5763
rect 20545 5729 20579 5763
rect 21005 5729 21039 5763
rect 22477 5729 22511 5763
rect 23029 5729 23063 5763
rect 23489 5729 23523 5763
rect 23581 5729 23615 5763
rect 27353 5729 27387 5763
rect 5181 5661 5215 5695
rect 10333 5661 10367 5695
rect 10425 5661 10459 5695
rect 10517 5661 10551 5695
rect 10609 5661 10643 5695
rect 10793 5661 10827 5695
rect 11069 5661 11103 5695
rect 12265 5661 12299 5695
rect 12449 5661 12483 5695
rect 12725 5661 12759 5695
rect 12909 5661 12943 5695
rect 13001 5661 13035 5695
rect 14749 5661 14783 5695
rect 14933 5661 14967 5695
rect 15209 5661 15243 5695
rect 17325 5661 17359 5695
rect 17509 5661 17543 5695
rect 18153 5661 18187 5695
rect 18337 5661 18371 5695
rect 19717 5661 19751 5695
rect 19901 5661 19935 5695
rect 20177 5661 20211 5695
rect 20637 5661 20671 5695
rect 22569 5661 22603 5695
rect 23305 5661 23339 5695
rect 23857 5661 23891 5695
rect 24501 5661 24535 5695
rect 24685 5661 24719 5695
rect 24961 5661 24995 5695
rect 26525 5661 26559 5695
rect 26709 5661 26743 5695
rect 27077 5661 27111 5695
rect 28181 5661 28215 5695
rect 28273 5661 28307 5695
rect 28457 5661 28491 5695
rect 28549 5661 28583 5695
rect 5457 5593 5491 5627
rect 8953 5593 8987 5627
rect 19809 5593 19843 5627
rect 18245 5525 18279 5559
rect 19993 5525 20027 5559
rect 23581 5525 23615 5559
rect 25145 5525 25179 5559
rect 27353 5525 27387 5559
rect 28733 5525 28767 5559
rect 15393 5321 15427 5355
rect 22937 5321 22971 5355
rect 26985 5321 27019 5355
rect 8493 5253 8527 5287
rect 12817 5253 12851 5287
rect 15761 5253 15795 5287
rect 28181 5253 28215 5287
rect 30389 5253 30423 5287
rect 11621 5185 11655 5219
rect 12357 5185 12391 5219
rect 13737 5185 13771 5219
rect 14657 5185 14691 5219
rect 15301 5185 15335 5219
rect 15577 5185 15611 5219
rect 15853 5185 15887 5219
rect 16037 5185 16071 5219
rect 16313 5185 16347 5219
rect 16497 5185 16531 5219
rect 16773 5185 16807 5219
rect 16957 5185 16991 5219
rect 19993 5185 20027 5219
rect 20177 5185 20211 5219
rect 21465 5185 21499 5219
rect 22293 5185 22327 5219
rect 22477 5185 22511 5219
rect 22753 5185 22787 5219
rect 23581 5185 23615 5219
rect 24317 5185 24351 5219
rect 25421 5185 25455 5219
rect 25881 5185 25915 5219
rect 26249 5185 26283 5219
rect 26433 5185 26467 5219
rect 27353 5185 27387 5219
rect 27629 5185 27663 5219
rect 27721 5185 27755 5219
rect 27905 5185 27939 5219
rect 27997 5185 28031 5219
rect 28365 5185 28399 5219
rect 28457 5185 28491 5219
rect 28641 5185 28675 5219
rect 28733 5185 28767 5219
rect 29377 5185 29411 5219
rect 6469 5117 6503 5151
rect 6745 5117 6779 5151
rect 11529 5117 11563 5151
rect 12081 5117 12115 5151
rect 12265 5117 12299 5151
rect 15209 5117 15243 5151
rect 16681 5117 16715 5151
rect 21189 5117 21223 5151
rect 23673 5117 23707 5151
rect 24409 5117 24443 5151
rect 25513 5117 25547 5151
rect 27445 5117 27479 5151
rect 29285 5117 29319 5151
rect 30113 5117 30147 5151
rect 24685 5049 24719 5083
rect 25789 5049 25823 5083
rect 28917 5049 28951 5083
rect 16037 4981 16071 5015
rect 16313 4981 16347 5015
rect 17141 4981 17175 5015
rect 19993 4981 20027 5015
rect 21281 4981 21315 5015
rect 21373 4981 21407 5015
rect 23949 4981 23983 5015
rect 25973 4981 26007 5015
rect 29009 4981 29043 5015
rect 31861 4981 31895 5015
rect 11161 4777 11195 4811
rect 27169 4777 27203 4811
rect 19901 4709 19935 4743
rect 20269 4709 20303 4743
rect 21189 4709 21223 4743
rect 27537 4709 27571 4743
rect 7205 4641 7239 4675
rect 8953 4641 8987 4675
rect 10977 4641 11011 4675
rect 12909 4641 12943 4675
rect 16405 4641 16439 4675
rect 17877 4641 17911 4675
rect 18705 4641 18739 4675
rect 19625 4641 19659 4675
rect 20913 4641 20947 4675
rect 22201 4641 22235 4675
rect 27261 4641 27295 4675
rect 27629 4641 27663 4675
rect 5181 4573 5215 4607
rect 14197 4573 14231 4607
rect 14749 4573 14783 4607
rect 16497 4573 16531 4607
rect 17785 4573 17819 4607
rect 18245 4573 18279 4607
rect 18613 4573 18647 4607
rect 18889 4573 18923 4607
rect 19533 4573 19567 4607
rect 19993 4573 20027 4607
rect 20821 4573 20855 4607
rect 22109 4573 22143 4607
rect 25605 4573 25639 4607
rect 27169 4573 27203 4607
rect 27813 4573 27847 4607
rect 5457 4505 5491 4539
rect 9229 4505 9263 4539
rect 12633 4505 12667 4539
rect 20269 4505 20303 4539
rect 24869 4505 24903 4539
rect 16865 4437 16899 4471
rect 18153 4437 18187 4471
rect 20085 4437 20119 4471
rect 22477 4437 22511 4471
rect 27997 4437 28031 4471
rect 8401 4165 8435 4199
rect 11989 4165 12023 4199
rect 15393 4097 15427 4131
rect 15853 4097 15887 4131
rect 16037 4097 16071 4131
rect 16773 4097 16807 4131
rect 18245 4097 18279 4131
rect 23581 4097 23615 4131
rect 23949 4097 23983 4131
rect 26525 4097 26559 4131
rect 26985 4097 27019 4131
rect 28825 4097 28859 4131
rect 6377 4029 6411 4063
rect 6653 4029 6687 4063
rect 8493 4029 8527 4063
rect 8769 4029 8803 4063
rect 10241 4029 10275 4063
rect 13737 4029 13771 4063
rect 14013 4029 14047 4063
rect 15301 4029 15335 4063
rect 15945 4029 15979 4063
rect 17233 4029 17267 4063
rect 18705 4029 18739 4063
rect 22477 4029 22511 4063
rect 24225 4029 24259 4063
rect 25513 4029 25547 4063
rect 27445 4029 27479 4063
rect 29101 4029 29135 4063
rect 14381 3893 14415 3927
rect 15669 3893 15703 3927
rect 30573 3893 30607 3927
rect 18061 3689 18095 3723
rect 23949 3689 23983 3723
rect 26157 3689 26191 3723
rect 4629 3553 4663 3587
rect 8769 3553 8803 3587
rect 11805 3553 11839 3587
rect 16589 3553 16623 3587
rect 19349 3553 19383 3587
rect 22201 3553 22235 3587
rect 22477 3553 22511 3587
rect 24685 3553 24719 3587
rect 26525 3553 26559 3587
rect 27997 3553 28031 3587
rect 30021 3553 30055 3587
rect 31493 3553 31527 3587
rect 32965 3553 32999 3587
rect 6653 3485 6687 3519
rect 6745 3485 6779 3519
rect 9781 3485 9815 3519
rect 11897 3485 11931 3519
rect 13921 3485 13955 3519
rect 16313 3485 16347 3519
rect 18613 3485 18647 3519
rect 19901 3485 19935 3519
rect 21925 3485 21959 3519
rect 24409 3485 24443 3519
rect 26249 3485 26283 3519
rect 28733 3485 28767 3519
rect 29561 3485 29595 3519
rect 31033 3485 31067 3519
rect 32505 3485 32539 3519
rect 4905 3417 4939 3451
rect 7021 3417 7055 3451
rect 10057 3417 10091 3451
rect 13645 3417 13679 3451
rect 18337 3417 18371 3451
rect 21097 3417 21131 3451
rect 28917 3349 28951 3383
rect 13185 3145 13219 3179
rect 21557 3145 21591 3179
rect 25421 3145 25455 3179
rect 28733 3145 28767 3179
rect 33609 3145 33643 3179
rect 8953 3077 8987 3111
rect 10793 3077 10827 3111
rect 13553 3077 13587 3111
rect 15301 3077 15335 3111
rect 18245 3077 18279 3111
rect 22109 3077 22143 3111
rect 23949 3077 23983 3111
rect 29101 3077 29135 3111
rect 30941 3077 30975 3111
rect 6929 3009 6963 3043
rect 11989 3009 12023 3043
rect 13369 3009 13403 3043
rect 15577 3009 15611 3043
rect 23673 3009 23707 3043
rect 28825 3009 28859 3043
rect 30665 3009 30699 3043
rect 32137 3009 32171 3043
rect 33793 3009 33827 3043
rect 4169 2941 4203 2975
rect 4445 2941 4479 2975
rect 6193 2941 6227 2975
rect 7205 2941 7239 2975
rect 9045 2941 9079 2975
rect 11069 2941 11103 2975
rect 17969 2941 18003 2975
rect 19809 2941 19843 2975
rect 20085 2941 20119 2975
rect 21833 2941 21867 2975
rect 26985 2941 27019 2975
rect 32597 2941 32631 2975
rect 23581 2873 23615 2907
rect 11805 2805 11839 2839
rect 19717 2805 19751 2839
rect 27242 2805 27276 2839
rect 30573 2805 30607 2839
rect 3249 2601 3283 2635
rect 5273 2601 5307 2635
rect 6561 2601 6595 2635
rect 7113 2601 7147 2635
rect 8125 2601 8159 2635
rect 9321 2601 9355 2635
rect 10149 2601 10183 2635
rect 11161 2601 11195 2635
rect 14197 2601 14231 2635
rect 14473 2601 14507 2635
rect 16497 2601 16531 2635
rect 26433 2601 26467 2635
rect 29285 2601 29319 2635
rect 1593 2533 1627 2567
rect 16681 2533 16715 2567
rect 34713 2533 34747 2567
rect 11529 2465 11563 2499
rect 11805 2465 11839 2499
rect 13553 2465 13587 2499
rect 14749 2465 14783 2499
rect 15025 2465 15059 2499
rect 17601 2465 17635 2499
rect 19073 2465 19107 2499
rect 19717 2465 19751 2499
rect 22293 2465 22327 2499
rect 24685 2465 24719 2499
rect 24961 2465 24995 2499
rect 27537 2465 27571 2499
rect 27813 2465 27847 2499
rect 32597 2465 32631 2499
rect 34253 2465 34287 2499
rect 1409 2397 1443 2431
rect 2053 2397 2087 2431
rect 3065 2397 3099 2431
rect 4077 2397 4111 2431
rect 5089 2397 5123 2431
rect 6377 2397 6411 2431
rect 7297 2397 7331 2431
rect 8309 2397 8343 2431
rect 9137 2397 9171 2431
rect 10333 2397 10367 2431
rect 11345 2397 11379 2431
rect 14381 2397 14415 2431
rect 14657 2397 14691 2431
rect 16865 2397 16899 2431
rect 17325 2397 17359 2431
rect 19257 2397 19291 2431
rect 21833 2397 21867 2431
rect 29561 2397 29595 2431
rect 32137 2397 32171 2431
rect 34529 2397 34563 2431
rect 34897 2397 34931 2431
rect 30481 2329 30515 2363
rect 2237 2261 2271 2295
rect 4261 2261 4295 2295
<< metal1 >>
rect 1104 36474 35248 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 35248 36474
rect 1104 36400 35248 36422
rect 1104 35930 35236 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 35236 35930
rect 1104 35856 35236 35878
rect 1104 35386 35248 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 35248 35386
rect 1104 35312 35248 35334
rect 1104 34842 35236 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 35236 34842
rect 1104 34768 35236 34790
rect 1104 34298 35248 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 35248 34298
rect 1104 34224 35248 34246
rect 1104 33754 35236 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 35236 33754
rect 1104 33680 35236 33702
rect 1104 33210 35248 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 35248 33210
rect 1104 33136 35248 33158
rect 1104 32666 35236 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 35236 32666
rect 1104 32592 35236 32614
rect 1104 32122 35248 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 35248 32122
rect 1104 32048 35248 32070
rect 1104 31578 35236 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 35236 31578
rect 1104 31504 35236 31526
rect 1104 31034 35248 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 35248 31034
rect 1104 30960 35248 30982
rect 1104 30490 35236 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 35236 30490
rect 1104 30416 35236 30438
rect 1104 29946 35248 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 35248 29946
rect 1104 29872 35248 29894
rect 1104 29402 35236 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 35236 29402
rect 1104 29328 35236 29350
rect 1104 28858 35248 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 35248 28858
rect 1104 28784 35248 28806
rect 1104 28314 35236 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 35236 28314
rect 1104 28240 35236 28262
rect 1104 27770 35248 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 35248 27770
rect 1104 27696 35248 27718
rect 1104 27226 35236 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 35236 27226
rect 1104 27152 35236 27174
rect 1104 26682 35248 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 35248 26682
rect 1104 26608 35248 26630
rect 1104 26138 35236 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 35236 26138
rect 1104 26064 35236 26086
rect 1104 25594 35248 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 35248 25594
rect 1104 25520 35248 25542
rect 1104 25050 35236 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 35236 25050
rect 1104 24976 35236 24998
rect 1104 24506 35248 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 35248 24506
rect 1104 24432 35248 24454
rect 1104 23962 35236 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 35236 23962
rect 1104 23888 35236 23910
rect 1104 23418 35248 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 35248 23418
rect 1104 23344 35248 23366
rect 1104 22874 35236 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 35236 22874
rect 1104 22800 35236 22822
rect 1104 22330 35248 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 35248 22330
rect 1104 22256 35248 22278
rect 1104 21786 35236 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 35236 21786
rect 1104 21712 35236 21734
rect 1104 21242 35248 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 35248 21242
rect 1104 21168 35248 21190
rect 1104 20698 35236 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 35236 20698
rect 1104 20624 35236 20646
rect 1104 20154 35248 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 35248 20154
rect 1104 20080 35248 20102
rect 1104 19610 35236 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 35236 19610
rect 1104 19536 35236 19558
rect 18046 19320 18052 19372
rect 18104 19360 18110 19372
rect 18233 19363 18291 19369
rect 18233 19360 18245 19363
rect 18104 19332 18245 19360
rect 18104 19320 18110 19332
rect 18233 19329 18245 19332
rect 18279 19329 18291 19363
rect 18233 19323 18291 19329
rect 18141 19295 18199 19301
rect 18141 19261 18153 19295
rect 18187 19292 18199 19295
rect 18187 19264 18276 19292
rect 18187 19261 18199 19264
rect 18141 19255 18199 19261
rect 18248 19168 18276 19264
rect 18230 19116 18236 19168
rect 18288 19116 18294 19168
rect 18506 19116 18512 19168
rect 18564 19116 18570 19168
rect 1104 19066 35248 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 35248 19066
rect 1104 18992 35248 19014
rect 20070 18884 20076 18896
rect 13280 18856 20076 18884
rect 13280 18825 13308 18856
rect 13265 18819 13323 18825
rect 13265 18785 13277 18819
rect 13311 18785 13323 18819
rect 13265 18779 13323 18785
rect 16393 18819 16451 18825
rect 16393 18785 16405 18819
rect 16439 18816 16451 18819
rect 16574 18816 16580 18828
rect 16439 18788 16580 18816
rect 16439 18785 16451 18788
rect 16393 18779 16451 18785
rect 16574 18776 16580 18788
rect 16632 18776 16638 18828
rect 18046 18776 18052 18828
rect 18104 18776 18110 18828
rect 18506 18776 18512 18828
rect 18564 18776 18570 18828
rect 19904 18825 19932 18856
rect 20070 18844 20076 18856
rect 20128 18884 20134 18896
rect 20990 18884 20996 18896
rect 20128 18856 20996 18884
rect 20128 18844 20134 18856
rect 20990 18844 20996 18856
rect 21048 18844 21054 18896
rect 19889 18819 19947 18825
rect 19889 18785 19901 18819
rect 19935 18785 19947 18819
rect 19889 18779 19947 18785
rect 19996 18788 21496 18816
rect 12618 18708 12624 18760
rect 12676 18708 12682 18760
rect 12710 18708 12716 18760
rect 12768 18708 12774 18760
rect 16482 18708 16488 18760
rect 16540 18708 16546 18760
rect 18230 18708 18236 18760
rect 18288 18708 18294 18760
rect 18524 18748 18552 18776
rect 19996 18760 20024 18788
rect 19978 18748 19984 18760
rect 18524 18720 19984 18748
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20622 18708 20628 18760
rect 20680 18708 20686 18760
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 20947 18720 21373 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 18248 18680 18276 18708
rect 16868 18652 18276 18680
rect 20441 18683 20499 18689
rect 16868 18621 16896 18652
rect 20441 18649 20453 18683
rect 20487 18680 20499 18683
rect 20487 18652 20944 18680
rect 20487 18649 20499 18652
rect 20441 18643 20499 18649
rect 20916 18624 20944 18652
rect 20990 18640 20996 18692
rect 21048 18640 21054 18692
rect 21177 18683 21235 18689
rect 21177 18649 21189 18683
rect 21223 18680 21235 18683
rect 21468 18680 21496 18788
rect 21223 18652 21496 18680
rect 21223 18649 21235 18652
rect 21177 18643 21235 18649
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18581 16911 18615
rect 16853 18575 16911 18581
rect 18414 18572 18420 18624
rect 18472 18572 18478 18624
rect 20346 18572 20352 18624
rect 20404 18572 20410 18624
rect 20806 18572 20812 18624
rect 20864 18572 20870 18624
rect 20898 18572 20904 18624
rect 20956 18572 20962 18624
rect 1104 18522 35236 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 35236 18522
rect 1104 18448 35236 18470
rect 12710 18368 12716 18420
rect 12768 18368 12774 18420
rect 19978 18368 19984 18420
rect 20036 18368 20042 18420
rect 20070 18368 20076 18420
rect 20128 18368 20134 18420
rect 20349 18411 20407 18417
rect 20349 18377 20361 18411
rect 20395 18408 20407 18411
rect 20622 18408 20628 18420
rect 20395 18380 20628 18408
rect 20395 18377 20407 18380
rect 20349 18371 20407 18377
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 12621 18343 12679 18349
rect 12621 18309 12633 18343
rect 12667 18340 12679 18343
rect 12728 18340 12756 18368
rect 12667 18312 12756 18340
rect 12667 18309 12679 18312
rect 12621 18303 12679 18309
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 12728 18272 12756 18312
rect 15565 18343 15623 18349
rect 15565 18309 15577 18343
rect 15611 18340 15623 18343
rect 16574 18340 16580 18352
rect 15611 18312 16580 18340
rect 15611 18309 15623 18312
rect 15565 18303 15623 18309
rect 16574 18300 16580 18312
rect 16632 18300 16638 18352
rect 17954 18300 17960 18352
rect 18012 18340 18018 18352
rect 18414 18340 18420 18352
rect 18012 18312 18420 18340
rect 18012 18300 18018 18312
rect 18414 18300 18420 18312
rect 18472 18300 18478 18352
rect 12897 18275 12955 18281
rect 12897 18272 12909 18275
rect 11388 18244 11730 18272
rect 12728 18244 12909 18272
rect 11388 18232 11394 18244
rect 12897 18241 12909 18244
rect 12943 18241 12955 18275
rect 12897 18235 12955 18241
rect 14274 18232 14280 18284
rect 14332 18272 14338 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14332 18244 14565 18272
rect 14332 18232 14338 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 15344 18244 15669 18272
rect 15344 18232 15350 18244
rect 15657 18241 15669 18244
rect 15703 18241 15715 18275
rect 15657 18235 15715 18241
rect 15746 18232 15752 18284
rect 15804 18232 15810 18284
rect 15933 18275 15991 18281
rect 15933 18241 15945 18275
rect 15979 18241 15991 18275
rect 15933 18235 15991 18241
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11793 18207 11851 18213
rect 11793 18204 11805 18207
rect 11572 18176 11805 18204
rect 11572 18164 11578 18176
rect 11793 18173 11805 18176
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12713 18207 12771 18213
rect 12713 18204 12725 18207
rect 12676 18176 12725 18204
rect 12676 18164 12682 18176
rect 12713 18173 12725 18176
rect 12759 18173 12771 18207
rect 15948 18204 15976 18235
rect 18506 18232 18512 18284
rect 18564 18272 18570 18284
rect 19996 18281 20024 18368
rect 18601 18275 18659 18281
rect 18601 18272 18613 18275
rect 18564 18244 18613 18272
rect 18564 18232 18570 18244
rect 18601 18241 18613 18244
rect 18647 18241 18659 18275
rect 18601 18235 18659 18241
rect 18693 18275 18751 18281
rect 18693 18241 18705 18275
rect 18739 18241 18751 18275
rect 18693 18235 18751 18241
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18241 20039 18275
rect 20088 18272 20116 18368
rect 20438 18300 20444 18352
rect 20496 18340 20502 18352
rect 20806 18340 20812 18352
rect 20496 18312 20812 18340
rect 20496 18300 20502 18312
rect 20806 18300 20812 18312
rect 20864 18340 20870 18352
rect 20864 18312 20944 18340
rect 20864 18300 20870 18312
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 20088 18244 20177 18272
rect 19981 18235 20039 18241
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20165 18235 20223 18241
rect 12713 18167 12771 18173
rect 15212 18176 15976 18204
rect 15212 18080 15240 18176
rect 18322 18164 18328 18216
rect 18380 18204 18386 18216
rect 18708 18204 18736 18235
rect 20346 18232 20352 18284
rect 20404 18272 20410 18284
rect 20916 18281 20944 18312
rect 20625 18275 20683 18281
rect 20625 18272 20637 18275
rect 20404 18244 20637 18272
rect 20404 18232 20410 18244
rect 20625 18241 20637 18244
rect 20671 18241 20683 18275
rect 20625 18235 20683 18241
rect 20901 18275 20959 18281
rect 20901 18241 20913 18275
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 18380 18176 18736 18204
rect 18380 18164 18386 18176
rect 21634 18164 21640 18216
rect 21692 18164 21698 18216
rect 13078 18028 13084 18080
rect 13136 18028 13142 18080
rect 15194 18028 15200 18080
rect 15252 18028 15258 18080
rect 15930 18028 15936 18080
rect 15988 18028 15994 18080
rect 18417 18071 18475 18077
rect 18417 18037 18429 18071
rect 18463 18068 18475 18071
rect 18690 18068 18696 18080
rect 18463 18040 18696 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 18690 18028 18696 18040
rect 18748 18028 18754 18080
rect 1104 17978 35248 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 35248 17978
rect 1104 17904 35248 17926
rect 14826 17824 14832 17876
rect 14884 17824 14890 17876
rect 15930 17824 15936 17876
rect 15988 17824 15994 17876
rect 16301 17867 16359 17873
rect 16301 17833 16313 17867
rect 16347 17864 16359 17867
rect 16482 17864 16488 17876
rect 16347 17836 16488 17864
rect 16347 17833 16359 17836
rect 16301 17827 16359 17833
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 16574 17824 16580 17876
rect 16632 17824 16638 17876
rect 19797 17867 19855 17873
rect 19797 17864 19809 17867
rect 18800 17836 19809 17864
rect 15746 17756 15752 17808
rect 15804 17756 15810 17808
rect 16592 17796 16620 17824
rect 15856 17768 16436 17796
rect 16592 17768 16804 17796
rect 10781 17731 10839 17737
rect 10781 17697 10793 17731
rect 10827 17728 10839 17731
rect 10827 17700 12112 17728
rect 10827 17697 10839 17700
rect 10781 17691 10839 17697
rect 12084 17672 12112 17700
rect 13078 17688 13084 17740
rect 13136 17728 13142 17740
rect 15013 17731 15071 17737
rect 13136 17700 13768 17728
rect 13136 17688 13142 17700
rect 10321 17663 10379 17669
rect 10321 17629 10333 17663
rect 10367 17629 10379 17663
rect 10321 17623 10379 17629
rect 10336 17592 10364 17623
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 10468 17632 10609 17660
rect 10468 17620 10474 17632
rect 10597 17629 10609 17632
rect 10643 17660 10655 17663
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 10643 17632 10885 17660
rect 10643 17629 10655 17632
rect 10597 17623 10655 17629
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 11330 17660 11336 17672
rect 10873 17623 10931 17629
rect 10980 17632 11336 17660
rect 10980 17592 11008 17632
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 11514 17620 11520 17672
rect 11572 17620 11578 17672
rect 12066 17620 12072 17672
rect 12124 17620 12130 17672
rect 12345 17663 12403 17669
rect 12345 17629 12357 17663
rect 12391 17629 12403 17663
rect 12345 17623 12403 17629
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12986 17660 12992 17672
rect 12575 17632 12992 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 10336 17564 11008 17592
rect 11054 17552 11060 17604
rect 11112 17592 11118 17604
rect 11425 17595 11483 17601
rect 11425 17592 11437 17595
rect 11112 17564 11437 17592
rect 11112 17552 11118 17564
rect 11425 17561 11437 17564
rect 11471 17592 11483 17595
rect 12158 17592 12164 17604
rect 11471 17564 12164 17592
rect 11471 17561 11483 17564
rect 11425 17555 11483 17561
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 10413 17527 10471 17533
rect 10413 17493 10425 17527
rect 10459 17524 10471 17527
rect 10686 17524 10692 17536
rect 10459 17496 10692 17524
rect 10459 17493 10471 17496
rect 10413 17487 10471 17493
rect 10686 17484 10692 17496
rect 10744 17524 10750 17536
rect 11514 17524 11520 17536
rect 10744 17496 11520 17524
rect 10744 17484 10750 17496
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 12360 17524 12388 17623
rect 12986 17620 12992 17632
rect 13044 17660 13050 17672
rect 13740 17669 13768 17700
rect 15013 17697 15025 17731
rect 15059 17728 15071 17731
rect 15473 17731 15531 17737
rect 15059 17700 15332 17728
rect 15059 17697 15071 17700
rect 15013 17691 15071 17697
rect 15304 17672 15332 17700
rect 15473 17697 15485 17731
rect 15519 17728 15531 17731
rect 15764 17728 15792 17756
rect 15519 17700 15792 17728
rect 15519 17697 15531 17700
rect 15473 17691 15531 17697
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 13044 17632 13185 17660
rect 13044 17620 13050 17632
rect 13173 17629 13185 17632
rect 13219 17660 13231 17663
rect 13449 17663 13507 17669
rect 13449 17660 13461 17663
rect 13219 17632 13461 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 13449 17629 13461 17632
rect 13495 17629 13507 17663
rect 13449 17623 13507 17629
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 15105 17663 15163 17669
rect 15105 17629 15117 17663
rect 15151 17660 15163 17663
rect 15194 17660 15200 17672
rect 15151 17632 15200 17660
rect 15151 17629 15163 17632
rect 15105 17623 15163 17629
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 15286 17620 15292 17672
rect 15344 17620 15350 17672
rect 15749 17663 15807 17669
rect 15749 17629 15761 17663
rect 15795 17660 15807 17663
rect 15856 17660 15884 17768
rect 16408 17740 16436 17768
rect 15795 17632 15884 17660
rect 15948 17700 16252 17728
rect 15795 17629 15807 17632
rect 15749 17623 15807 17629
rect 12713 17595 12771 17601
rect 12713 17561 12725 17595
rect 12759 17592 12771 17595
rect 13541 17595 13599 17601
rect 13541 17592 13553 17595
rect 12759 17564 13553 17592
rect 12759 17561 12771 17564
rect 12713 17555 12771 17561
rect 13188 17536 13216 17564
rect 13541 17561 13553 17564
rect 13587 17561 13599 17595
rect 13541 17555 13599 17561
rect 13909 17595 13967 17601
rect 13909 17561 13921 17595
rect 13955 17592 13967 17595
rect 15948 17592 15976 17700
rect 16025 17663 16083 17669
rect 16025 17629 16037 17663
rect 16071 17629 16083 17663
rect 16025 17623 16083 17629
rect 13955 17564 15976 17592
rect 13955 17561 13967 17564
rect 13909 17555 13967 17561
rect 16040 17536 16068 17623
rect 16224 17592 16252 17700
rect 16390 17688 16396 17740
rect 16448 17728 16454 17740
rect 16776 17737 16804 17768
rect 17696 17768 18552 17796
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16448 17700 16681 17728
rect 16448 17688 16454 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 16761 17731 16819 17737
rect 16761 17697 16773 17731
rect 16807 17728 16819 17731
rect 16850 17728 16856 17740
rect 16807 17700 16856 17728
rect 16807 17697 16819 17700
rect 16761 17691 16819 17697
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 17696 17737 17724 17768
rect 18524 17740 18552 17768
rect 16945 17731 17003 17737
rect 16945 17697 16957 17731
rect 16991 17697 17003 17731
rect 16945 17691 17003 17697
rect 17681 17731 17739 17737
rect 17681 17697 17693 17731
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 16298 17620 16304 17672
rect 16356 17660 16362 17672
rect 16485 17663 16543 17669
rect 16485 17660 16497 17663
rect 16356 17632 16497 17660
rect 16356 17620 16362 17632
rect 16485 17629 16497 17632
rect 16531 17629 16543 17663
rect 16485 17623 16543 17629
rect 16574 17620 16580 17672
rect 16632 17620 16638 17672
rect 16960 17660 16988 17691
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18049 17731 18107 17737
rect 18049 17728 18061 17731
rect 18012 17700 18061 17728
rect 18012 17688 18018 17700
rect 18049 17697 18061 17700
rect 18095 17697 18107 17731
rect 18049 17691 18107 17697
rect 18506 17688 18512 17740
rect 18564 17688 18570 17740
rect 17034 17660 17040 17672
rect 16960 17632 17040 17660
rect 17034 17620 17040 17632
rect 17092 17620 17098 17672
rect 17126 17620 17132 17672
rect 17184 17660 17190 17672
rect 17313 17663 17371 17669
rect 17313 17660 17325 17663
rect 17184 17632 17325 17660
rect 17184 17620 17190 17632
rect 17313 17629 17325 17632
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 18141 17663 18199 17669
rect 18141 17660 18153 17663
rect 17543 17632 18153 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 18141 17629 18153 17632
rect 18187 17660 18199 17663
rect 18322 17660 18328 17672
rect 18187 17632 18328 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18322 17620 18328 17632
rect 18380 17620 18386 17672
rect 18414 17620 18420 17672
rect 18472 17620 18478 17672
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 18800 17669 18828 17836
rect 19797 17833 19809 17836
rect 19843 17833 19855 17867
rect 19797 17827 19855 17833
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 18932 17700 19840 17728
rect 18932 17688 18938 17700
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 18748 17632 18797 17660
rect 18748 17620 18754 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 18966 17620 18972 17672
rect 19024 17660 19030 17672
rect 19812 17669 19840 17700
rect 19337 17663 19395 17669
rect 19337 17660 19349 17663
rect 19024 17632 19349 17660
rect 19024 17620 19030 17632
rect 19337 17629 19349 17632
rect 19383 17629 19395 17663
rect 19337 17623 19395 17629
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19797 17663 19855 17669
rect 19797 17629 19809 17663
rect 19843 17629 19855 17663
rect 19797 17623 19855 17629
rect 18509 17595 18567 17601
rect 18509 17592 18521 17595
rect 16224 17564 18521 17592
rect 18509 17561 18521 17564
rect 18555 17592 18567 17595
rect 19444 17592 19472 17623
rect 18555 17564 19472 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 12526 17524 12532 17536
rect 12360 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13170 17484 13176 17536
rect 13228 17484 13234 17536
rect 13354 17484 13360 17536
rect 13412 17484 13418 17536
rect 16022 17484 16028 17536
rect 16080 17484 16086 17536
rect 16666 17484 16672 17536
rect 16724 17524 16730 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 16724 17496 17141 17524
rect 16724 17484 16730 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 18322 17484 18328 17536
rect 18380 17484 18386 17536
rect 18414 17484 18420 17536
rect 18472 17524 18478 17536
rect 18966 17524 18972 17536
rect 18472 17496 18972 17524
rect 18472 17484 18478 17496
rect 18966 17484 18972 17496
rect 19024 17484 19030 17536
rect 19058 17484 19064 17536
rect 19116 17484 19122 17536
rect 19978 17484 19984 17536
rect 20036 17484 20042 17536
rect 1104 17434 35236 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 35236 17434
rect 1104 17360 35236 17382
rect 10505 17323 10563 17329
rect 10505 17289 10517 17323
rect 10551 17320 10563 17323
rect 11330 17320 11336 17332
rect 10551 17292 11336 17320
rect 10551 17289 10563 17292
rect 10505 17283 10563 17289
rect 11330 17280 11336 17292
rect 11388 17280 11394 17332
rect 12066 17280 12072 17332
rect 12124 17320 12130 17332
rect 12124 17292 12296 17320
rect 12124 17280 12130 17292
rect 10689 17255 10747 17261
rect 10689 17252 10701 17255
rect 9876 17224 10701 17252
rect 9876 17193 9904 17224
rect 10689 17221 10701 17224
rect 10735 17221 10747 17255
rect 10689 17215 10747 17221
rect 12158 17212 12164 17264
rect 12216 17212 12222 17264
rect 12268 17261 12296 17292
rect 12986 17280 12992 17332
rect 13044 17280 13050 17332
rect 13078 17280 13084 17332
rect 13136 17280 13142 17332
rect 15286 17280 15292 17332
rect 15344 17320 15350 17332
rect 15581 17323 15639 17329
rect 15581 17320 15593 17323
rect 15344 17292 15593 17320
rect 15344 17280 15350 17292
rect 15581 17289 15593 17292
rect 15627 17289 15639 17323
rect 15581 17283 15639 17289
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17289 15807 17323
rect 15749 17283 15807 17289
rect 12253 17255 12311 17261
rect 12253 17221 12265 17255
rect 12299 17221 12311 17255
rect 12253 17215 12311 17221
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 9950 17144 9956 17196
rect 10008 17184 10014 17196
rect 10597 17187 10655 17193
rect 10597 17184 10609 17187
rect 10008 17156 10609 17184
rect 10008 17144 10014 17156
rect 10597 17153 10609 17156
rect 10643 17153 10655 17187
rect 10597 17147 10655 17153
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 12176 17184 12204 17212
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12176 17156 12449 17184
rect 10781 17147 10839 17153
rect 12437 17153 12449 17156
rect 12483 17153 12495 17187
rect 12437 17147 12495 17153
rect 9674 17076 9680 17128
rect 9732 17076 9738 17128
rect 10042 17076 10048 17128
rect 10100 17116 10106 17128
rect 10796 17116 10824 17147
rect 12526 17144 12532 17196
rect 12584 17144 12590 17196
rect 13004 17193 13032 17280
rect 13096 17252 13124 17280
rect 13096 17224 13308 17252
rect 12989 17187 13047 17193
rect 12989 17153 13001 17187
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13170 17144 13176 17196
rect 13228 17144 13234 17196
rect 13280 17193 13308 17224
rect 15194 17212 15200 17264
rect 15252 17252 15258 17264
rect 15378 17252 15384 17264
rect 15252 17224 15384 17252
rect 15252 17212 15258 17224
rect 15378 17212 15384 17224
rect 15436 17212 15442 17264
rect 13265 17187 13323 17193
rect 13265 17153 13277 17187
rect 13311 17153 13323 17187
rect 15764 17184 15792 17283
rect 15930 17280 15936 17332
rect 15988 17280 15994 17332
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 16850 17320 16856 17332
rect 16356 17292 16856 17320
rect 16356 17280 16362 17292
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 17034 17280 17040 17332
rect 17092 17320 17098 17332
rect 17092 17292 17264 17320
rect 17092 17280 17098 17292
rect 15948 17252 15976 17280
rect 15948 17224 16436 17252
rect 16022 17184 16028 17196
rect 15764 17156 16028 17184
rect 13265 17147 13323 17153
rect 16022 17144 16028 17156
rect 16080 17184 16086 17196
rect 16408 17193 16436 17224
rect 16666 17212 16672 17264
rect 16724 17252 16730 17264
rect 17236 17261 17264 17292
rect 18230 17280 18236 17332
rect 18288 17320 18294 17332
rect 18709 17323 18767 17329
rect 18709 17320 18721 17323
rect 18288 17292 18721 17320
rect 18288 17280 18294 17292
rect 18709 17289 18721 17292
rect 18755 17289 18767 17323
rect 18709 17283 18767 17289
rect 18874 17280 18880 17332
rect 18932 17280 18938 17332
rect 19058 17280 19064 17332
rect 19116 17280 19122 17332
rect 17129 17255 17187 17261
rect 17129 17252 17141 17255
rect 16724 17224 17141 17252
rect 16724 17212 16730 17224
rect 17129 17221 17141 17224
rect 17175 17221 17187 17255
rect 17129 17215 17187 17221
rect 17221 17255 17279 17261
rect 17221 17221 17233 17255
rect 17267 17221 17279 17255
rect 17221 17215 17279 17221
rect 16209 17187 16267 17193
rect 16209 17184 16221 17187
rect 16080 17156 16221 17184
rect 16080 17144 16086 17156
rect 16209 17153 16221 17156
rect 16255 17153 16267 17187
rect 16209 17147 16267 17153
rect 16393 17187 16451 17193
rect 16393 17153 16405 17187
rect 16439 17153 16451 17187
rect 16393 17147 16451 17153
rect 16482 17144 16488 17196
rect 16540 17184 16546 17196
rect 16761 17187 16819 17193
rect 16761 17184 16773 17187
rect 16540 17156 16773 17184
rect 16540 17144 16546 17156
rect 16761 17153 16773 17156
rect 16807 17153 16819 17187
rect 16761 17147 16819 17153
rect 16850 17144 16856 17196
rect 16908 17144 16914 17196
rect 16942 17144 16948 17196
rect 17000 17144 17006 17196
rect 17144 17184 17172 17215
rect 17954 17212 17960 17264
rect 18012 17252 18018 17264
rect 18509 17255 18567 17261
rect 18509 17252 18521 17255
rect 18012 17224 18521 17252
rect 18012 17212 18018 17224
rect 18509 17221 18521 17224
rect 18555 17221 18567 17255
rect 19076 17252 19104 17280
rect 20625 17255 20683 17261
rect 20625 17252 20637 17255
rect 19076 17224 20637 17252
rect 18509 17215 18567 17221
rect 20625 17221 20637 17224
rect 20671 17252 20683 17255
rect 21821 17255 21879 17261
rect 21821 17252 21833 17255
rect 20671 17224 21833 17252
rect 20671 17221 20683 17224
rect 20625 17215 20683 17221
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 17144 17156 17417 17184
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17405 17147 17463 17153
rect 17497 17187 17555 17193
rect 17497 17153 17509 17187
rect 17543 17153 17555 17187
rect 17497 17147 17555 17153
rect 10100 17088 10824 17116
rect 10100 17076 10106 17088
rect 12529 17051 12587 17057
rect 12529 17017 12541 17051
rect 12575 17048 12587 17051
rect 13188 17048 13216 17144
rect 17126 17076 17132 17128
rect 17184 17116 17190 17128
rect 17512 17116 17540 17147
rect 19978 17144 19984 17196
rect 20036 17184 20042 17196
rect 20809 17187 20867 17193
rect 20809 17184 20821 17187
rect 20036 17156 20821 17184
rect 20036 17144 20042 17156
rect 20809 17153 20821 17156
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 17184 17088 17540 17116
rect 20824 17116 20852 17147
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 21008 17193 21036 17224
rect 21821 17221 21833 17224
rect 21867 17221 21879 17255
rect 21821 17215 21879 17221
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 21100 17116 21128 17147
rect 21174 17144 21180 17196
rect 21232 17184 21238 17196
rect 21269 17187 21327 17193
rect 21269 17184 21281 17187
rect 21232 17156 21281 17184
rect 21232 17144 21238 17156
rect 21269 17153 21281 17156
rect 21315 17184 21327 17187
rect 22373 17187 22431 17193
rect 22373 17184 22385 17187
rect 21315 17156 22385 17184
rect 21315 17153 21327 17156
rect 21269 17147 21327 17153
rect 22373 17153 22385 17156
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 22465 17119 22523 17125
rect 22465 17116 22477 17119
rect 20824 17088 22477 17116
rect 17184 17076 17190 17088
rect 22465 17085 22477 17088
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 12575 17020 13216 17048
rect 13265 17051 13323 17057
rect 12575 17017 12587 17020
rect 12529 17011 12587 17017
rect 13265 17017 13277 17051
rect 13311 17048 13323 17051
rect 18414 17048 18420 17060
rect 13311 17020 18420 17048
rect 13311 17017 13323 17020
rect 13265 17011 13323 17017
rect 18414 17008 18420 17020
rect 18472 17008 18478 17060
rect 22094 17008 22100 17060
rect 22152 17008 22158 17060
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 15746 16980 15752 16992
rect 15611 16952 15752 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 15746 16940 15752 16952
rect 15804 16940 15810 16992
rect 16393 16983 16451 16989
rect 16393 16949 16405 16983
rect 16439 16980 16451 16983
rect 16574 16980 16580 16992
rect 16439 16952 16580 16980
rect 16439 16949 16451 16952
rect 16393 16943 16451 16949
rect 16574 16940 16580 16952
rect 16632 16980 16638 16992
rect 16942 16980 16948 16992
rect 16632 16952 16948 16980
rect 16632 16940 16638 16952
rect 16942 16940 16948 16952
rect 17000 16940 17006 16992
rect 17497 16983 17555 16989
rect 17497 16949 17509 16983
rect 17543 16980 17555 16983
rect 18506 16980 18512 16992
rect 17543 16952 18512 16980
rect 17543 16949 17555 16952
rect 17497 16943 17555 16949
rect 18506 16940 18512 16952
rect 18564 16980 18570 16992
rect 18693 16983 18751 16989
rect 18693 16980 18705 16983
rect 18564 16952 18705 16980
rect 18564 16940 18570 16952
rect 18693 16949 18705 16952
rect 18739 16949 18751 16983
rect 18693 16943 18751 16949
rect 20898 16940 20904 16992
rect 20956 16940 20962 16992
rect 21174 16940 21180 16992
rect 21232 16980 21238 16992
rect 21453 16983 21511 16989
rect 21453 16980 21465 16983
rect 21232 16952 21465 16980
rect 21232 16940 21238 16952
rect 21453 16949 21465 16952
rect 21499 16949 21511 16983
rect 21453 16943 21511 16949
rect 1104 16890 35248 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 35248 16890
rect 1104 16816 35248 16838
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 10410 16776 10416 16788
rect 9723 16748 10416 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 10410 16736 10416 16748
rect 10468 16736 10474 16788
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 15746 16776 15752 16788
rect 14875 16748 15752 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16708 9551 16711
rect 9539 16680 9628 16708
rect 9539 16677 9551 16680
rect 9493 16671 9551 16677
rect 9214 16600 9220 16652
rect 9272 16600 9278 16652
rect 9600 16649 9628 16680
rect 14734 16668 14740 16720
rect 14792 16708 14798 16720
rect 17678 16708 17684 16720
rect 14792 16680 15332 16708
rect 14792 16668 14798 16680
rect 9585 16643 9643 16649
rect 9585 16609 9597 16643
rect 9631 16609 9643 16643
rect 9585 16603 9643 16609
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9815 16612 10057 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 10045 16609 10057 16612
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 13740 16612 15238 16640
rect 9125 16575 9183 16581
rect 9125 16541 9137 16575
rect 9171 16572 9183 16575
rect 9861 16575 9919 16581
rect 9171 16544 9812 16572
rect 9171 16541 9183 16544
rect 9125 16535 9183 16541
rect 9784 16516 9812 16544
rect 9861 16541 9873 16575
rect 9907 16541 9919 16575
rect 9861 16535 9919 16541
rect 9766 16464 9772 16516
rect 9824 16464 9830 16516
rect 9876 16448 9904 16535
rect 9950 16532 9956 16584
rect 10008 16532 10014 16584
rect 10137 16575 10195 16581
rect 10137 16572 10149 16575
rect 10060 16544 10149 16572
rect 10060 16448 10088 16544
rect 10137 16541 10149 16544
rect 10183 16541 10195 16575
rect 10137 16535 10195 16541
rect 13740 16516 13768 16612
rect 14553 16575 14611 16581
rect 14553 16572 14565 16575
rect 14476 16544 14565 16572
rect 13722 16464 13728 16516
rect 13780 16464 13786 16516
rect 14476 16448 14504 16544
rect 14553 16541 14565 16544
rect 14599 16541 14611 16575
rect 14553 16535 14611 16541
rect 14734 16532 14740 16584
rect 14792 16572 14798 16584
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14792 16544 14933 16572
rect 14792 16532 14798 16544
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15105 16575 15163 16581
rect 15105 16541 15117 16575
rect 15151 16541 15163 16575
rect 15105 16535 15163 16541
rect 15119 16504 15147 16535
rect 14660 16476 15147 16504
rect 15210 16504 15238 16612
rect 15304 16581 15332 16680
rect 15396 16680 17684 16708
rect 15396 16652 15424 16680
rect 17678 16668 17684 16680
rect 17736 16668 17742 16720
rect 22094 16668 22100 16720
rect 22152 16708 22158 16720
rect 22152 16680 22692 16708
rect 22152 16668 22158 16680
rect 15378 16600 15384 16652
rect 15436 16600 15442 16652
rect 16298 16600 16304 16652
rect 16356 16640 16362 16652
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16356 16612 16865 16640
rect 16356 16600 16362 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 19242 16640 19248 16652
rect 17819 16612 19248 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 19242 16600 19248 16612
rect 19300 16600 19306 16652
rect 22664 16649 22692 16680
rect 22649 16643 22707 16649
rect 22649 16609 22661 16643
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 15289 16575 15347 16581
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 16942 16532 16948 16584
rect 17000 16532 17006 16584
rect 20990 16532 20996 16584
rect 21048 16532 21054 16584
rect 21100 16504 21128 16558
rect 22094 16532 22100 16584
rect 22152 16532 22158 16584
rect 22465 16575 22523 16581
rect 22465 16541 22477 16575
rect 22511 16541 22523 16575
rect 22465 16535 22523 16541
rect 21358 16504 21364 16516
rect 15210 16476 21364 16504
rect 14660 16448 14688 16476
rect 21358 16464 21364 16476
rect 21416 16464 21422 16516
rect 22002 16464 22008 16516
rect 22060 16504 22066 16516
rect 22480 16504 22508 16535
rect 22060 16476 22508 16504
rect 22060 16464 22066 16476
rect 9858 16396 9864 16448
rect 9916 16396 9922 16448
rect 10042 16396 10048 16448
rect 10100 16396 10106 16448
rect 14458 16396 14464 16448
rect 14516 16396 14522 16448
rect 14642 16396 14648 16448
rect 14700 16396 14706 16448
rect 14737 16439 14795 16445
rect 14737 16405 14749 16439
rect 14783 16436 14795 16439
rect 14826 16436 14832 16448
rect 14783 16408 14832 16436
rect 14783 16405 14795 16408
rect 14737 16399 14795 16405
rect 14826 16396 14832 16408
rect 14884 16396 14890 16448
rect 15289 16439 15347 16445
rect 15289 16405 15301 16439
rect 15335 16436 15347 16439
rect 15470 16436 15476 16448
rect 15335 16408 15476 16436
rect 15335 16405 15347 16408
rect 15289 16399 15347 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 22465 16439 22523 16445
rect 22465 16405 22477 16439
rect 22511 16436 22523 16439
rect 26050 16436 26056 16448
rect 22511 16408 26056 16436
rect 22511 16405 22523 16408
rect 22465 16399 22523 16405
rect 26050 16396 26056 16408
rect 26108 16396 26114 16448
rect 1104 16346 35236 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 35236 16346
rect 1104 16272 35236 16294
rect 11333 16235 11391 16241
rect 10704 16204 11192 16232
rect 10704 16108 10732 16204
rect 10781 16167 10839 16173
rect 10781 16133 10793 16167
rect 10827 16164 10839 16167
rect 11054 16164 11060 16176
rect 10827 16136 11060 16164
rect 10827 16133 10839 16136
rect 10781 16127 10839 16133
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 11164 16173 11192 16204
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11379 16204 14228 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11149 16167 11207 16173
rect 11149 16133 11161 16167
rect 11195 16133 11207 16167
rect 11149 16127 11207 16133
rect 13722 16124 13728 16176
rect 13780 16124 13786 16176
rect 14200 16164 14228 16204
rect 14274 16192 14280 16244
rect 14332 16192 14338 16244
rect 14645 16235 14703 16241
rect 14645 16201 14657 16235
rect 14691 16232 14703 16235
rect 14826 16232 14832 16244
rect 14691 16204 14832 16232
rect 14691 16201 14703 16204
rect 14645 16195 14703 16201
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 19337 16235 19395 16241
rect 14936 16204 18644 16232
rect 14936 16164 14964 16204
rect 14200 16136 14964 16164
rect 15013 16167 15071 16173
rect 15013 16133 15025 16167
rect 15059 16164 15071 16167
rect 15289 16167 15347 16173
rect 15289 16164 15301 16167
rect 15059 16136 15301 16164
rect 15059 16133 15071 16136
rect 15013 16127 15071 16133
rect 15289 16133 15301 16136
rect 15335 16133 15347 16167
rect 15289 16127 15347 16133
rect 15381 16167 15439 16173
rect 15381 16133 15393 16167
rect 15427 16164 15439 16167
rect 15749 16167 15807 16173
rect 15749 16164 15761 16167
rect 15427 16136 15761 16164
rect 15427 16133 15439 16136
rect 15381 16127 15439 16133
rect 15749 16133 15761 16136
rect 15795 16133 15807 16167
rect 15749 16127 15807 16133
rect 13360 16108 13412 16114
rect 10318 16056 10324 16108
rect 10376 16096 10382 16108
rect 10413 16099 10471 16105
rect 10413 16096 10425 16099
rect 10376 16068 10425 16096
rect 10376 16056 10382 16068
rect 10413 16065 10425 16068
rect 10459 16065 10471 16099
rect 10413 16059 10471 16065
rect 10686 16056 10692 16108
rect 10744 16056 10750 16108
rect 10965 16099 11023 16105
rect 10965 16065 10977 16099
rect 11011 16065 11023 16099
rect 10965 16059 11023 16065
rect 9766 15988 9772 16040
rect 9824 16028 9830 16040
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 9824 16000 10241 16028
rect 9824 15988 9830 16000
rect 10229 15997 10241 16000
rect 10275 15997 10287 16031
rect 10980 16028 11008 16059
rect 15105 16099 15163 16105
rect 15105 16096 15117 16099
rect 13360 16050 13412 16056
rect 14200 16068 15117 16096
rect 10980 16000 11468 16028
rect 10229 15991 10287 15997
rect 11440 15904 11468 16000
rect 12894 15988 12900 16040
rect 12952 15988 12958 16040
rect 13814 15988 13820 16040
rect 13872 15988 13878 16040
rect 14200 15969 14228 16068
rect 15105 16065 15117 16068
rect 15151 16065 15163 16099
rect 15105 16059 15163 16065
rect 15470 16056 15476 16108
rect 15528 16056 15534 16108
rect 15930 16056 15936 16108
rect 15988 16056 15994 16108
rect 16022 16056 16028 16108
rect 16080 16096 16086 16108
rect 16117 16099 16175 16105
rect 16117 16096 16129 16099
rect 16080 16068 16129 16096
rect 16080 16056 16086 16068
rect 16117 16065 16129 16068
rect 16163 16065 16175 16099
rect 16117 16059 16175 16065
rect 17954 16056 17960 16108
rect 18012 16096 18018 16108
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18012 16068 18521 16096
rect 18012 16056 18018 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18509 16059 18567 16065
rect 14369 16031 14427 16037
rect 14369 15997 14381 16031
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 14461 16031 14519 16037
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 14642 16028 14648 16040
rect 14507 16000 14648 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 14185 15963 14243 15969
rect 14185 15929 14197 15963
rect 14231 15929 14243 15963
rect 14384 15960 14412 15991
rect 14642 15988 14648 16000
rect 14700 15988 14706 16040
rect 14734 15988 14740 16040
rect 14792 15988 14798 16040
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 16028 14887 16031
rect 15010 16028 15016 16040
rect 14875 16000 15016 16028
rect 14875 15997 14887 16000
rect 14829 15991 14887 15997
rect 15010 15988 15016 16000
rect 15068 15988 15074 16040
rect 17402 15988 17408 16040
rect 17460 15988 17466 16040
rect 18049 16031 18107 16037
rect 18049 15997 18061 16031
rect 18095 16028 18107 16031
rect 18322 16028 18328 16040
rect 18095 16000 18328 16028
rect 18095 15997 18107 16000
rect 18049 15991 18107 15997
rect 18322 15988 18328 16000
rect 18380 16028 18386 16040
rect 18417 16031 18475 16037
rect 18417 16028 18429 16031
rect 18380 16000 18429 16028
rect 18380 15988 18386 16000
rect 18417 15997 18429 16000
rect 18463 15997 18475 16031
rect 18616 16028 18644 16204
rect 19337 16201 19349 16235
rect 19383 16232 19395 16235
rect 20990 16232 20996 16244
rect 19383 16204 20996 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 20990 16192 20996 16204
rect 21048 16232 21054 16244
rect 21361 16235 21419 16241
rect 21048 16204 21312 16232
rect 21048 16192 21054 16204
rect 21085 16167 21143 16173
rect 21085 16164 21097 16167
rect 20640 16136 21097 16164
rect 19242 16056 19248 16108
rect 19300 16096 19306 16108
rect 19794 16096 19800 16108
rect 19300 16068 19800 16096
rect 19300 16056 19306 16068
rect 19794 16056 19800 16068
rect 19852 16056 19858 16108
rect 20257 16099 20315 16105
rect 20257 16065 20269 16099
rect 20303 16065 20315 16099
rect 20257 16059 20315 16065
rect 19705 16031 19763 16037
rect 19705 16028 19717 16031
rect 18616 16000 19717 16028
rect 18417 15991 18475 15997
rect 19705 15997 19717 16000
rect 19751 16028 19763 16031
rect 19751 16000 20024 16028
rect 19751 15997 19763 16000
rect 19705 15991 19763 15997
rect 14660 15960 14688 15988
rect 15657 15963 15715 15969
rect 14384 15932 14504 15960
rect 14660 15932 14964 15960
rect 14185 15923 14243 15929
rect 10689 15895 10747 15901
rect 10689 15861 10701 15895
rect 10735 15892 10747 15895
rect 11330 15892 11336 15904
rect 10735 15864 11336 15892
rect 10735 15861 10747 15864
rect 10689 15855 10747 15861
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 11422 15852 11428 15904
rect 11480 15852 11486 15904
rect 14200 15892 14228 15923
rect 14476 15904 14504 15932
rect 14936 15904 14964 15932
rect 15657 15929 15669 15963
rect 15703 15960 15715 15963
rect 16850 15960 16856 15972
rect 15703 15932 16856 15960
rect 15703 15929 15715 15932
rect 15657 15923 15715 15929
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 17681 15963 17739 15969
rect 17681 15929 17693 15963
rect 17727 15960 17739 15963
rect 19996 15960 20024 16000
rect 20070 15988 20076 16040
rect 20128 15988 20134 16040
rect 20272 16028 20300 16059
rect 20438 16056 20444 16108
rect 20496 16096 20502 16108
rect 20640 16105 20668 16136
rect 21085 16133 21097 16136
rect 21131 16133 21143 16167
rect 21085 16127 21143 16133
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20496 16068 20545 16096
rect 20496 16056 20502 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 20714 16056 20720 16108
rect 20772 16056 20778 16108
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 20990 16096 20996 16108
rect 20947 16068 20996 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21284 16105 21312 16204
rect 21361 16201 21373 16235
rect 21407 16232 21419 16235
rect 22094 16232 22100 16244
rect 21407 16204 22100 16232
rect 21407 16201 21419 16204
rect 21361 16195 21419 16201
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 24121 16235 24179 16241
rect 24121 16201 24133 16235
rect 24167 16232 24179 16235
rect 24167 16204 26556 16232
rect 24167 16201 24179 16204
rect 24121 16195 24179 16201
rect 22002 16124 22008 16176
rect 22060 16164 22066 16176
rect 22060 16136 22232 16164
rect 22060 16124 22066 16136
rect 21177 16099 21235 16105
rect 21177 16065 21189 16099
rect 21223 16065 21235 16099
rect 21177 16059 21235 16065
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 20809 16031 20867 16037
rect 20809 16028 20821 16031
rect 20272 16000 20821 16028
rect 20809 15997 20821 16000
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 20714 15960 20720 15972
rect 17727 15932 19932 15960
rect 19996 15932 20720 15960
rect 17727 15929 17739 15932
rect 17681 15923 17739 15929
rect 14366 15892 14372 15904
rect 14200 15864 14372 15892
rect 14366 15852 14372 15864
rect 14424 15852 14430 15904
rect 14458 15852 14464 15904
rect 14516 15852 14522 15904
rect 14918 15852 14924 15904
rect 14976 15852 14982 15904
rect 19426 15852 19432 15904
rect 19484 15852 19490 15904
rect 19904 15892 19932 15932
rect 20714 15920 20720 15932
rect 20772 15960 20778 15972
rect 21192 15960 21220 16059
rect 21358 16056 21364 16108
rect 21416 16096 21422 16108
rect 22204 16105 22232 16136
rect 22480 16136 24716 16164
rect 21453 16099 21511 16105
rect 21453 16096 21465 16099
rect 21416 16068 21465 16096
rect 21416 16056 21422 16068
rect 21453 16065 21465 16068
rect 21499 16065 21511 16099
rect 21453 16059 21511 16065
rect 22189 16099 22247 16105
rect 22189 16065 22201 16099
rect 22235 16065 22247 16099
rect 22189 16059 22247 16065
rect 22094 15988 22100 16040
rect 22152 15988 22158 16040
rect 20772 15932 21220 15960
rect 20772 15920 20778 15932
rect 22480 15892 22508 16136
rect 24688 16108 24716 16136
rect 26050 16124 26056 16176
rect 26108 16124 26114 16176
rect 23290 16056 23296 16108
rect 23348 16096 23354 16108
rect 23753 16099 23811 16105
rect 23753 16096 23765 16099
rect 23348 16068 23765 16096
rect 23348 16056 23354 16068
rect 23753 16065 23765 16068
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 23846 16099 23904 16105
rect 23846 16065 23858 16099
rect 23892 16065 23904 16099
rect 23846 16059 23904 16065
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 16028 23443 16031
rect 23860 16028 23888 16059
rect 24670 16056 24676 16108
rect 24728 16056 24734 16108
rect 24854 16056 24860 16108
rect 24912 16056 24918 16108
rect 26528 16096 26556 16204
rect 26970 16124 26976 16176
rect 27028 16164 27034 16176
rect 27028 16136 28212 16164
rect 27028 16124 27034 16136
rect 27065 16099 27123 16105
rect 27065 16096 27077 16099
rect 26528 16068 27077 16096
rect 27065 16065 27077 16068
rect 27111 16065 27123 16099
rect 27172 16082 27200 16136
rect 28184 16105 28212 16136
rect 28169 16099 28227 16105
rect 27065 16059 27123 16065
rect 28169 16065 28181 16099
rect 28215 16065 28227 16099
rect 28169 16059 28227 16065
rect 28353 16099 28411 16105
rect 28353 16065 28365 16099
rect 28399 16065 28411 16099
rect 28353 16059 28411 16065
rect 23431 16000 23888 16028
rect 23431 15997 23443 16000
rect 23385 15991 23443 15997
rect 19904 15864 22508 15892
rect 22557 15895 22615 15901
rect 22557 15861 22569 15895
rect 22603 15892 22615 15895
rect 23400 15892 23428 15991
rect 25682 15988 25688 16040
rect 25740 16028 25746 16040
rect 25740 16000 26372 16028
rect 25740 15988 25746 16000
rect 23661 15963 23719 15969
rect 23661 15929 23673 15963
rect 23707 15960 23719 15963
rect 24302 15960 24308 15972
rect 23707 15932 24308 15960
rect 23707 15929 23719 15932
rect 23661 15923 23719 15929
rect 24302 15920 24308 15932
rect 24360 15920 24366 15972
rect 26344 15969 26372 16000
rect 26329 15963 26387 15969
rect 26329 15929 26341 15963
rect 26375 15929 26387 15963
rect 27080 15960 27108 16059
rect 28074 15988 28080 16040
rect 28132 15988 28138 16040
rect 28368 15960 28396 16059
rect 27080 15932 28396 15960
rect 26329 15923 26387 15929
rect 22603 15864 23428 15892
rect 22603 15861 22615 15864
rect 22557 15855 22615 15861
rect 26510 15852 26516 15904
rect 26568 15852 26574 15904
rect 28166 15852 28172 15904
rect 28224 15852 28230 15904
rect 1104 15802 35248 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 35248 15802
rect 1104 15728 35248 15750
rect 9674 15648 9680 15700
rect 9732 15648 9738 15700
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10873 15691 10931 15697
rect 10873 15688 10885 15691
rect 10284 15660 10885 15688
rect 10284 15648 10290 15660
rect 10873 15657 10885 15660
rect 10919 15657 10931 15691
rect 10873 15651 10931 15657
rect 10686 15580 10692 15632
rect 10744 15580 10750 15632
rect 9401 15487 9459 15493
rect 9401 15453 9413 15487
rect 9447 15453 9459 15487
rect 9401 15447 9459 15453
rect 9677 15487 9735 15493
rect 9677 15453 9689 15487
rect 9723 15484 9735 15487
rect 9950 15484 9956 15496
rect 9723 15456 9956 15484
rect 9723 15453 9735 15456
rect 9677 15447 9735 15453
rect 9416 15416 9444 15447
rect 9950 15444 9956 15456
rect 10008 15444 10014 15496
rect 10888 15484 10916 15651
rect 11422 15648 11428 15700
rect 11480 15648 11486 15700
rect 12894 15648 12900 15700
rect 12952 15648 12958 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 15010 15688 15016 15700
rect 13872 15660 15016 15688
rect 13872 15648 13878 15660
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 15286 15648 15292 15700
rect 15344 15648 15350 15700
rect 17954 15648 17960 15700
rect 18012 15648 18018 15700
rect 19794 15648 19800 15700
rect 19852 15688 19858 15700
rect 20990 15688 20996 15700
rect 19852 15660 20996 15688
rect 19852 15648 19858 15660
rect 20990 15648 20996 15660
rect 21048 15648 21054 15700
rect 21545 15691 21603 15697
rect 21545 15657 21557 15691
rect 21591 15688 21603 15691
rect 22094 15688 22100 15700
rect 21591 15660 22100 15688
rect 21591 15657 21603 15660
rect 21545 15651 21603 15657
rect 22094 15648 22100 15660
rect 22152 15688 22158 15700
rect 23290 15688 23296 15700
rect 22152 15660 23296 15688
rect 22152 15648 22158 15660
rect 23290 15648 23296 15660
rect 23348 15648 23354 15700
rect 25682 15648 25688 15700
rect 25740 15648 25746 15700
rect 26050 15648 26056 15700
rect 26108 15648 26114 15700
rect 26510 15648 26516 15700
rect 26568 15648 26574 15700
rect 27709 15691 27767 15697
rect 27709 15657 27721 15691
rect 27755 15688 27767 15691
rect 28166 15688 28172 15700
rect 27755 15660 28172 15688
rect 27755 15657 27767 15660
rect 27709 15651 27767 15657
rect 11330 15512 11336 15564
rect 11388 15512 11394 15564
rect 12158 15512 12164 15564
rect 12216 15512 12222 15564
rect 12805 15555 12863 15561
rect 12805 15521 12817 15555
rect 12851 15552 12863 15555
rect 12912 15552 12940 15648
rect 13354 15580 13360 15632
rect 13412 15580 13418 15632
rect 14734 15580 14740 15632
rect 14792 15620 14798 15632
rect 14792 15592 15238 15620
rect 14792 15580 14798 15592
rect 13725 15555 13783 15561
rect 13725 15552 13737 15555
rect 12851 15524 13737 15552
rect 12851 15521 12863 15524
rect 12805 15515 12863 15521
rect 13725 15521 13737 15524
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 11149 15487 11207 15493
rect 11149 15484 11161 15487
rect 10888 15456 11161 15484
rect 11149 15453 11161 15456
rect 11195 15453 11207 15487
rect 11348 15484 11376 15512
rect 11974 15484 11980 15496
rect 11348 15456 11980 15484
rect 11149 15447 11207 15453
rect 11974 15444 11980 15456
rect 12032 15444 12038 15496
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 14737 15487 14795 15493
rect 14737 15484 14749 15487
rect 14516 15456 14749 15484
rect 14516 15444 14522 15456
rect 14737 15453 14749 15456
rect 14783 15453 14795 15487
rect 14737 15447 14795 15453
rect 14826 15444 14832 15496
rect 14884 15484 14890 15496
rect 15102 15484 15108 15496
rect 14884 15456 15108 15484
rect 14884 15444 14890 15456
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 9766 15416 9772 15428
rect 9416 15388 9772 15416
rect 9766 15376 9772 15388
rect 9824 15416 9830 15428
rect 10410 15416 10416 15428
rect 9824 15388 10416 15416
rect 9824 15376 9830 15388
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 11054 15376 11060 15428
rect 11112 15416 11118 15428
rect 11241 15419 11299 15425
rect 11241 15416 11253 15419
rect 11112 15388 11253 15416
rect 11112 15376 11118 15388
rect 11241 15385 11253 15388
rect 11287 15385 11299 15419
rect 11241 15379 11299 15385
rect 11330 15376 11336 15428
rect 11388 15416 11394 15428
rect 11425 15419 11483 15425
rect 11425 15416 11437 15419
rect 11388 15388 11437 15416
rect 11388 15376 11394 15388
rect 11425 15385 11437 15388
rect 11471 15385 11483 15419
rect 11425 15379 11483 15385
rect 14918 15376 14924 15428
rect 14976 15376 14982 15428
rect 15013 15419 15071 15425
rect 15013 15385 15025 15419
rect 15059 15416 15071 15419
rect 15210 15416 15238 15592
rect 16393 15555 16451 15561
rect 16393 15521 16405 15555
rect 16439 15552 16451 15555
rect 17773 15555 17831 15561
rect 16439 15524 16988 15552
rect 16439 15521 16451 15524
rect 16393 15515 16451 15521
rect 15930 15484 15936 15496
rect 15488 15456 15936 15484
rect 15488 15428 15516 15456
rect 15930 15444 15936 15456
rect 15988 15444 15994 15496
rect 16022 15444 16028 15496
rect 16080 15444 16086 15496
rect 16209 15487 16267 15493
rect 16209 15453 16221 15487
rect 16255 15484 16267 15487
rect 16666 15484 16672 15496
rect 16255 15456 16672 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 16666 15444 16672 15456
rect 16724 15444 16730 15496
rect 16758 15444 16764 15496
rect 16816 15444 16822 15496
rect 16960 15493 16988 15524
rect 17773 15521 17785 15555
rect 17819 15552 17831 15555
rect 17972 15552 18000 15648
rect 17819 15524 18000 15552
rect 17819 15521 17831 15524
rect 17773 15515 17831 15521
rect 24854 15512 24860 15564
rect 24912 15552 24918 15564
rect 25700 15561 25728 15648
rect 25685 15555 25743 15561
rect 24912 15524 25176 15552
rect 24912 15512 24918 15524
rect 16945 15487 17003 15493
rect 16945 15453 16957 15487
rect 16991 15484 17003 15487
rect 17586 15484 17592 15496
rect 16991 15456 17592 15484
rect 16991 15453 17003 15456
rect 16945 15447 17003 15453
rect 17586 15444 17592 15456
rect 17644 15444 17650 15496
rect 20898 15444 20904 15496
rect 20956 15484 20962 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20956 15456 21097 15484
rect 20956 15444 20962 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 21174 15444 21180 15496
rect 21232 15444 21238 15496
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15484 21419 15487
rect 21818 15484 21824 15496
rect 21407 15456 21824 15484
rect 21407 15453 21419 15456
rect 21361 15447 21419 15453
rect 21818 15444 21824 15456
rect 21876 15444 21882 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 25148 15493 25176 15524
rect 25685 15521 25697 15555
rect 25731 15521 25743 15555
rect 25685 15515 25743 15521
rect 24949 15487 25007 15493
rect 24949 15484 24961 15487
rect 24728 15456 24961 15484
rect 24728 15444 24734 15456
rect 24949 15453 24961 15456
rect 24995 15453 25007 15487
rect 24949 15447 25007 15453
rect 25133 15487 25191 15493
rect 25133 15453 25145 15487
rect 25179 15453 25191 15487
rect 26068 15470 26096 15648
rect 26528 15620 26556 15648
rect 27157 15623 27215 15629
rect 27157 15620 27169 15623
rect 26528 15592 27169 15620
rect 27157 15589 27169 15592
rect 27203 15589 27215 15623
rect 27157 15583 27215 15589
rect 27249 15623 27307 15629
rect 27249 15589 27261 15623
rect 27295 15620 27307 15623
rect 27724 15620 27752 15651
rect 28166 15648 28172 15660
rect 28224 15648 28230 15700
rect 27295 15592 27752 15620
rect 27295 15589 27307 15592
rect 27249 15583 27307 15589
rect 26513 15555 26571 15561
rect 26513 15521 26525 15555
rect 26559 15552 26571 15555
rect 26970 15552 26976 15564
rect 26559 15524 26976 15552
rect 26559 15521 26571 15524
rect 26513 15515 26571 15521
rect 26970 15512 26976 15524
rect 27028 15512 27034 15564
rect 27172 15552 27200 15583
rect 27617 15555 27675 15561
rect 27617 15552 27629 15555
rect 27172 15524 27629 15552
rect 27617 15521 27629 15524
rect 27663 15521 27675 15555
rect 27617 15515 27675 15521
rect 27065 15487 27123 15493
rect 27065 15484 27077 15487
rect 25133 15447 25191 15453
rect 26620 15456 27077 15484
rect 15470 15416 15476 15428
rect 15059 15388 15476 15416
rect 15059 15385 15071 15388
rect 15013 15379 15071 15385
rect 15470 15376 15476 15388
rect 15528 15376 15534 15428
rect 16040 15416 16068 15444
rect 15948 15388 16068 15416
rect 9493 15351 9551 15357
rect 9493 15317 9505 15351
rect 9539 15348 9551 15351
rect 10686 15348 10692 15360
rect 9539 15320 10692 15348
rect 9539 15317 9551 15320
rect 9493 15311 9551 15317
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 10873 15351 10931 15357
rect 10873 15317 10885 15351
rect 10919 15348 10931 15351
rect 11348 15348 11376 15376
rect 10919 15320 11376 15348
rect 10919 15317 10931 15320
rect 10873 15311 10931 15317
rect 12894 15308 12900 15360
rect 12952 15348 12958 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 12952 15320 13093 15348
rect 12952 15308 12958 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13081 15311 13139 15317
rect 13262 15308 13268 15360
rect 13320 15308 13326 15360
rect 14936 15348 14964 15376
rect 15948 15348 15976 15388
rect 14936 15320 15976 15348
rect 25041 15351 25099 15357
rect 25041 15317 25053 15351
rect 25087 15348 25099 15351
rect 26620 15348 26648 15456
rect 27065 15453 27077 15456
rect 27111 15453 27123 15487
rect 27065 15447 27123 15453
rect 27341 15487 27399 15493
rect 27341 15453 27353 15487
rect 27387 15484 27399 15487
rect 27430 15484 27436 15496
rect 27387 15456 27436 15484
rect 27387 15453 27399 15456
rect 27341 15447 27399 15453
rect 27080 15416 27108 15447
rect 27430 15444 27436 15456
rect 27488 15484 27494 15496
rect 27893 15487 27951 15493
rect 27893 15484 27905 15487
rect 27488 15456 27905 15484
rect 27488 15444 27494 15456
rect 27893 15453 27905 15456
rect 27939 15453 27951 15487
rect 27893 15447 27951 15453
rect 27525 15419 27583 15425
rect 27525 15416 27537 15419
rect 27080 15388 27537 15416
rect 27525 15385 27537 15388
rect 27571 15385 27583 15419
rect 28166 15416 28172 15428
rect 27525 15379 27583 15385
rect 27724 15388 28172 15416
rect 25087 15320 26648 15348
rect 26881 15351 26939 15357
rect 25087 15317 25099 15320
rect 25041 15311 25099 15317
rect 26881 15317 26893 15351
rect 26927 15348 26939 15351
rect 27724 15348 27752 15388
rect 28166 15376 28172 15388
rect 28224 15376 28230 15428
rect 26927 15320 27752 15348
rect 26927 15317 26939 15320
rect 26881 15311 26939 15317
rect 27798 15308 27804 15360
rect 27856 15308 27862 15360
rect 1104 15258 35236 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 35236 15258
rect 1104 15184 35236 15206
rect 9309 15147 9367 15153
rect 9309 15113 9321 15147
rect 9355 15144 9367 15147
rect 9490 15144 9496 15156
rect 9355 15116 9496 15144
rect 9355 15113 9367 15116
rect 9309 15107 9367 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 9677 15147 9735 15153
rect 9677 15113 9689 15147
rect 9723 15144 9735 15147
rect 9950 15144 9956 15156
rect 9723 15116 9956 15144
rect 9723 15113 9735 15116
rect 9677 15107 9735 15113
rect 9950 15104 9956 15116
rect 10008 15104 10014 15156
rect 10226 15104 10232 15156
rect 10284 15104 10290 15156
rect 10410 15144 10416 15156
rect 10336 15116 10416 15144
rect 9401 15079 9459 15085
rect 9401 15076 9413 15079
rect 9232 15048 9413 15076
rect 9232 15020 9260 15048
rect 9401 15045 9413 15048
rect 9447 15045 9459 15079
rect 9401 15039 9459 15045
rect 9766 15036 9772 15088
rect 9824 15036 9830 15088
rect 10336 15085 10364 15116
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10597 15147 10655 15153
rect 10597 15113 10609 15147
rect 10643 15144 10655 15147
rect 11054 15144 11060 15156
rect 10643 15116 11060 15144
rect 10643 15113 10655 15116
rect 10597 15107 10655 15113
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11974 15104 11980 15156
rect 12032 15104 12038 15156
rect 17126 15104 17132 15156
rect 17184 15104 17190 15156
rect 17221 15147 17279 15153
rect 17221 15113 17233 15147
rect 17267 15144 17279 15147
rect 17402 15144 17408 15156
rect 17267 15116 17408 15144
rect 17267 15113 17279 15116
rect 17221 15107 17279 15113
rect 17402 15104 17408 15116
rect 17460 15104 17466 15156
rect 21174 15104 21180 15156
rect 21232 15104 21238 15156
rect 9861 15079 9919 15085
rect 9861 15045 9873 15079
rect 9907 15076 9919 15079
rect 10321 15079 10379 15085
rect 9907 15048 10180 15076
rect 9907 15045 9919 15048
rect 9861 15039 9919 15045
rect 9772 15033 9830 15036
rect 9214 14968 9220 15020
rect 9272 14968 9278 15020
rect 9493 15011 9551 15017
rect 9493 14977 9505 15011
rect 9539 15008 9551 15011
rect 9582 15008 9588 15020
rect 9539 14980 9588 15008
rect 9539 14977 9551 14980
rect 9493 14971 9551 14977
rect 9582 14968 9588 14980
rect 9640 14968 9646 15020
rect 9674 14968 9680 15020
rect 9732 14968 9738 15020
rect 9772 14999 9784 15033
rect 9818 14999 9830 15033
rect 10152 15020 10180 15048
rect 10321 15045 10333 15079
rect 10367 15045 10379 15079
rect 10505 15079 10563 15085
rect 10505 15076 10517 15079
rect 10321 15039 10379 15045
rect 10428 15048 10517 15076
rect 9772 14993 9830 14999
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14940 9183 14943
rect 9692 14940 9720 14968
rect 9171 14912 9720 14940
rect 10060 14940 10088 14971
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10192 14998 10364 15008
rect 10428 14998 10456 15048
rect 10505 15045 10517 15048
rect 10551 15045 10563 15079
rect 11992 15076 12020 15104
rect 12621 15079 12679 15085
rect 11992 15048 12296 15076
rect 10505 15039 10563 15045
rect 10192 14980 10456 14998
rect 10192 14968 10198 14980
rect 10336 14970 10456 14980
rect 10597 15011 10655 15017
rect 10597 14977 10609 15011
rect 10643 15008 10655 15011
rect 10686 15008 10692 15020
rect 10643 14980 10692 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 10612 14940 10640 14971
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 11698 14968 11704 15020
rect 11756 15008 11762 15020
rect 11977 15011 12035 15017
rect 11977 15008 11989 15011
rect 11756 14980 11989 15008
rect 11756 14968 11762 14980
rect 11977 14977 11989 14980
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 12066 14968 12072 15020
rect 12124 15008 12130 15020
rect 12268 15017 12296 15048
rect 12360 15048 12572 15076
rect 12360 15017 12388 15048
rect 12161 15011 12219 15017
rect 12161 15008 12173 15011
rect 12124 14980 12173 15008
rect 12124 14968 12130 14980
rect 12161 14977 12173 14980
rect 12207 14977 12219 15011
rect 12161 14971 12219 14977
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 12345 15011 12403 15017
rect 12345 14977 12357 15011
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 10060 14912 10640 14940
rect 12544 14940 12572 15048
rect 12621 15045 12633 15079
rect 12667 15045 12679 15079
rect 12621 15039 12679 15045
rect 12636 15008 12664 15039
rect 15194 15036 15200 15088
rect 15252 15076 15258 15088
rect 15838 15076 15844 15088
rect 15252 15048 15844 15076
rect 15252 15036 15258 15048
rect 15838 15036 15844 15048
rect 15896 15076 15902 15088
rect 15896 15048 20760 15076
rect 15896 15036 15902 15048
rect 20732 15020 20760 15048
rect 20898 15036 20904 15088
rect 20956 15036 20962 15088
rect 21192 15076 21220 15104
rect 21361 15079 21419 15085
rect 21361 15076 21373 15079
rect 21192 15048 21373 15076
rect 21361 15045 21373 15048
rect 21407 15045 21419 15079
rect 21361 15039 21419 15045
rect 13081 15011 13139 15017
rect 13081 15008 13093 15011
rect 12636 14980 13093 15008
rect 13081 14977 13093 14980
rect 13127 14977 13139 15011
rect 13081 14971 13139 14977
rect 13262 14968 13268 15020
rect 13320 14968 13326 15020
rect 16942 14968 16948 15020
rect 17000 14968 17006 15020
rect 17494 15008 17500 15020
rect 17236 14980 17500 15008
rect 12618 14940 12624 14952
rect 12544 14912 12624 14940
rect 9171 14909 9183 14912
rect 9125 14903 9183 14909
rect 9692 14872 9720 14912
rect 12618 14900 12624 14912
rect 12676 14900 12682 14952
rect 16761 14943 16819 14949
rect 16761 14909 16773 14943
rect 16807 14940 16819 14943
rect 17236 14940 17264 14980
rect 17494 14968 17500 14980
rect 17552 14968 17558 15020
rect 17586 14968 17592 15020
rect 17644 14968 17650 15020
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 17957 15011 18015 15017
rect 17957 15008 17969 15011
rect 17920 14980 17969 15008
rect 17920 14968 17926 14980
rect 17957 14977 17969 14980
rect 18003 14977 18015 15011
rect 17957 14971 18015 14977
rect 18046 14968 18052 15020
rect 18104 14968 18110 15020
rect 19613 15011 19671 15017
rect 19613 14977 19625 15011
rect 19659 15008 19671 15011
rect 20070 15008 20076 15020
rect 19659 14980 20076 15008
rect 19659 14977 19671 14980
rect 19613 14971 19671 14977
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 20714 14968 20720 15020
rect 20772 14968 20778 15020
rect 20916 15008 20944 15036
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20916 14980 21189 15008
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 21453 15011 21511 15017
rect 21453 14977 21465 15011
rect 21499 15008 21511 15011
rect 21818 15008 21824 15020
rect 21499 14980 21824 15008
rect 21499 14977 21511 14980
rect 21453 14971 21511 14977
rect 21818 14968 21824 14980
rect 21876 14968 21882 15020
rect 16807 14912 17264 14940
rect 17681 14943 17739 14949
rect 16807 14909 16819 14912
rect 16761 14903 16819 14909
rect 17681 14909 17693 14943
rect 17727 14940 17739 14943
rect 18064 14940 18092 14968
rect 17727 14912 18092 14940
rect 17727 14909 17739 14912
rect 17681 14903 17739 14909
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19521 14943 19579 14949
rect 19521 14940 19533 14943
rect 19484 14912 19533 14940
rect 19484 14900 19490 14912
rect 19521 14909 19533 14912
rect 19567 14909 19579 14943
rect 24854 14940 24860 14952
rect 19521 14903 19579 14909
rect 19628 14912 24860 14940
rect 9950 14872 9956 14884
rect 9692 14844 9956 14872
rect 9950 14832 9956 14844
rect 10008 14832 10014 14884
rect 13081 14875 13139 14881
rect 13081 14841 13093 14875
rect 13127 14872 13139 14875
rect 19628 14872 19656 14912
rect 24854 14900 24860 14912
rect 24912 14900 24918 14952
rect 13127 14844 19656 14872
rect 13127 14841 13139 14844
rect 13081 14835 13139 14841
rect 19978 14832 19984 14884
rect 20036 14832 20042 14884
rect 20806 14832 20812 14884
rect 20864 14872 20870 14884
rect 23934 14872 23940 14884
rect 20864 14844 23940 14872
rect 20864 14832 20870 14844
rect 23934 14832 23940 14844
rect 23992 14832 23998 14884
rect 15286 14764 15292 14816
rect 15344 14804 15350 14816
rect 16022 14804 16028 14816
rect 15344 14776 16028 14804
rect 15344 14764 15350 14776
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 17773 14807 17831 14813
rect 17773 14773 17785 14807
rect 17819 14804 17831 14807
rect 17954 14804 17960 14816
rect 17819 14776 17960 14804
rect 17819 14773 17831 14776
rect 17773 14767 17831 14773
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 21450 14764 21456 14816
rect 21508 14764 21514 14816
rect 1104 14714 35248 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 35248 14714
rect 1104 14640 35248 14662
rect 9677 14603 9735 14609
rect 9677 14569 9689 14603
rect 9723 14600 9735 14603
rect 9766 14600 9772 14612
rect 9723 14572 9772 14600
rect 9723 14569 9735 14572
rect 9677 14563 9735 14569
rect 9766 14560 9772 14572
rect 9824 14560 9830 14612
rect 10045 14603 10103 14609
rect 10045 14569 10057 14603
rect 10091 14600 10103 14603
rect 10134 14600 10140 14612
rect 10091 14572 10140 14600
rect 10091 14569 10103 14572
rect 10045 14563 10103 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 12158 14560 12164 14612
rect 12216 14560 12222 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14976 14572 15117 14600
rect 14976 14560 14982 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 15565 14603 15623 14609
rect 15565 14569 15577 14603
rect 15611 14600 15623 14603
rect 15654 14600 15660 14612
rect 15611 14572 15660 14600
rect 15611 14569 15623 14572
rect 15565 14563 15623 14569
rect 15654 14560 15660 14572
rect 15712 14600 15718 14612
rect 16301 14603 16359 14609
rect 15712 14572 16252 14600
rect 15712 14560 15718 14572
rect 9214 14492 9220 14544
rect 9272 14532 9278 14544
rect 10318 14532 10324 14544
rect 9272 14504 10324 14532
rect 9272 14492 9278 14504
rect 9582 14464 9588 14476
rect 9140 14436 9588 14464
rect 9140 14408 9168 14436
rect 9582 14424 9588 14436
rect 9640 14464 9646 14476
rect 9640 14436 9812 14464
rect 9640 14424 9646 14436
rect 9122 14356 9128 14408
rect 9180 14356 9186 14408
rect 9490 14356 9496 14408
rect 9548 14356 9554 14408
rect 9784 14405 9812 14436
rect 9876 14405 9904 14504
rect 10318 14492 10324 14504
rect 10376 14492 10382 14544
rect 11606 14492 11612 14544
rect 11664 14532 11670 14544
rect 12066 14532 12072 14544
rect 11664 14504 12072 14532
rect 11664 14492 11670 14504
rect 12066 14492 12072 14504
rect 12124 14532 12130 14544
rect 12345 14535 12403 14541
rect 12124 14504 12296 14532
rect 12124 14492 12130 14504
rect 9950 14424 9956 14476
rect 10008 14464 10014 14476
rect 10137 14467 10195 14473
rect 10137 14464 10149 14467
rect 10008 14436 10149 14464
rect 10008 14424 10014 14436
rect 10137 14433 10149 14436
rect 10183 14433 10195 14467
rect 10137 14427 10195 14433
rect 10502 14424 10508 14476
rect 10560 14464 10566 14476
rect 12268 14464 12296 14504
rect 12345 14501 12357 14535
rect 12391 14532 12403 14535
rect 12526 14532 12532 14544
rect 12391 14504 12532 14532
rect 12391 14501 12403 14504
rect 12345 14495 12403 14501
rect 12526 14492 12532 14504
rect 12584 14492 12590 14544
rect 16114 14532 16120 14544
rect 13648 14504 16120 14532
rect 10560 14436 11928 14464
rect 12268 14436 12572 14464
rect 10560 14424 10566 14436
rect 9769 14399 9827 14405
rect 9769 14365 9781 14399
rect 9815 14365 9827 14399
rect 9769 14359 9827 14365
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14365 9919 14399
rect 9861 14359 9919 14365
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 11606 14396 11612 14408
rect 11563 14368 11612 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 11606 14356 11612 14368
rect 11664 14356 11670 14408
rect 11698 14356 11704 14408
rect 11756 14356 11762 14408
rect 11900 14405 11928 14436
rect 11793 14399 11851 14405
rect 11793 14365 11805 14399
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 12345 14399 12403 14405
rect 12345 14365 12357 14399
rect 12391 14396 12403 14399
rect 12434 14396 12440 14408
rect 12391 14368 12440 14396
rect 12391 14365 12403 14368
rect 12345 14359 12403 14365
rect 9214 14288 9220 14340
rect 9272 14328 9278 14340
rect 9309 14331 9367 14337
rect 9309 14328 9321 14331
rect 9272 14300 9321 14328
rect 9272 14288 9278 14300
rect 9309 14297 9321 14300
rect 9355 14297 9367 14331
rect 9309 14291 9367 14297
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14297 9459 14331
rect 9508 14328 9536 14356
rect 11716 14328 11744 14356
rect 9508 14300 9996 14328
rect 9401 14291 9459 14297
rect 9416 14260 9444 14291
rect 9674 14260 9680 14272
rect 9416 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 9968 14269 9996 14300
rect 11348 14300 11744 14328
rect 9953 14263 10011 14269
rect 9953 14229 9965 14263
rect 9999 14229 10011 14263
rect 9953 14223 10011 14229
rect 11054 14220 11060 14272
rect 11112 14220 11118 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 11348 14269 11376 14300
rect 11808 14272 11836 14359
rect 11900 14328 11928 14359
rect 12434 14356 12440 14368
rect 12492 14356 12498 14408
rect 12544 14405 12572 14436
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12676 14436 13001 14464
rect 12676 14424 12682 14436
rect 12989 14433 13001 14436
rect 13035 14464 13047 14467
rect 13173 14467 13231 14473
rect 13173 14464 13185 14467
rect 13035 14436 13185 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 13173 14433 13185 14436
rect 13219 14433 13231 14467
rect 13173 14427 13231 14433
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12894 14356 12900 14408
rect 12952 14356 12958 14408
rect 13262 14356 13268 14408
rect 13320 14356 13326 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 13648 14396 13676 14504
rect 16114 14492 16120 14504
rect 16172 14492 16178 14544
rect 16224 14532 16252 14572
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 16758 14600 16764 14612
rect 16347 14572 16764 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 16758 14560 16764 14572
rect 16816 14560 16822 14612
rect 17494 14560 17500 14612
rect 17552 14560 17558 14612
rect 17862 14560 17868 14612
rect 17920 14560 17926 14612
rect 18046 14560 18052 14612
rect 18104 14600 18110 14612
rect 18233 14603 18291 14609
rect 18233 14600 18245 14603
rect 18104 14572 18245 14600
rect 18104 14560 18110 14572
rect 18233 14569 18245 14572
rect 18279 14569 18291 14603
rect 22094 14600 22100 14612
rect 18233 14563 18291 14569
rect 21284 14572 22100 14600
rect 17880 14532 17908 14560
rect 16224 14504 17908 14532
rect 17773 14467 17831 14473
rect 17773 14464 17785 14467
rect 14108 14436 15700 14464
rect 13587 14368 13676 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 13556 14328 13584 14359
rect 13998 14356 14004 14408
rect 14056 14396 14062 14408
rect 14108 14405 14136 14436
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 14056 14368 14105 14396
rect 14056 14356 14062 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14369 14399 14427 14405
rect 14369 14365 14381 14399
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14461 14399 14519 14405
rect 14461 14365 14473 14399
rect 14507 14396 14519 14399
rect 15286 14396 15292 14408
rect 14507 14368 15292 14396
rect 14507 14365 14519 14368
rect 14461 14359 14519 14365
rect 14292 14328 14320 14359
rect 11900 14300 13584 14328
rect 13924 14300 14320 14328
rect 14384 14328 14412 14359
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15672 14405 15700 14436
rect 15948 14436 17785 14464
rect 15948 14408 15976 14436
rect 17773 14433 17785 14436
rect 17819 14464 17831 14467
rect 17819 14436 18276 14464
rect 17819 14433 17831 14436
rect 17773 14427 17831 14433
rect 15381 14399 15439 14405
rect 15381 14365 15393 14399
rect 15427 14365 15439 14399
rect 15381 14359 15439 14365
rect 15657 14399 15715 14405
rect 15657 14365 15669 14399
rect 15703 14365 15715 14399
rect 15657 14359 15715 14365
rect 15396 14328 15424 14359
rect 15838 14356 15844 14408
rect 15896 14356 15902 14408
rect 15930 14356 15936 14408
rect 15988 14356 15994 14408
rect 16022 14356 16028 14408
rect 16080 14396 16086 14408
rect 17681 14399 17739 14405
rect 17681 14396 17693 14399
rect 16080 14368 17693 14396
rect 16080 14356 16086 14368
rect 17681 14365 17693 14368
rect 17727 14396 17739 14399
rect 18049 14399 18107 14405
rect 18049 14396 18061 14399
rect 17727 14368 18061 14396
rect 17727 14365 17739 14368
rect 17681 14359 17739 14365
rect 18049 14365 18061 14368
rect 18095 14396 18107 14399
rect 18138 14396 18144 14408
rect 18095 14368 18144 14396
rect 18095 14365 18107 14368
rect 18049 14359 18107 14365
rect 18138 14356 18144 14368
rect 18196 14356 18202 14408
rect 18248 14405 18276 14436
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14365 18291 14399
rect 18233 14359 18291 14365
rect 20806 14356 20812 14408
rect 20864 14356 20870 14408
rect 14384 14300 15424 14328
rect 15565 14331 15623 14337
rect 13924 14272 13952 14300
rect 14568 14272 14596 14300
rect 15565 14297 15577 14331
rect 15611 14328 15623 14331
rect 15746 14328 15752 14340
rect 15611 14300 15752 14328
rect 15611 14297 15623 14300
rect 15565 14291 15623 14297
rect 15746 14288 15752 14300
rect 15804 14328 15810 14340
rect 15804 14300 16436 14328
rect 15804 14288 15810 14300
rect 11333 14263 11391 14269
rect 11333 14260 11345 14263
rect 11204 14232 11345 14260
rect 11204 14220 11210 14232
rect 11333 14229 11345 14232
rect 11379 14229 11391 14263
rect 11333 14223 11391 14229
rect 11790 14220 11796 14272
rect 11848 14220 11854 14272
rect 13630 14220 13636 14272
rect 13688 14260 13694 14272
rect 13817 14263 13875 14269
rect 13817 14260 13829 14263
rect 13688 14232 13829 14260
rect 13688 14220 13694 14232
rect 13817 14229 13829 14232
rect 13863 14229 13875 14263
rect 13817 14223 13875 14229
rect 13906 14220 13912 14272
rect 13964 14220 13970 14272
rect 14550 14220 14556 14272
rect 14608 14220 14614 14272
rect 14734 14220 14740 14272
rect 14792 14220 14798 14272
rect 16408 14260 16436 14300
rect 17954 14288 17960 14340
rect 18012 14328 18018 14340
rect 20824 14328 20852 14356
rect 18012 14300 20852 14328
rect 21284 14328 21312 14572
rect 22094 14560 22100 14572
rect 22152 14560 22158 14612
rect 23658 14560 23664 14612
rect 23716 14560 23722 14612
rect 23934 14560 23940 14612
rect 23992 14600 23998 14612
rect 24397 14603 24455 14609
rect 24397 14600 24409 14603
rect 23992 14572 24409 14600
rect 23992 14560 23998 14572
rect 24397 14569 24409 14572
rect 24443 14569 24455 14603
rect 24397 14563 24455 14569
rect 21821 14535 21879 14541
rect 21821 14501 21833 14535
rect 21867 14532 21879 14535
rect 22186 14532 22192 14544
rect 21867 14504 22192 14532
rect 21867 14501 21879 14504
rect 21821 14495 21879 14501
rect 22186 14492 22192 14504
rect 22244 14492 22250 14544
rect 24029 14535 24087 14541
rect 24029 14501 24041 14535
rect 24075 14501 24087 14535
rect 24029 14495 24087 14501
rect 24765 14535 24823 14541
rect 24765 14501 24777 14535
rect 24811 14501 24823 14535
rect 24765 14495 24823 14501
rect 21450 14424 21456 14476
rect 21508 14424 21514 14476
rect 21542 14424 21548 14476
rect 21600 14464 21606 14476
rect 21600 14436 22156 14464
rect 21600 14424 21606 14436
rect 21361 14399 21419 14405
rect 21361 14365 21373 14399
rect 21407 14396 21419 14399
rect 21468 14396 21496 14424
rect 21407 14368 21496 14396
rect 21637 14399 21695 14405
rect 21407 14365 21419 14368
rect 21361 14359 21419 14365
rect 21637 14365 21649 14399
rect 21683 14396 21695 14399
rect 21683 14368 21956 14396
rect 21683 14365 21695 14368
rect 21637 14359 21695 14365
rect 21928 14340 21956 14368
rect 21453 14331 21511 14337
rect 21453 14328 21465 14331
rect 21284 14300 21465 14328
rect 18012 14288 18018 14300
rect 21453 14297 21465 14300
rect 21499 14297 21511 14331
rect 21453 14291 21511 14297
rect 21910 14288 21916 14340
rect 21968 14337 21974 14340
rect 22128 14337 22156 14436
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 23753 14467 23811 14473
rect 23753 14464 23765 14467
rect 23440 14436 23765 14464
rect 23440 14424 23446 14436
rect 23753 14433 23765 14436
rect 23799 14433 23811 14467
rect 24044 14464 24072 14495
rect 24780 14464 24808 14495
rect 25038 14464 25044 14476
rect 24044 14436 24716 14464
rect 24780 14436 25044 14464
rect 23753 14427 23811 14433
rect 23014 14356 23020 14408
rect 23072 14396 23078 14408
rect 23477 14399 23535 14405
rect 23477 14396 23489 14399
rect 23072 14368 23489 14396
rect 23072 14356 23078 14368
rect 23477 14365 23489 14368
rect 23523 14365 23535 14399
rect 23477 14359 23535 14365
rect 23566 14356 23572 14408
rect 23624 14396 23630 14408
rect 24394 14396 24400 14408
rect 23624 14368 24400 14396
rect 23624 14356 23630 14368
rect 24394 14356 24400 14368
rect 24452 14356 24458 14408
rect 24486 14356 24492 14408
rect 24544 14356 24550 14408
rect 24688 14396 24716 14436
rect 25038 14424 25044 14436
rect 25096 14464 25102 14476
rect 25777 14467 25835 14473
rect 25777 14464 25789 14467
rect 25096 14436 25789 14464
rect 25096 14424 25102 14436
rect 24854 14396 24860 14408
rect 24688 14368 24860 14396
rect 24854 14356 24860 14368
rect 24912 14396 24918 14408
rect 25148 14405 25176 14436
rect 25777 14433 25789 14436
rect 25823 14433 25835 14467
rect 25777 14427 25835 14433
rect 24949 14399 25007 14405
rect 24949 14396 24961 14399
rect 24912 14368 24961 14396
rect 24912 14356 24918 14368
rect 24949 14365 24961 14368
rect 24995 14365 25007 14399
rect 24949 14359 25007 14365
rect 25133 14399 25191 14405
rect 25133 14365 25145 14399
rect 25179 14365 25191 14399
rect 25593 14399 25651 14405
rect 25593 14396 25605 14399
rect 25133 14359 25191 14365
rect 25240 14368 25605 14396
rect 21968 14331 21997 14337
rect 21985 14297 21997 14331
rect 21968 14291 21997 14297
rect 22113 14331 22171 14337
rect 22113 14297 22125 14331
rect 22159 14297 22171 14331
rect 22370 14328 22376 14340
rect 22113 14291 22171 14297
rect 22204 14300 22376 14328
rect 21968 14288 21974 14291
rect 21174 14260 21180 14272
rect 16408 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 21266 14220 21272 14272
rect 21324 14260 21330 14272
rect 22204 14260 22232 14300
rect 22370 14288 22376 14300
rect 22428 14328 22434 14340
rect 24964 14328 24992 14359
rect 25240 14328 25268 14368
rect 25593 14365 25605 14368
rect 25639 14365 25651 14399
rect 25593 14359 25651 14365
rect 25869 14399 25927 14405
rect 25869 14365 25881 14399
rect 25915 14365 25927 14399
rect 25869 14359 25927 14365
rect 22428 14300 24164 14328
rect 24964 14300 25268 14328
rect 22428 14288 22434 14300
rect 24136 14272 24164 14300
rect 25314 14288 25320 14340
rect 25372 14328 25378 14340
rect 25884 14328 25912 14359
rect 26050 14356 26056 14408
rect 26108 14356 26114 14408
rect 25372 14300 25912 14328
rect 25372 14288 25378 14300
rect 21324 14232 22232 14260
rect 21324 14220 21330 14232
rect 22278 14220 22284 14272
rect 22336 14220 22342 14272
rect 23014 14220 23020 14272
rect 23072 14260 23078 14272
rect 23293 14263 23351 14269
rect 23293 14260 23305 14263
rect 23072 14232 23305 14260
rect 23072 14220 23078 14232
rect 23293 14229 23305 14232
rect 23339 14229 23351 14263
rect 23293 14223 23351 14229
rect 24118 14220 24124 14272
rect 24176 14220 24182 14272
rect 25406 14220 25412 14272
rect 25464 14220 25470 14272
rect 25866 14220 25872 14272
rect 25924 14220 25930 14272
rect 1104 14170 35236 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 35236 14170
rect 1104 14096 35236 14118
rect 9401 14059 9459 14065
rect 9401 14025 9413 14059
rect 9447 14056 9459 14059
rect 9490 14056 9496 14068
rect 9447 14028 9496 14056
rect 9447 14025 9459 14028
rect 9401 14019 9459 14025
rect 9490 14016 9496 14028
rect 9548 14016 9554 14068
rect 9674 14016 9680 14068
rect 9732 14056 9738 14068
rect 10229 14059 10287 14065
rect 10229 14056 10241 14059
rect 9732 14028 10241 14056
rect 9732 14016 9738 14028
rect 10229 14025 10241 14028
rect 10275 14025 10287 14059
rect 10229 14019 10287 14025
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11790 14056 11796 14068
rect 11112 14028 11796 14056
rect 11112 14016 11118 14028
rect 11790 14016 11796 14028
rect 11848 14056 11854 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 11848 14028 12173 14056
rect 11848 14016 11854 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 12434 14016 12440 14068
rect 12492 14056 12498 14068
rect 12713 14059 12771 14065
rect 12713 14056 12725 14059
rect 12492 14028 12725 14056
rect 12492 14016 12498 14028
rect 12713 14025 12725 14028
rect 12759 14025 12771 14059
rect 12713 14019 12771 14025
rect 13262 14016 13268 14068
rect 13320 14016 13326 14068
rect 14458 14016 14464 14068
rect 14516 14016 14522 14068
rect 15841 14059 15899 14065
rect 14660 14028 15332 14056
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13988 10011 13991
rect 12805 13991 12863 13997
rect 12805 13988 12817 13991
rect 9999 13960 12817 13988
rect 9999 13957 10011 13960
rect 9953 13951 10011 13957
rect 9677 13923 9735 13929
rect 9677 13889 9689 13923
rect 9723 13920 9735 13923
rect 9723 13892 9996 13920
rect 9723 13889 9735 13892
rect 9677 13883 9735 13889
rect 9968 13864 9996 13892
rect 10428 13892 10640 13920
rect 9585 13855 9643 13861
rect 9585 13821 9597 13855
rect 9631 13821 9643 13855
rect 9585 13815 9643 13821
rect 8846 13744 8852 13796
rect 8904 13784 8910 13796
rect 9600 13784 9628 13815
rect 9950 13812 9956 13864
rect 10008 13812 10014 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13852 10103 13855
rect 10318 13852 10324 13864
rect 10091 13824 10324 13852
rect 10091 13821 10103 13824
rect 10045 13815 10103 13821
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 10428 13784 10456 13892
rect 10502 13812 10508 13864
rect 10560 13812 10566 13864
rect 10612 13793 10640 13892
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 10873 13923 10931 13929
rect 10873 13920 10885 13923
rect 10836 13892 10885 13920
rect 10836 13880 10842 13892
rect 10873 13889 10885 13892
rect 10919 13889 10931 13923
rect 10873 13883 10931 13889
rect 12452 13864 12480 13960
rect 12805 13957 12817 13960
rect 12851 13957 12863 13991
rect 12805 13951 12863 13957
rect 12529 13923 12587 13929
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 13280 13920 13308 14016
rect 13817 13991 13875 13997
rect 13817 13957 13829 13991
rect 13863 13988 13875 13991
rect 13906 13988 13912 14000
rect 13863 13960 13912 13988
rect 13863 13957 13875 13960
rect 13817 13951 13875 13957
rect 13906 13948 13912 13960
rect 13964 13948 13970 14000
rect 14660 13988 14688 14028
rect 14108 13960 14688 13988
rect 12575 13892 13308 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 12345 13855 12403 13861
rect 12345 13852 12357 13855
rect 10796 13824 12357 13852
rect 8904 13756 10456 13784
rect 10597 13787 10655 13793
rect 8904 13744 8910 13756
rect 10597 13753 10609 13787
rect 10643 13784 10655 13787
rect 10796 13784 10824 13824
rect 12345 13821 12357 13824
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 12434 13812 12440 13864
rect 12492 13812 12498 13864
rect 10870 13784 10876 13796
rect 10643 13756 10876 13784
rect 10643 13753 10655 13756
rect 10597 13747 10655 13753
rect 10870 13744 10876 13756
rect 10928 13744 10934 13796
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 12544 13784 12572 13883
rect 12894 13812 12900 13864
rect 12952 13852 12958 13864
rect 13630 13852 13636 13864
rect 12952 13824 13636 13852
rect 12952 13812 12958 13824
rect 13630 13812 13636 13824
rect 13688 13812 13694 13864
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 14108 13852 14136 13960
rect 14734 13948 14740 14000
rect 14792 13988 14798 14000
rect 14792 13960 15056 13988
rect 14792 13948 14798 13960
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 14458 13920 14464 13932
rect 14231 13892 14464 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14642 13880 14648 13932
rect 14700 13920 14706 13932
rect 14829 13923 14887 13929
rect 14829 13920 14841 13923
rect 14700 13892 14841 13920
rect 14700 13880 14706 13892
rect 14829 13889 14841 13892
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 14918 13880 14924 13932
rect 14976 13880 14982 13932
rect 15028 13929 15056 13960
rect 15194 13948 15200 14000
rect 15252 13948 15258 14000
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15013 13883 15071 13889
rect 13955 13824 14136 13852
rect 14277 13855 14335 13861
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 14277 13821 14289 13855
rect 14323 13821 14335 13855
rect 14277 13815 14335 13821
rect 11848 13756 12572 13784
rect 14292 13784 14320 13815
rect 14366 13812 14372 13864
rect 14424 13852 14430 13864
rect 14553 13855 14611 13861
rect 14553 13852 14565 13855
rect 14424 13824 14565 13852
rect 14424 13812 14430 13824
rect 14553 13821 14565 13824
rect 14599 13821 14611 13855
rect 14553 13815 14611 13821
rect 14737 13855 14795 13861
rect 14737 13821 14749 13855
rect 14783 13852 14795 13855
rect 15212 13852 15240 13948
rect 15304 13864 15332 14028
rect 15841 14025 15853 14059
rect 15887 14056 15899 14059
rect 16942 14056 16948 14068
rect 15887 14028 16948 14056
rect 15887 14025 15899 14028
rect 15841 14019 15899 14025
rect 16942 14016 16948 14028
rect 17000 14016 17006 14068
rect 18693 14059 18751 14065
rect 18693 14025 18705 14059
rect 18739 14056 18751 14059
rect 19061 14059 19119 14065
rect 18739 14028 19012 14056
rect 18739 14025 18751 14028
rect 18693 14019 18751 14025
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 18417 13991 18475 13997
rect 18417 13988 18429 13991
rect 17736 13960 18429 13988
rect 17736 13948 17742 13960
rect 18417 13957 18429 13960
rect 18463 13988 18475 13991
rect 18463 13960 18828 13988
rect 18463 13957 18475 13960
rect 18417 13951 18475 13957
rect 18800 13929 18828 13960
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13920 15623 13923
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 15611 13892 15976 13920
rect 15611 13889 15623 13892
rect 15565 13883 15623 13889
rect 14783 13824 15240 13852
rect 14783 13821 14795 13824
rect 14737 13815 14795 13821
rect 15286 13812 15292 13864
rect 15344 13812 15350 13864
rect 15654 13852 15660 13864
rect 15396 13824 15660 13852
rect 15396 13784 15424 13824
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15948 13796 15976 13892
rect 17972 13892 18705 13920
rect 17972 13796 18000 13892
rect 18616 13852 18644 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13889 18843 13923
rect 18984 13920 19012 14028
rect 19061 14025 19073 14059
rect 19107 14056 19119 14059
rect 19705 14059 19763 14065
rect 19107 14028 19472 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 19444 13932 19472 14028
rect 19705 14025 19717 14059
rect 19751 14056 19763 14059
rect 20070 14056 20076 14068
rect 19751 14028 20076 14056
rect 19751 14025 19763 14028
rect 19705 14019 19763 14025
rect 20070 14016 20076 14028
rect 20128 14016 20134 14068
rect 20806 14016 20812 14068
rect 20864 14016 20870 14068
rect 21910 14016 21916 14068
rect 21968 14016 21974 14068
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 22741 14059 22799 14065
rect 22741 14056 22753 14059
rect 22520 14028 22753 14056
rect 22520 14016 22526 14028
rect 22741 14025 22753 14028
rect 22787 14025 22799 14059
rect 22741 14019 22799 14025
rect 23106 14016 23112 14068
rect 23164 14056 23170 14068
rect 23164 14028 23612 14056
rect 23164 14016 23170 14028
rect 22189 13991 22247 13997
rect 22189 13988 22201 13991
rect 21100 13960 22201 13988
rect 19334 13920 19340 13932
rect 18984 13892 19340 13920
rect 18785 13883 18843 13889
rect 19334 13880 19340 13892
rect 19392 13880 19398 13932
rect 19426 13880 19432 13932
rect 19484 13920 19490 13932
rect 19521 13923 19579 13929
rect 19521 13920 19533 13923
rect 19484 13892 19533 13920
rect 19484 13880 19490 13892
rect 19521 13889 19533 13892
rect 19567 13889 19579 13923
rect 19521 13883 19579 13889
rect 20714 13880 20720 13932
rect 20772 13880 20778 13932
rect 21100 13929 21128 13960
rect 22189 13957 22201 13960
rect 22235 13957 22247 13991
rect 22189 13951 22247 13957
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 21008 13892 21097 13920
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18616 13824 19073 13852
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19061 13815 19119 13821
rect 19245 13855 19303 13861
rect 19245 13821 19257 13855
rect 19291 13852 19303 13855
rect 19886 13852 19892 13864
rect 19291 13824 19892 13852
rect 19291 13821 19303 13824
rect 19245 13815 19303 13821
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 14292 13756 15424 13784
rect 11848 13744 11854 13756
rect 15930 13744 15936 13796
rect 15988 13744 15994 13796
rect 17954 13744 17960 13796
rect 18012 13744 18018 13796
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 18877 13787 18935 13793
rect 18877 13784 18889 13787
rect 18656 13756 18889 13784
rect 18656 13744 18662 13756
rect 18877 13753 18889 13756
rect 18923 13753 18935 13787
rect 18877 13747 18935 13753
rect 18966 13744 18972 13796
rect 19024 13784 19030 13796
rect 21008 13784 21036 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21266 13880 21272 13932
rect 21324 13920 21330 13932
rect 21361 13923 21419 13929
rect 21361 13920 21373 13923
rect 21324 13892 21373 13920
rect 21324 13880 21330 13892
rect 21361 13889 21373 13892
rect 21407 13889 21419 13923
rect 21361 13883 21419 13889
rect 21451 13923 21509 13929
rect 21451 13889 21463 13923
rect 21497 13889 21509 13923
rect 21451 13883 21509 13889
rect 21637 13923 21695 13929
rect 21637 13889 21649 13923
rect 21683 13920 21695 13923
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21683 13892 21833 13920
rect 21683 13889 21695 13892
rect 21637 13883 21695 13889
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 21462 13852 21490 13883
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 21968 13892 22017 13920
rect 21968 13880 21974 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22094 13852 22100 13864
rect 19024 13756 21036 13784
rect 21100 13824 22100 13852
rect 19024 13744 19030 13756
rect 10735 13719 10793 13725
rect 10735 13685 10747 13719
rect 10781 13716 10793 13719
rect 11054 13716 11060 13728
rect 10781 13688 11060 13716
rect 10781 13685 10793 13688
rect 10735 13679 10793 13685
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 21100 13716 21128 13824
rect 22094 13812 22100 13824
rect 22152 13812 22158 13864
rect 22204 13784 22232 13951
rect 22370 13948 22376 14000
rect 22428 13948 22434 14000
rect 22572 13960 23428 13988
rect 22572 13864 22600 13960
rect 23032 13929 23060 13960
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 23017 13923 23075 13929
rect 23017 13889 23029 13923
rect 23063 13889 23075 13923
rect 23017 13883 23075 13889
rect 22554 13812 22560 13864
rect 22612 13812 22618 13864
rect 22940 13852 22968 13883
rect 23106 13880 23112 13932
rect 23164 13880 23170 13932
rect 23400 13929 23428 13960
rect 23584 13929 23612 14028
rect 23658 14016 23664 14068
rect 23716 14016 23722 14068
rect 24394 14056 24400 14068
rect 23861 14028 24400 14056
rect 23676 13929 23704 14016
rect 23201 13923 23259 13929
rect 23201 13889 23213 13923
rect 23247 13889 23259 13923
rect 23201 13883 23259 13889
rect 23293 13923 23351 13929
rect 23293 13889 23305 13923
rect 23339 13889 23351 13923
rect 23293 13883 23351 13889
rect 23385 13923 23443 13929
rect 23385 13889 23397 13923
rect 23431 13889 23443 13923
rect 23385 13883 23443 13889
rect 23569 13923 23627 13929
rect 23569 13889 23581 13923
rect 23615 13889 23627 13923
rect 23569 13883 23627 13889
rect 23661 13923 23719 13929
rect 23661 13889 23673 13923
rect 23707 13889 23719 13923
rect 23661 13883 23719 13889
rect 23753 13923 23811 13929
rect 23753 13889 23765 13923
rect 23799 13920 23811 13923
rect 23861 13920 23889 14028
rect 24394 14016 24400 14028
rect 24452 14056 24458 14068
rect 24452 14028 24624 14056
rect 24452 14016 24458 14028
rect 24213 13991 24271 13997
rect 24213 13988 24225 13991
rect 23799 13892 23889 13920
rect 23952 13960 24225 13988
rect 23799 13889 23811 13892
rect 23753 13883 23811 13889
rect 23124 13852 23152 13880
rect 22940 13824 23152 13852
rect 23216 13784 23244 13883
rect 23308 13852 23336 13883
rect 23474 13852 23480 13864
rect 23308 13824 23480 13852
rect 23474 13812 23480 13824
rect 23532 13812 23538 13864
rect 23676 13852 23704 13883
rect 23952 13852 23980 13960
rect 24213 13957 24225 13960
rect 24259 13988 24271 13991
rect 24259 13960 24440 13988
rect 24259 13957 24271 13960
rect 24213 13951 24271 13957
rect 24026 13880 24032 13932
rect 24084 13880 24090 13932
rect 24118 13880 24124 13932
rect 24176 13880 24182 13932
rect 24412 13929 24440 13960
rect 24596 13929 24624 14028
rect 25314 14016 25320 14068
rect 25372 14016 25378 14068
rect 25406 14016 25412 14068
rect 25464 14016 25470 14068
rect 25866 14016 25872 14068
rect 25924 14016 25930 14068
rect 25332 13988 25360 14016
rect 25148 13960 25360 13988
rect 25148 13929 25176 13960
rect 24305 13923 24363 13929
rect 24305 13889 24317 13923
rect 24351 13889 24363 13923
rect 24305 13883 24363 13889
rect 24397 13923 24455 13929
rect 24397 13889 24409 13923
rect 24443 13889 24455 13923
rect 24397 13883 24455 13889
rect 24581 13923 24639 13929
rect 24581 13889 24593 13923
rect 24627 13889 24639 13923
rect 24581 13883 24639 13889
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 23676 13824 23980 13852
rect 24044 13852 24072 13880
rect 24320 13852 24348 13883
rect 24872 13852 24900 13883
rect 25222 13880 25228 13932
rect 25280 13880 25286 13932
rect 25424 13929 25452 14016
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25685 13923 25743 13929
rect 25685 13889 25697 13923
rect 25731 13920 25743 13923
rect 25884 13920 25912 14016
rect 25731 13892 25912 13920
rect 25731 13889 25743 13892
rect 25685 13883 25743 13889
rect 24044 13824 24348 13852
rect 24412 13824 25728 13852
rect 23676 13784 23704 13824
rect 24412 13784 24440 13824
rect 22204 13756 23152 13784
rect 23216 13756 23704 13784
rect 24044 13756 24440 13784
rect 25700 13784 25728 13824
rect 25774 13812 25780 13864
rect 25832 13812 25838 13864
rect 26970 13852 26976 13864
rect 25884 13824 26976 13852
rect 25884 13784 25912 13824
rect 26970 13812 26976 13824
rect 27028 13812 27034 13864
rect 25700 13756 25912 13784
rect 26053 13787 26111 13793
rect 14884 13688 21128 13716
rect 14884 13676 14890 13688
rect 21174 13676 21180 13728
rect 21232 13676 21238 13728
rect 23124 13716 23152 13756
rect 23290 13716 23296 13728
rect 23124 13688 23296 13716
rect 23290 13676 23296 13688
rect 23348 13676 23354 13728
rect 24044 13725 24072 13756
rect 26053 13753 26065 13787
rect 26099 13784 26111 13787
rect 26418 13784 26424 13796
rect 26099 13756 26424 13784
rect 26099 13753 26111 13756
rect 26053 13747 26111 13753
rect 26418 13744 26424 13756
rect 26476 13744 26482 13796
rect 24029 13719 24087 13725
rect 24029 13685 24041 13719
rect 24075 13685 24087 13719
rect 24029 13679 24087 13685
rect 24486 13676 24492 13728
rect 24544 13676 24550 13728
rect 24670 13676 24676 13728
rect 24728 13716 24734 13728
rect 24765 13719 24823 13725
rect 24765 13716 24777 13719
rect 24728 13688 24777 13716
rect 24728 13676 24734 13688
rect 24765 13685 24777 13688
rect 24811 13685 24823 13719
rect 24765 13679 24823 13685
rect 25406 13676 25412 13728
rect 25464 13676 25470 13728
rect 1104 13626 35248 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 35248 13626
rect 1104 13552 35248 13574
rect 10778 13512 10784 13524
rect 8956 13484 10784 13512
rect 8956 13184 8984 13484
rect 10778 13472 10784 13484
rect 10836 13512 10842 13524
rect 11974 13512 11980 13524
rect 10836 13484 11980 13512
rect 10836 13472 10842 13484
rect 11974 13472 11980 13484
rect 12032 13512 12038 13524
rect 14826 13512 14832 13524
rect 12032 13484 14832 13512
rect 12032 13472 12038 13484
rect 14826 13472 14832 13484
rect 14884 13472 14890 13524
rect 14921 13515 14979 13521
rect 14921 13481 14933 13515
rect 14967 13481 14979 13515
rect 14921 13475 14979 13481
rect 14185 13447 14243 13453
rect 14185 13413 14197 13447
rect 14231 13444 14243 13447
rect 14458 13444 14464 13456
rect 14231 13416 14464 13444
rect 14231 13413 14243 13416
rect 14185 13407 14243 13413
rect 14458 13404 14464 13416
rect 14516 13404 14522 13456
rect 14936 13444 14964 13475
rect 15010 13472 15016 13524
rect 15068 13472 15074 13524
rect 16960 13484 18644 13512
rect 16960 13444 16988 13484
rect 14936 13416 16988 13444
rect 17037 13447 17095 13453
rect 17037 13413 17049 13447
rect 17083 13413 17095 13447
rect 17037 13407 17095 13413
rect 17221 13447 17279 13453
rect 17221 13413 17233 13447
rect 17267 13444 17279 13447
rect 18616 13444 18644 13484
rect 23106 13472 23112 13524
rect 23164 13512 23170 13524
rect 23201 13515 23259 13521
rect 23201 13512 23213 13515
rect 23164 13484 23213 13512
rect 23164 13472 23170 13484
rect 23201 13481 23213 13484
rect 23247 13481 23259 13515
rect 23201 13475 23259 13481
rect 23474 13472 23480 13524
rect 23532 13472 23538 13524
rect 24486 13472 24492 13524
rect 24544 13512 24550 13524
rect 24581 13515 24639 13521
rect 24581 13512 24593 13515
rect 24544 13484 24593 13512
rect 24544 13472 24550 13484
rect 24581 13481 24593 13484
rect 24627 13481 24639 13515
rect 24581 13475 24639 13481
rect 21910 13444 21916 13456
rect 17267 13416 18552 13444
rect 18616 13416 21916 13444
rect 17267 13413 17279 13416
rect 17221 13407 17279 13413
rect 10502 13376 10508 13388
rect 9876 13348 10508 13376
rect 9876 13317 9904 13348
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 14826 13376 14832 13388
rect 14200 13348 14832 13376
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13277 9919 13311
rect 9861 13271 9919 13277
rect 9950 13268 9956 13320
rect 10008 13308 10014 13320
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 10008 13280 10057 13308
rect 10008 13268 10014 13280
rect 10045 13277 10057 13280
rect 10091 13308 10103 13311
rect 11054 13308 11060 13320
rect 10091 13280 11060 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 11054 13268 11060 13280
rect 11112 13268 11118 13320
rect 9677 13243 9735 13249
rect 9677 13209 9689 13243
rect 9723 13240 9735 13243
rect 9766 13240 9772 13252
rect 9723 13212 9772 13240
rect 9723 13209 9735 13212
rect 9677 13203 9735 13209
rect 9766 13200 9772 13212
rect 9824 13200 9830 13252
rect 10962 13240 10968 13252
rect 10336 13212 10968 13240
rect 8938 13132 8944 13184
rect 8996 13132 9002 13184
rect 10226 13132 10232 13184
rect 10284 13172 10290 13184
rect 10336 13181 10364 13212
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 13814 13200 13820 13252
rect 13872 13240 13878 13252
rect 14200 13249 14228 13348
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 14918 13336 14924 13388
rect 14976 13376 14982 13388
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 14976 13348 15577 13376
rect 14976 13336 14982 13348
rect 15565 13345 15577 13348
rect 15611 13345 15623 13379
rect 15565 13339 15623 13345
rect 16298 13336 16304 13388
rect 16356 13336 16362 13388
rect 14642 13268 14648 13320
rect 14700 13268 14706 13320
rect 14734 13268 14740 13320
rect 14792 13308 14798 13320
rect 15197 13311 15255 13317
rect 15197 13308 15209 13311
rect 14792 13280 15209 13308
rect 14792 13268 14798 13280
rect 15197 13277 15209 13280
rect 15243 13277 15255 13311
rect 15197 13271 15255 13277
rect 15289 13311 15347 13317
rect 15289 13277 15301 13311
rect 15335 13308 15347 13311
rect 15838 13308 15844 13320
rect 15335 13280 15844 13308
rect 15335 13277 15347 13280
rect 15289 13271 15347 13277
rect 15838 13268 15844 13280
rect 15896 13268 15902 13320
rect 16390 13268 16396 13320
rect 16448 13268 16454 13320
rect 16666 13268 16672 13320
rect 16724 13308 16730 13320
rect 17052 13308 17080 13407
rect 17328 13348 17816 13376
rect 17328 13320 17356 13348
rect 16724 13280 17080 13308
rect 16724 13268 16730 13280
rect 17310 13268 17316 13320
rect 17368 13268 17374 13320
rect 17586 13268 17592 13320
rect 17644 13268 17650 13320
rect 17788 13317 17816 13348
rect 18524 13317 18552 13416
rect 21910 13404 21916 13416
rect 21968 13404 21974 13456
rect 23382 13444 23388 13456
rect 23124 13416 23388 13444
rect 18598 13336 18604 13388
rect 18656 13336 18662 13388
rect 19978 13336 19984 13388
rect 20036 13336 20042 13388
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 18049 13311 18107 13317
rect 18049 13308 18061 13311
rect 17819 13280 18061 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 18049 13277 18061 13280
rect 18095 13277 18107 13311
rect 18049 13271 18107 13277
rect 18509 13311 18567 13317
rect 18509 13277 18521 13311
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 19886 13268 19892 13320
rect 19944 13308 19950 13320
rect 20070 13308 20076 13320
rect 19944 13280 20076 13308
rect 19944 13268 19950 13280
rect 20070 13268 20076 13280
rect 20128 13268 20134 13320
rect 21174 13268 21180 13320
rect 21232 13308 21238 13320
rect 23017 13311 23075 13317
rect 23017 13308 23029 13311
rect 21232 13280 23029 13308
rect 21232 13268 21238 13280
rect 23017 13277 23029 13280
rect 23063 13308 23075 13311
rect 23124 13308 23152 13416
rect 23382 13404 23388 13416
rect 23440 13404 23446 13456
rect 24394 13376 24400 13388
rect 23216 13348 24400 13376
rect 23216 13320 23244 13348
rect 24394 13336 24400 13348
rect 24452 13336 24458 13388
rect 24596 13376 24624 13475
rect 25774 13472 25780 13524
rect 25832 13512 25838 13524
rect 25961 13515 26019 13521
rect 25961 13512 25973 13515
rect 25832 13484 25973 13512
rect 25832 13472 25838 13484
rect 25961 13481 25973 13484
rect 26007 13481 26019 13515
rect 25961 13475 26019 13481
rect 26050 13472 26056 13524
rect 26108 13472 26114 13524
rect 26970 13472 26976 13524
rect 27028 13472 27034 13524
rect 24949 13447 25007 13453
rect 24949 13413 24961 13447
rect 24995 13444 25007 13447
rect 26068 13444 26096 13472
rect 24995 13416 26096 13444
rect 27341 13447 27399 13453
rect 24995 13413 25007 13416
rect 24949 13407 25007 13413
rect 27341 13413 27353 13447
rect 27387 13413 27399 13447
rect 27341 13407 27399 13413
rect 25501 13379 25559 13385
rect 25501 13376 25513 13379
rect 24596 13348 25513 13376
rect 25501 13345 25513 13348
rect 25547 13376 25559 13379
rect 25547 13348 26280 13376
rect 25547 13345 25559 13348
rect 25501 13339 25559 13345
rect 23063 13280 23152 13308
rect 23063 13277 23075 13280
rect 23017 13271 23075 13277
rect 23198 13268 23204 13320
rect 23256 13268 23262 13320
rect 23290 13268 23296 13320
rect 23348 13268 23354 13320
rect 23477 13311 23535 13317
rect 23477 13277 23489 13311
rect 23523 13308 23535 13311
rect 24026 13308 24032 13320
rect 23523 13280 24032 13308
rect 23523 13277 23535 13280
rect 23477 13271 23535 13277
rect 24026 13268 24032 13280
rect 24084 13268 24090 13320
rect 24854 13268 24860 13320
rect 24912 13268 24918 13320
rect 25038 13268 25044 13320
rect 25096 13268 25102 13320
rect 25590 13268 25596 13320
rect 25648 13268 25654 13320
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13308 25835 13311
rect 26142 13308 26148 13320
rect 25823 13280 26148 13308
rect 25823 13277 25835 13280
rect 25777 13271 25835 13277
rect 14185 13243 14243 13249
rect 14185 13240 14197 13243
rect 13872 13212 14197 13240
rect 13872 13200 13878 13212
rect 14185 13209 14197 13212
rect 14231 13209 14243 13243
rect 14660 13240 14688 13268
rect 15378 13240 15384 13252
rect 14660 13212 15384 13240
rect 14185 13203 14243 13209
rect 15378 13200 15384 13212
rect 15436 13200 15442 13252
rect 16758 13200 16764 13252
rect 16816 13200 16822 13252
rect 17604 13212 18092 13240
rect 10321 13175 10379 13181
rect 10321 13172 10333 13175
rect 10284 13144 10333 13172
rect 10284 13132 10290 13144
rect 10321 13141 10333 13144
rect 10367 13141 10379 13175
rect 10321 13135 10379 13141
rect 10410 13132 10416 13184
rect 10468 13172 10474 13184
rect 10689 13175 10747 13181
rect 10689 13172 10701 13175
rect 10468 13144 10701 13172
rect 10468 13132 10474 13144
rect 10689 13141 10701 13144
rect 10735 13172 10747 13175
rect 11146 13172 11152 13184
rect 10735 13144 11152 13172
rect 10735 13141 10747 13144
rect 10689 13135 10747 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11422 13132 11428 13184
rect 11480 13172 11486 13184
rect 12250 13172 12256 13184
rect 11480 13144 12256 13172
rect 11480 13132 11486 13144
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 14645 13175 14703 13181
rect 14645 13172 14657 13175
rect 13964 13144 14657 13172
rect 13964 13132 13970 13144
rect 14645 13141 14657 13144
rect 14691 13141 14703 13175
rect 14645 13135 14703 13141
rect 14734 13132 14740 13184
rect 14792 13132 14798 13184
rect 14826 13132 14832 13184
rect 14884 13172 14890 13184
rect 17604 13172 17632 13212
rect 14884 13144 17632 13172
rect 14884 13132 14890 13144
rect 17678 13132 17684 13184
rect 17736 13132 17742 13184
rect 18064 13172 18092 13212
rect 18138 13200 18144 13252
rect 18196 13240 18202 13252
rect 18233 13243 18291 13249
rect 18233 13240 18245 13243
rect 18196 13212 18245 13240
rect 18196 13200 18202 13212
rect 18233 13209 18245 13212
rect 18279 13240 18291 13243
rect 18322 13240 18328 13252
rect 18279 13212 18328 13240
rect 18279 13209 18291 13212
rect 18233 13203 18291 13209
rect 18322 13200 18328 13212
rect 18380 13200 18386 13252
rect 18414 13200 18420 13252
rect 18472 13240 18478 13252
rect 21266 13240 21272 13252
rect 18472 13212 21272 13240
rect 18472 13200 18478 13212
rect 21266 13200 21272 13212
rect 21324 13200 21330 13252
rect 22094 13200 22100 13252
rect 22152 13200 22158 13252
rect 22462 13200 22468 13252
rect 22520 13240 22526 13252
rect 24670 13249 24676 13252
rect 24397 13243 24455 13249
rect 24397 13240 24409 13243
rect 22520 13212 24409 13240
rect 22520 13200 22526 13212
rect 24397 13209 24409 13212
rect 24443 13209 24455 13243
rect 24397 13203 24455 13209
rect 24613 13243 24676 13249
rect 24613 13209 24625 13243
rect 24659 13209 24676 13243
rect 24613 13203 24676 13209
rect 24670 13200 24676 13203
rect 24728 13200 24734 13252
rect 25222 13200 25228 13252
rect 25280 13240 25286 13252
rect 25792 13240 25820 13271
rect 26142 13268 26148 13280
rect 26200 13268 26206 13320
rect 26252 13317 26280 13348
rect 26326 13336 26332 13388
rect 26384 13336 26390 13388
rect 27065 13379 27123 13385
rect 27065 13376 27077 13379
rect 26528 13348 27077 13376
rect 26237 13311 26295 13317
rect 26237 13277 26249 13311
rect 26283 13277 26295 13311
rect 26237 13271 26295 13277
rect 25280 13212 25820 13240
rect 25280 13200 25286 13212
rect 18966 13172 18972 13184
rect 18064 13144 18972 13172
rect 18966 13132 18972 13144
rect 19024 13132 19030 13184
rect 20257 13175 20315 13181
rect 20257 13141 20269 13175
rect 20303 13172 20315 13175
rect 21174 13172 21180 13184
rect 20303 13144 21180 13172
rect 20303 13141 20315 13144
rect 20257 13135 20315 13141
rect 21174 13132 21180 13144
rect 21232 13132 21238 13184
rect 22112 13172 22140 13200
rect 26528 13184 26556 13348
rect 27065 13345 27077 13348
rect 27111 13345 27123 13379
rect 27356 13376 27384 13407
rect 27356 13348 27660 13376
rect 27065 13339 27123 13345
rect 26973 13311 27031 13317
rect 26973 13308 26985 13311
rect 26620 13280 26985 13308
rect 26620 13184 26648 13280
rect 26973 13277 26985 13280
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 27430 13268 27436 13320
rect 27488 13268 27494 13320
rect 27632 13317 27660 13348
rect 27617 13311 27675 13317
rect 27617 13277 27629 13311
rect 27663 13277 27675 13311
rect 27617 13271 27675 13277
rect 22922 13172 22928 13184
rect 22112 13144 22928 13172
rect 22922 13132 22928 13144
rect 22980 13172 22986 13184
rect 23198 13172 23204 13184
rect 22980 13144 23204 13172
rect 22980 13132 22986 13144
rect 23198 13132 23204 13144
rect 23256 13132 23262 13184
rect 24029 13175 24087 13181
rect 24029 13141 24041 13175
rect 24075 13172 24087 13175
rect 24118 13172 24124 13184
rect 24075 13144 24124 13172
rect 24075 13141 24087 13144
rect 24029 13135 24087 13141
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 24762 13132 24768 13184
rect 24820 13132 24826 13184
rect 26510 13132 26516 13184
rect 26568 13132 26574 13184
rect 26602 13132 26608 13184
rect 26660 13132 26666 13184
rect 27798 13132 27804 13184
rect 27856 13132 27862 13184
rect 1104 13082 35236 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 35236 13082
rect 1104 13008 35236 13030
rect 9766 12968 9772 12980
rect 9048 12940 9772 12968
rect 9048 12909 9076 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 11146 12928 11152 12980
rect 11204 12928 11210 12980
rect 15194 12968 15200 12980
rect 11256 12940 12204 12968
rect 9033 12903 9091 12909
rect 9033 12869 9045 12903
rect 9079 12869 9091 12903
rect 9033 12863 9091 12869
rect 9214 12860 9220 12912
rect 9272 12909 9278 12912
rect 9272 12903 9291 12909
rect 9279 12869 9291 12903
rect 9272 12863 9291 12869
rect 9272 12860 9278 12863
rect 8757 12835 8815 12841
rect 8757 12801 8769 12835
rect 8803 12832 8815 12835
rect 8846 12832 8852 12844
rect 8803 12804 8852 12832
rect 8803 12801 8815 12804
rect 8757 12795 8815 12801
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 8938 12792 8944 12844
rect 8996 12792 9002 12844
rect 9677 12835 9735 12841
rect 9677 12832 9689 12835
rect 9232 12804 9689 12832
rect 9232 12637 9260 12804
rect 9677 12801 9689 12804
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12733 9551 12767
rect 9493 12727 9551 12733
rect 9508 12696 9536 12727
rect 9784 12696 9812 12928
rect 9858 12860 9864 12912
rect 9916 12860 9922 12912
rect 10686 12860 10692 12912
rect 10744 12900 10750 12912
rect 10965 12903 11023 12909
rect 10965 12900 10977 12903
rect 10744 12872 10977 12900
rect 10744 12860 10750 12872
rect 10965 12869 10977 12872
rect 11011 12900 11023 12903
rect 11256 12900 11284 12940
rect 11011 12872 11284 12900
rect 11011 12869 11023 12872
rect 10965 12863 11023 12869
rect 10321 12835 10379 12841
rect 10321 12801 10333 12835
rect 10367 12832 10379 12835
rect 10778 12832 10784 12844
rect 10367 12804 10784 12832
rect 10367 12801 10379 12804
rect 10321 12795 10379 12801
rect 10778 12792 10784 12804
rect 10836 12832 10842 12844
rect 10873 12835 10931 12841
rect 10873 12832 10885 12835
rect 10836 12804 10885 12832
rect 10836 12792 10842 12804
rect 10873 12801 10885 12804
rect 10919 12801 10931 12835
rect 11057 12835 11115 12841
rect 11057 12832 11069 12835
rect 10873 12795 10931 12801
rect 10980 12804 11069 12832
rect 9950 12724 9956 12776
rect 10008 12724 10014 12776
rect 10410 12724 10416 12776
rect 10468 12724 10474 12776
rect 10980 12696 11008 12804
rect 11057 12801 11069 12804
rect 11103 12801 11115 12835
rect 11057 12795 11115 12801
rect 11146 12792 11152 12844
rect 11204 12792 11210 12844
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 11422 12832 11428 12844
rect 11379 12804 11428 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 11422 12792 11428 12804
rect 11480 12792 11486 12844
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11701 12835 11759 12841
rect 11701 12801 11713 12835
rect 11747 12801 11759 12835
rect 11701 12795 11759 12801
rect 11532 12764 11560 12795
rect 11256 12736 11560 12764
rect 11256 12708 11284 12736
rect 9508 12668 11008 12696
rect 8941 12631 8999 12637
rect 8941 12597 8953 12631
rect 8987 12628 8999 12631
rect 9217 12631 9275 12637
rect 9217 12628 9229 12631
rect 8987 12600 9229 12628
rect 8987 12597 8999 12600
rect 8941 12591 8999 12597
rect 9217 12597 9229 12600
rect 9263 12597 9275 12631
rect 9217 12591 9275 12597
rect 9401 12631 9459 12637
rect 9401 12597 9413 12631
rect 9447 12628 9459 12631
rect 10042 12628 10048 12640
rect 9447 12600 10048 12628
rect 9447 12597 9459 12600
rect 9401 12591 9459 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 10980 12628 11008 12668
rect 11238 12656 11244 12708
rect 11296 12656 11302 12708
rect 11514 12656 11520 12708
rect 11572 12696 11578 12708
rect 11716 12696 11744 12795
rect 11790 12792 11796 12844
rect 11848 12832 11854 12844
rect 11977 12835 12035 12841
rect 11977 12832 11989 12835
rect 11848 12804 11989 12832
rect 11848 12792 11854 12804
rect 11977 12801 11989 12804
rect 12023 12801 12035 12835
rect 12176 12832 12204 12940
rect 14660 12940 15200 12968
rect 11977 12795 12035 12801
rect 12084 12804 12204 12832
rect 11808 12736 12020 12764
rect 11808 12705 11836 12736
rect 11992 12708 12020 12736
rect 11572 12668 11744 12696
rect 11793 12699 11851 12705
rect 11572 12656 11578 12668
rect 11793 12665 11805 12699
rect 11839 12665 11851 12699
rect 11793 12659 11851 12665
rect 11882 12656 11888 12708
rect 11940 12656 11946 12708
rect 11974 12656 11980 12708
rect 12032 12656 12038 12708
rect 12084 12696 12112 12804
rect 12250 12792 12256 12844
rect 12308 12792 12314 12844
rect 14366 12792 14372 12844
rect 14424 12832 14430 12844
rect 14660 12841 14688 12940
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 15378 12928 15384 12980
rect 15436 12928 15442 12980
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 16666 12928 16672 12980
rect 16724 12928 16730 12980
rect 19889 12971 19947 12977
rect 19889 12937 19901 12971
rect 19935 12968 19947 12971
rect 19978 12968 19984 12980
rect 19935 12940 19984 12968
rect 19935 12937 19947 12940
rect 19889 12931 19947 12937
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 26602 12928 26608 12980
rect 26660 12928 26666 12980
rect 26786 12928 26792 12980
rect 26844 12968 26850 12980
rect 27430 12968 27436 12980
rect 26844 12940 27436 12968
rect 26844 12928 26850 12940
rect 27430 12928 27436 12940
rect 27488 12928 27494 12980
rect 15396 12900 15424 12928
rect 15657 12903 15715 12909
rect 15657 12900 15669 12903
rect 15396 12872 15669 12900
rect 15657 12869 15669 12872
rect 15703 12900 15715 12903
rect 17586 12900 17592 12912
rect 15703 12872 17592 12900
rect 15703 12869 15715 12872
rect 15657 12863 15715 12869
rect 17236 12844 17264 12872
rect 17586 12860 17592 12872
rect 17644 12860 17650 12912
rect 19334 12860 19340 12912
rect 19392 12900 19398 12912
rect 19429 12903 19487 12909
rect 19429 12900 19441 12903
rect 19392 12872 19441 12900
rect 19392 12860 19398 12872
rect 19429 12869 19441 12872
rect 19475 12869 19487 12903
rect 19429 12863 19487 12869
rect 21913 12903 21971 12909
rect 21913 12869 21925 12903
rect 21959 12900 21971 12903
rect 22278 12900 22284 12912
rect 21959 12872 22284 12900
rect 21959 12869 21971 12872
rect 21913 12863 21971 12869
rect 22278 12860 22284 12872
rect 22336 12860 22342 12912
rect 14645 12835 14703 12841
rect 14645 12832 14657 12835
rect 14424 12804 14657 12832
rect 14424 12792 14430 12804
rect 14645 12801 14657 12804
rect 14691 12801 14703 12835
rect 14645 12795 14703 12801
rect 15838 12792 15844 12844
rect 15896 12792 15902 12844
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 16025 12835 16083 12841
rect 16025 12832 16037 12835
rect 15988 12804 16037 12832
rect 15988 12792 15994 12804
rect 16025 12801 16037 12804
rect 16071 12801 16083 12835
rect 16025 12795 16083 12801
rect 16776 12804 17172 12832
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12764 12219 12767
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 12207 12736 12541 12764
rect 12207 12733 12219 12736
rect 12161 12727 12219 12733
rect 12529 12733 12541 12736
rect 12575 12733 12587 12767
rect 12529 12727 12587 12733
rect 15194 12724 15200 12776
rect 15252 12724 15258 12776
rect 16776 12764 16804 12804
rect 16040 12736 16804 12764
rect 12084 12668 12388 12696
rect 11532 12628 11560 12656
rect 12360 12637 12388 12668
rect 14734 12656 14740 12708
rect 14792 12696 14798 12708
rect 15010 12696 15016 12708
rect 14792 12668 15016 12696
rect 14792 12656 14798 12668
rect 15010 12656 15016 12668
rect 15068 12656 15074 12708
rect 15105 12699 15163 12705
rect 15105 12665 15117 12699
rect 15151 12696 15163 12699
rect 15470 12696 15476 12708
rect 15151 12668 15476 12696
rect 15151 12665 15163 12668
rect 15105 12659 15163 12665
rect 15470 12656 15476 12668
rect 15528 12656 15534 12708
rect 10980 12600 11560 12628
rect 12345 12631 12403 12637
rect 12345 12597 12357 12631
rect 12391 12597 12403 12631
rect 12345 12591 12403 12597
rect 12805 12631 12863 12637
rect 12805 12597 12817 12631
rect 12851 12628 12863 12631
rect 16040 12628 16068 12736
rect 16850 12724 16856 12776
rect 16908 12764 16914 12776
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 16908 12736 17049 12764
rect 16908 12724 16914 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17144 12764 17172 12804
rect 17218 12792 17224 12844
rect 17276 12792 17282 12844
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17368 12804 17417 12832
rect 17368 12792 17374 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 18966 12792 18972 12844
rect 19024 12792 19030 12844
rect 26510 12832 26516 12844
rect 22066 12804 26516 12832
rect 17954 12764 17960 12776
rect 17144 12736 17960 12764
rect 17037 12727 17095 12733
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 21910 12724 21916 12776
rect 21968 12764 21974 12776
rect 22066 12764 22094 12804
rect 26510 12792 26516 12804
rect 26568 12792 26574 12844
rect 21968 12736 22094 12764
rect 26620 12764 26648 12928
rect 27893 12835 27951 12841
rect 27893 12801 27905 12835
rect 27939 12832 27951 12835
rect 28074 12832 28080 12844
rect 27939 12804 28080 12832
rect 27939 12801 27951 12804
rect 27893 12795 27951 12801
rect 28074 12792 28080 12804
rect 28132 12832 28138 12844
rect 28350 12832 28356 12844
rect 28132 12804 28356 12832
rect 28132 12792 28138 12804
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 26789 12767 26847 12773
rect 26789 12764 26801 12767
rect 26620 12736 26801 12764
rect 21968 12724 21974 12736
rect 26789 12733 26801 12736
rect 26835 12733 26847 12767
rect 26789 12727 26847 12733
rect 27798 12724 27804 12776
rect 27856 12724 27862 12776
rect 16666 12656 16672 12708
rect 16724 12696 16730 12708
rect 17129 12699 17187 12705
rect 17129 12696 17141 12699
rect 16724 12668 17141 12696
rect 16724 12656 16730 12668
rect 17129 12665 17141 12668
rect 17175 12665 17187 12699
rect 17129 12659 17187 12665
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 19705 12699 19763 12705
rect 19705 12696 19717 12699
rect 19484 12668 19717 12696
rect 19484 12656 19490 12668
rect 19705 12665 19717 12668
rect 19751 12665 19763 12699
rect 19705 12659 19763 12665
rect 22186 12656 22192 12708
rect 22244 12656 22250 12708
rect 12851 12600 16068 12628
rect 12851 12597 12863 12600
rect 12805 12591 12863 12597
rect 16574 12588 16580 12640
rect 16632 12628 16638 12640
rect 16945 12631 17003 12637
rect 16945 12628 16957 12631
rect 16632 12600 16957 12628
rect 16632 12588 16638 12600
rect 16945 12597 16957 12600
rect 16991 12597 17003 12631
rect 16945 12591 17003 12597
rect 19061 12631 19119 12637
rect 19061 12597 19073 12631
rect 19107 12628 19119 12631
rect 19334 12628 19340 12640
rect 19107 12600 19340 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19334 12588 19340 12600
rect 19392 12588 19398 12640
rect 22373 12631 22431 12637
rect 22373 12597 22385 12631
rect 22419 12628 22431 12631
rect 22646 12628 22652 12640
rect 22419 12600 22652 12628
rect 22419 12597 22431 12600
rect 22373 12591 22431 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 26605 12631 26663 12637
rect 26605 12597 26617 12631
rect 26651 12628 26663 12631
rect 26970 12628 26976 12640
rect 26651 12600 26976 12628
rect 26651 12597 26663 12600
rect 26605 12591 26663 12597
rect 26970 12588 26976 12600
rect 27028 12588 27034 12640
rect 28261 12631 28319 12637
rect 28261 12597 28273 12631
rect 28307 12628 28319 12631
rect 28534 12628 28540 12640
rect 28307 12600 28540 12628
rect 28307 12597 28319 12600
rect 28261 12591 28319 12597
rect 28534 12588 28540 12600
rect 28592 12588 28598 12640
rect 1104 12538 35248 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 35248 12538
rect 1104 12464 35248 12486
rect 9306 12384 9312 12436
rect 9364 12384 9370 12436
rect 10778 12384 10784 12436
rect 10836 12424 10842 12436
rect 11238 12424 11244 12436
rect 10836 12396 11244 12424
rect 10836 12384 10842 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11701 12427 11759 12433
rect 11701 12393 11713 12427
rect 11747 12424 11759 12427
rect 11882 12424 11888 12436
rect 11747 12396 11888 12424
rect 11747 12393 11759 12396
rect 11701 12387 11759 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12069 12427 12127 12433
rect 12069 12393 12081 12427
rect 12115 12424 12127 12427
rect 12250 12424 12256 12436
rect 12115 12396 12256 12424
rect 12115 12393 12127 12396
rect 12069 12387 12127 12393
rect 12250 12384 12256 12396
rect 12308 12384 12314 12436
rect 15013 12427 15071 12433
rect 15013 12393 15025 12427
rect 15059 12424 15071 12427
rect 15102 12424 15108 12436
rect 15059 12396 15108 12424
rect 15059 12393 15071 12396
rect 15013 12387 15071 12393
rect 15102 12384 15108 12396
rect 15160 12384 15166 12436
rect 15933 12427 15991 12433
rect 15933 12424 15945 12427
rect 15488 12396 15945 12424
rect 9677 12359 9735 12365
rect 9677 12356 9689 12359
rect 9324 12328 9689 12356
rect 9324 12232 9352 12328
rect 9677 12325 9689 12328
rect 9723 12325 9735 12359
rect 9677 12319 9735 12325
rect 9769 12359 9827 12365
rect 9769 12325 9781 12359
rect 9815 12356 9827 12359
rect 9858 12356 9864 12368
rect 9815 12328 9864 12356
rect 9815 12325 9827 12328
rect 9769 12319 9827 12325
rect 9858 12316 9864 12328
rect 9916 12316 9922 12368
rect 11054 12316 11060 12368
rect 11112 12356 11118 12368
rect 11606 12356 11612 12368
rect 11112 12328 11612 12356
rect 11112 12316 11118 12328
rect 11606 12316 11612 12328
rect 11664 12316 11670 12368
rect 11790 12316 11796 12368
rect 11848 12316 11854 12368
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 11808 12288 11836 12316
rect 9640 12260 11100 12288
rect 9640 12248 9646 12260
rect 11072 12232 11100 12260
rect 11440 12260 11836 12288
rect 11900 12288 11928 12384
rect 15488 12368 15516 12396
rect 15933 12393 15945 12396
rect 15979 12424 15991 12427
rect 15979 12396 16344 12424
rect 15979 12393 15991 12396
rect 15933 12387 15991 12393
rect 15470 12356 15476 12368
rect 15028 12328 15476 12356
rect 11900 12260 12112 12288
rect 11440 12232 11468 12260
rect 9306 12180 9312 12232
rect 9364 12180 9370 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 10137 12223 10195 12229
rect 10137 12220 10149 12223
rect 9824 12192 10149 12220
rect 9824 12180 9830 12192
rect 10137 12189 10149 12192
rect 10183 12220 10195 12223
rect 10410 12220 10416 12232
rect 10183 12192 10416 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11054 12180 11060 12232
rect 11112 12180 11118 12232
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11296 12192 11345 12220
rect 11296 12180 11302 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11422 12180 11428 12232
rect 11480 12180 11486 12232
rect 11514 12180 11520 12232
rect 11572 12180 11578 12232
rect 11624 12229 11652 12260
rect 11609 12223 11667 12229
rect 11609 12189 11621 12223
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12220 11851 12223
rect 11974 12220 11980 12232
rect 11839 12192 11980 12220
rect 11839 12189 11851 12192
rect 11793 12183 11851 12189
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10704 12124 10885 12152
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9858 12084 9864 12096
rect 9456 12056 9864 12084
rect 9456 12044 9462 12056
rect 9858 12044 9864 12056
rect 9916 12084 9922 12096
rect 10226 12084 10232 12096
rect 9916 12056 10232 12084
rect 9916 12044 9922 12056
rect 10226 12044 10232 12056
rect 10284 12084 10290 12096
rect 10704 12093 10732 12124
rect 10873 12121 10885 12124
rect 10919 12121 10931 12155
rect 11808 12152 11836 12183
rect 11974 12180 11980 12192
rect 12032 12180 12038 12232
rect 10873 12115 10931 12121
rect 11256 12124 11836 12152
rect 11256 12096 11284 12124
rect 10689 12087 10747 12093
rect 10689 12084 10701 12087
rect 10284 12056 10701 12084
rect 10284 12044 10290 12056
rect 10689 12053 10701 12056
rect 10735 12053 10747 12087
rect 10689 12047 10747 12053
rect 11238 12044 11244 12096
rect 11296 12044 11302 12096
rect 12084 12084 12112 12260
rect 14458 12248 14464 12300
rect 14516 12288 14522 12300
rect 14516 12260 14688 12288
rect 14516 12248 14522 12260
rect 12342 12180 12348 12232
rect 12400 12220 12406 12232
rect 13265 12223 13323 12229
rect 13265 12220 13277 12223
rect 12400 12192 13277 12220
rect 12400 12180 12406 12192
rect 13265 12189 13277 12192
rect 13311 12189 13323 12223
rect 13265 12183 13323 12189
rect 13280 12152 13308 12183
rect 13354 12180 13360 12232
rect 13412 12220 13418 12232
rect 13449 12223 13507 12229
rect 13449 12220 13461 12223
rect 13412 12192 13461 12220
rect 13412 12180 13418 12192
rect 13449 12189 13461 12192
rect 13495 12189 13507 12223
rect 13449 12183 13507 12189
rect 13814 12180 13820 12232
rect 13872 12180 13878 12232
rect 14200 12192 14504 12220
rect 13832 12152 13860 12180
rect 14200 12164 14228 12192
rect 13280 12124 13860 12152
rect 14182 12112 14188 12164
rect 14240 12112 14246 12164
rect 14366 12112 14372 12164
rect 14424 12112 14430 12164
rect 14476 12161 14504 12192
rect 14461 12155 14519 12161
rect 14461 12121 14473 12155
rect 14507 12121 14519 12155
rect 14660 12152 14688 12260
rect 15028 12232 15056 12328
rect 15470 12316 15476 12328
rect 15528 12316 15534 12368
rect 15838 12316 15844 12368
rect 15896 12356 15902 12368
rect 15896 12328 16252 12356
rect 15896 12316 15902 12328
rect 16022 12288 16028 12300
rect 15120 12260 16028 12288
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 15010 12220 15016 12232
rect 14875 12192 15016 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 15120 12152 15148 12260
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 16224 12232 16252 12328
rect 16206 12180 16212 12232
rect 16264 12180 16270 12232
rect 16316 12220 16344 12396
rect 16390 12384 16396 12436
rect 16448 12384 16454 12436
rect 16485 12427 16543 12433
rect 16485 12393 16497 12427
rect 16531 12424 16543 12427
rect 16758 12424 16764 12436
rect 16531 12396 16764 12424
rect 16531 12393 16543 12396
rect 16485 12387 16543 12393
rect 16758 12384 16764 12396
rect 16816 12384 16822 12436
rect 19245 12427 19303 12433
rect 19245 12393 19257 12427
rect 19291 12424 19303 12427
rect 20070 12424 20076 12436
rect 19291 12396 20076 12424
rect 19291 12393 19303 12396
rect 19245 12387 19303 12393
rect 20070 12384 20076 12396
rect 20128 12384 20134 12436
rect 22278 12384 22284 12436
rect 22336 12384 22342 12436
rect 25774 12384 25780 12436
rect 25832 12384 25838 12436
rect 26326 12384 26332 12436
rect 26384 12424 26390 12436
rect 26513 12427 26571 12433
rect 26513 12424 26525 12427
rect 26384 12396 26525 12424
rect 26384 12384 26390 12396
rect 26513 12393 26525 12396
rect 26559 12393 26571 12427
rect 26513 12387 26571 12393
rect 16408 12288 16436 12384
rect 16574 12316 16580 12368
rect 16632 12356 16638 12368
rect 16853 12359 16911 12365
rect 16853 12356 16865 12359
rect 16632 12328 16865 12356
rect 16632 12316 16638 12328
rect 16853 12325 16865 12328
rect 16899 12325 16911 12359
rect 28258 12356 28264 12368
rect 16853 12319 16911 12325
rect 18340 12328 19656 12356
rect 18340 12297 18368 12328
rect 17221 12291 17279 12297
rect 17221 12288 17233 12291
rect 16408 12260 17233 12288
rect 17221 12257 17233 12260
rect 17267 12257 17279 12291
rect 18325 12291 18383 12297
rect 17221 12251 17279 12257
rect 17328 12260 18184 12288
rect 16390 12220 16396 12232
rect 16316 12192 16396 12220
rect 16390 12180 16396 12192
rect 16448 12220 16454 12232
rect 16666 12220 16672 12232
rect 16448 12192 16672 12220
rect 16448 12180 16454 12192
rect 16666 12180 16672 12192
rect 16724 12180 16730 12232
rect 16761 12223 16819 12229
rect 16761 12189 16773 12223
rect 16807 12220 16819 12223
rect 16850 12220 16856 12232
rect 16807 12192 16856 12220
rect 16807 12189 16819 12192
rect 16761 12183 16819 12189
rect 16850 12180 16856 12192
rect 16908 12180 16914 12232
rect 16942 12180 16948 12232
rect 17000 12180 17006 12232
rect 17126 12180 17132 12232
rect 17184 12180 17190 12232
rect 14660 12124 15148 12152
rect 14461 12115 14519 12121
rect 15838 12112 15844 12164
rect 15896 12152 15902 12164
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 15896 12124 15945 12152
rect 15896 12112 15902 12124
rect 15933 12121 15945 12124
rect 15979 12152 15991 12155
rect 16574 12152 16580 12164
rect 15979 12124 16580 12152
rect 15979 12121 15991 12124
rect 15933 12115 15991 12121
rect 16574 12112 16580 12124
rect 16632 12112 16638 12164
rect 16868 12152 16896 12180
rect 17328 12152 17356 12260
rect 17402 12180 17408 12232
rect 17460 12180 17466 12232
rect 18156 12229 18184 12260
rect 18325 12257 18337 12291
rect 18371 12257 18383 12291
rect 18325 12251 18383 12257
rect 18969 12291 19027 12297
rect 18969 12257 18981 12291
rect 19015 12288 19027 12291
rect 19015 12260 19564 12288
rect 19015 12257 19027 12260
rect 18969 12251 19027 12257
rect 17957 12223 18015 12229
rect 17957 12220 17969 12223
rect 17512 12192 17969 12220
rect 16868 12124 17356 12152
rect 13357 12087 13415 12093
rect 13357 12084 13369 12087
rect 12084 12056 13369 12084
rect 13357 12053 13369 12056
rect 13403 12084 13415 12087
rect 17512 12084 17540 12192
rect 17957 12189 17969 12192
rect 18003 12189 18015 12223
rect 17957 12183 18015 12189
rect 18141 12223 18199 12229
rect 18141 12189 18153 12223
rect 18187 12220 18199 12223
rect 18187 12192 18644 12220
rect 18187 12189 18199 12192
rect 18141 12183 18199 12189
rect 17972 12152 18000 12183
rect 18616 12161 18644 12192
rect 18782 12180 18788 12232
rect 18840 12180 18846 12232
rect 18874 12180 18880 12232
rect 18932 12180 18938 12232
rect 19061 12223 19119 12229
rect 19061 12189 19073 12223
rect 19107 12220 19119 12223
rect 19107 12192 19380 12220
rect 19107 12189 19119 12192
rect 19061 12183 19119 12189
rect 18417 12155 18475 12161
rect 18417 12152 18429 12155
rect 17972 12124 18429 12152
rect 18417 12121 18429 12124
rect 18463 12121 18475 12155
rect 18417 12115 18475 12121
rect 18601 12155 18659 12161
rect 18601 12121 18613 12155
rect 18647 12121 18659 12155
rect 18601 12115 18659 12121
rect 18690 12112 18696 12164
rect 18748 12152 18754 12164
rect 19245 12155 19303 12161
rect 19245 12152 19257 12155
rect 18748 12124 19257 12152
rect 18748 12112 18754 12124
rect 19245 12121 19257 12124
rect 19291 12121 19303 12155
rect 19245 12115 19303 12121
rect 13403 12056 17540 12084
rect 13403 12053 13415 12056
rect 13357 12047 13415 12053
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 19352 12084 19380 12192
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19536 12229 19564 12260
rect 19521 12223 19579 12229
rect 19521 12220 19533 12223
rect 19484 12192 19533 12220
rect 19484 12180 19490 12192
rect 19521 12189 19533 12192
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 17644 12056 19380 12084
rect 19429 12087 19487 12093
rect 17644 12044 17650 12056
rect 19429 12053 19441 12087
rect 19475 12084 19487 12087
rect 19628 12084 19656 12328
rect 28000 12328 28264 12356
rect 22373 12291 22431 12297
rect 22373 12257 22385 12291
rect 22419 12288 22431 12291
rect 23198 12288 23204 12300
rect 22419 12260 23204 12288
rect 22419 12257 22431 12260
rect 22373 12251 22431 12257
rect 22097 12223 22155 12229
rect 22097 12189 22109 12223
rect 22143 12220 22155 12223
rect 22186 12220 22192 12232
rect 22143 12192 22192 12220
rect 22143 12189 22155 12192
rect 22097 12183 22155 12189
rect 22186 12180 22192 12192
rect 22244 12180 22250 12232
rect 22646 12180 22652 12232
rect 22704 12180 22710 12232
rect 23032 12229 23060 12260
rect 23198 12248 23204 12260
rect 23256 12288 23262 12300
rect 23845 12291 23903 12297
rect 23845 12288 23857 12291
rect 23256 12260 23857 12288
rect 23256 12248 23262 12260
rect 23845 12257 23857 12260
rect 23891 12257 23903 12291
rect 25225 12291 25283 12297
rect 25225 12288 25237 12291
rect 23845 12251 23903 12257
rect 24596 12260 25237 12288
rect 23017 12223 23075 12229
rect 23017 12189 23029 12223
rect 23063 12189 23075 12223
rect 23017 12183 23075 12189
rect 23106 12180 23112 12232
rect 23164 12220 23170 12232
rect 23753 12223 23811 12229
rect 23753 12220 23765 12223
rect 23164 12192 23765 12220
rect 23164 12180 23170 12192
rect 23753 12189 23765 12192
rect 23799 12189 23811 12223
rect 23753 12183 23811 12189
rect 23937 12223 23995 12229
rect 23937 12189 23949 12223
rect 23983 12189 23995 12223
rect 23937 12183 23995 12189
rect 22554 12112 22560 12164
rect 22612 12152 22618 12164
rect 23952 12152 23980 12183
rect 24302 12180 24308 12232
rect 24360 12220 24366 12232
rect 24596 12229 24624 12260
rect 25225 12257 25237 12260
rect 25271 12257 25283 12291
rect 25225 12251 25283 12257
rect 24581 12223 24639 12229
rect 24581 12220 24593 12223
rect 24360 12192 24593 12220
rect 24360 12180 24366 12192
rect 24581 12189 24593 12192
rect 24627 12189 24639 12223
rect 24581 12183 24639 12189
rect 24762 12180 24768 12232
rect 24820 12220 24826 12232
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 24820 12192 25053 12220
rect 24820 12180 24826 12192
rect 25041 12189 25053 12192
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 25498 12180 25504 12232
rect 25556 12220 25562 12232
rect 25593 12223 25651 12229
rect 25593 12220 25605 12223
rect 25556 12192 25605 12220
rect 25556 12180 25562 12192
rect 25593 12189 25605 12192
rect 25639 12189 25651 12223
rect 25593 12183 25651 12189
rect 25777 12223 25835 12229
rect 25777 12189 25789 12223
rect 25823 12189 25835 12223
rect 25777 12183 25835 12189
rect 25792 12152 25820 12183
rect 26142 12180 26148 12232
rect 26200 12180 26206 12232
rect 26326 12180 26332 12232
rect 26384 12180 26390 12232
rect 27798 12180 27804 12232
rect 27856 12180 27862 12232
rect 27893 12223 27951 12229
rect 27893 12189 27905 12223
rect 27939 12220 27951 12223
rect 28000 12220 28028 12328
rect 28258 12316 28264 12328
rect 28316 12356 28322 12368
rect 28721 12359 28779 12365
rect 28721 12356 28733 12359
rect 28316 12328 28733 12356
rect 28316 12316 28322 12328
rect 28721 12325 28733 12328
rect 28767 12325 28779 12359
rect 28721 12319 28779 12325
rect 29089 12291 29147 12297
rect 29089 12288 29101 12291
rect 28460 12260 29101 12288
rect 27939 12192 28028 12220
rect 27939 12189 27951 12192
rect 27893 12183 27951 12189
rect 28074 12180 28080 12232
rect 28132 12220 28138 12232
rect 28169 12223 28227 12229
rect 28169 12220 28181 12223
rect 28132 12192 28181 12220
rect 28132 12180 28138 12192
rect 28169 12189 28181 12192
rect 28215 12220 28227 12223
rect 28261 12223 28319 12229
rect 28261 12220 28273 12223
rect 28215 12192 28273 12220
rect 28215 12189 28227 12192
rect 28169 12183 28227 12189
rect 28261 12189 28273 12192
rect 28307 12189 28319 12223
rect 28261 12183 28319 12189
rect 28350 12180 28356 12232
rect 28408 12220 28414 12232
rect 28460 12229 28488 12260
rect 29089 12257 29101 12260
rect 29135 12257 29147 12291
rect 29089 12251 29147 12257
rect 28445 12223 28503 12229
rect 28445 12220 28457 12223
rect 28408 12192 28457 12220
rect 28408 12180 28414 12192
rect 28445 12189 28457 12192
rect 28491 12189 28503 12223
rect 28445 12183 28503 12189
rect 28905 12223 28963 12229
rect 28905 12189 28917 12223
rect 28951 12189 28963 12223
rect 28905 12183 28963 12189
rect 22612 12124 23980 12152
rect 25608 12124 25820 12152
rect 27816 12152 27844 12180
rect 28629 12155 28687 12161
rect 28629 12152 28641 12155
rect 27816 12124 28641 12152
rect 22612 12112 22618 12124
rect 25608 12096 25636 12124
rect 28629 12121 28641 12124
rect 28675 12152 28687 12155
rect 28920 12152 28948 12183
rect 28675 12124 28948 12152
rect 28675 12121 28687 12124
rect 28629 12115 28687 12121
rect 19978 12084 19984 12096
rect 19475 12056 19984 12084
rect 19475 12053 19487 12056
rect 19429 12047 19487 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 21913 12087 21971 12093
rect 21913 12053 21925 12087
rect 21959 12084 21971 12087
rect 23566 12084 23572 12096
rect 21959 12056 23572 12084
rect 21959 12053 21971 12056
rect 21913 12047 21971 12053
rect 23566 12044 23572 12056
rect 23624 12044 23630 12096
rect 23661 12087 23719 12093
rect 23661 12053 23673 12087
rect 23707 12084 23719 12087
rect 24302 12084 24308 12096
rect 23707 12056 24308 12084
rect 23707 12053 23719 12056
rect 23661 12047 23719 12053
rect 24302 12044 24308 12056
rect 24360 12044 24366 12096
rect 24397 12087 24455 12093
rect 24397 12053 24409 12087
rect 24443 12084 24455 12087
rect 24578 12084 24584 12096
rect 24443 12056 24584 12084
rect 24443 12053 24455 12056
rect 24397 12047 24455 12053
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 24854 12044 24860 12096
rect 24912 12044 24918 12096
rect 25590 12044 25596 12096
rect 25648 12044 25654 12096
rect 27706 12044 27712 12096
rect 27764 12044 27770 12096
rect 27890 12044 27896 12096
rect 27948 12084 27954 12096
rect 28077 12087 28135 12093
rect 28077 12084 28089 12087
rect 27948 12056 28089 12084
rect 27948 12044 27954 12056
rect 28077 12053 28089 12056
rect 28123 12053 28135 12087
rect 28077 12047 28135 12053
rect 1104 11994 35236 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 35236 11994
rect 1104 11920 35236 11942
rect 9214 11840 9220 11892
rect 9272 11880 9278 11892
rect 9309 11883 9367 11889
rect 9309 11880 9321 11883
rect 9272 11852 9321 11880
rect 9272 11840 9278 11852
rect 9309 11849 9321 11852
rect 9355 11849 9367 11883
rect 9309 11843 9367 11849
rect 9582 11840 9588 11892
rect 9640 11840 9646 11892
rect 11146 11840 11152 11892
rect 11204 11880 11210 11892
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11204 11852 11989 11880
rect 11204 11840 11210 11852
rect 11977 11849 11989 11852
rect 12023 11849 12035 11883
rect 11977 11843 12035 11849
rect 9600 11753 9628 11840
rect 9784 11784 11008 11812
rect 9784 11756 9812 11784
rect 9585 11747 9643 11753
rect 9585 11713 9597 11747
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 9677 11747 9735 11753
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 9217 11679 9275 11685
rect 9217 11645 9229 11679
rect 9263 11676 9275 11679
rect 9398 11676 9404 11688
rect 9263 11648 9404 11676
rect 9263 11645 9275 11648
rect 9217 11639 9275 11645
rect 9398 11636 9404 11648
rect 9456 11676 9462 11688
rect 9692 11676 9720 11707
rect 9766 11704 9772 11756
rect 9824 11704 9830 11756
rect 9950 11704 9956 11756
rect 10008 11704 10014 11756
rect 10413 11747 10471 11753
rect 10413 11713 10425 11747
rect 10459 11744 10471 11747
rect 10778 11744 10784 11756
rect 10459 11716 10784 11744
rect 10459 11713 10471 11716
rect 10413 11707 10471 11713
rect 10778 11704 10784 11716
rect 10836 11704 10842 11756
rect 9456 11648 9720 11676
rect 9456 11636 9462 11648
rect 10502 11636 10508 11688
rect 10560 11636 10566 11688
rect 10980 11617 11008 11784
rect 11072 11784 11836 11812
rect 11072 11756 11100 11784
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 11808 11753 11836 11784
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 11296 11716 11529 11744
rect 11296 11704 11302 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 11517 11707 11575 11713
rect 11793 11747 11851 11753
rect 11793 11713 11805 11747
rect 11839 11713 11851 11747
rect 11992 11744 12020 11843
rect 14182 11840 14188 11892
rect 14240 11840 14246 11892
rect 14461 11883 14519 11889
rect 14461 11849 14473 11883
rect 14507 11880 14519 11883
rect 17402 11880 17408 11892
rect 14507 11852 17408 11880
rect 14507 11849 14519 11852
rect 14461 11843 14519 11849
rect 17402 11840 17408 11852
rect 17460 11840 17466 11892
rect 17586 11840 17592 11892
rect 17644 11840 17650 11892
rect 18417 11883 18475 11889
rect 18417 11849 18429 11883
rect 18463 11880 18475 11883
rect 18690 11880 18696 11892
rect 18463 11852 18696 11880
rect 18463 11849 18475 11852
rect 18417 11843 18475 11849
rect 18690 11840 18696 11852
rect 18748 11840 18754 11892
rect 18782 11840 18788 11892
rect 18840 11840 18846 11892
rect 19978 11840 19984 11892
rect 20036 11840 20042 11892
rect 22373 11883 22431 11889
rect 22373 11849 22385 11883
rect 22419 11880 22431 11883
rect 22419 11852 22692 11880
rect 22419 11849 22431 11852
rect 22373 11843 22431 11849
rect 14200 11812 14228 11840
rect 14200 11784 15056 11812
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11992 11716 12081 11744
rect 11793 11707 11851 11713
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12069 11707 12127 11713
rect 11606 11636 11612 11688
rect 11664 11636 11670 11688
rect 11808 11676 11836 11707
rect 12158 11704 12164 11756
rect 12216 11744 12222 11756
rect 12253 11747 12311 11753
rect 12253 11744 12265 11747
rect 12216 11716 12265 11744
rect 12216 11704 12222 11716
rect 12253 11713 12265 11716
rect 12299 11713 12311 11747
rect 12253 11707 12311 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 14185 11747 14243 11753
rect 12483 11716 14044 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 13354 11676 13360 11688
rect 11808 11648 13360 11676
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 13814 11636 13820 11688
rect 13872 11636 13878 11688
rect 13909 11679 13967 11685
rect 13909 11645 13921 11679
rect 13955 11645 13967 11679
rect 13909 11639 13967 11645
rect 10965 11611 11023 11617
rect 9324 11580 10916 11608
rect 9324 11552 9352 11580
rect 9306 11500 9312 11552
rect 9364 11500 9370 11552
rect 10137 11543 10195 11549
rect 10137 11509 10149 11543
rect 10183 11540 10195 11543
rect 10226 11540 10232 11552
rect 10183 11512 10232 11540
rect 10183 11509 10195 11512
rect 10137 11503 10195 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 10888 11540 10916 11580
rect 10965 11577 10977 11611
rect 11011 11608 11023 11611
rect 11333 11611 11391 11617
rect 11333 11608 11345 11611
rect 11011 11580 11345 11608
rect 11011 11577 11023 11580
rect 10965 11571 11023 11577
rect 11333 11577 11345 11580
rect 11379 11608 11391 11611
rect 11379 11580 11744 11608
rect 11379 11577 11391 11580
rect 11333 11571 11391 11577
rect 11716 11552 11744 11580
rect 11514 11540 11520 11552
rect 10888 11512 11520 11540
rect 11514 11500 11520 11512
rect 11572 11500 11578 11552
rect 11698 11500 11704 11552
rect 11756 11540 11762 11552
rect 12618 11540 12624 11552
rect 11756 11512 12624 11540
rect 11756 11500 11762 11512
rect 12618 11500 12624 11512
rect 12676 11540 12682 11552
rect 13630 11540 13636 11552
rect 12676 11512 13636 11540
rect 12676 11500 12682 11512
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13924 11540 13952 11639
rect 14016 11608 14044 11716
rect 14185 11713 14197 11747
rect 14231 11744 14243 11747
rect 14458 11744 14464 11756
rect 14231 11716 14464 11744
rect 14231 11713 14243 11716
rect 14185 11707 14243 11713
rect 14458 11704 14464 11716
rect 14516 11704 14522 11756
rect 15028 11753 15056 11784
rect 16022 11772 16028 11824
rect 16080 11812 16086 11824
rect 16080 11784 16896 11812
rect 16080 11772 16086 11784
rect 15013 11747 15071 11753
rect 15013 11713 15025 11747
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 16298 11704 16304 11756
rect 16356 11744 16362 11756
rect 16868 11753 16896 11784
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 16356 11716 16681 11744
rect 16356 11704 16362 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 16853 11747 16911 11753
rect 16853 11713 16865 11747
rect 16899 11713 16911 11747
rect 17604 11744 17632 11840
rect 18325 11747 18383 11753
rect 18325 11744 18337 11747
rect 17604 11716 18337 11744
rect 16853 11707 16911 11713
rect 18325 11713 18337 11716
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 18509 11747 18567 11753
rect 18509 11713 18521 11747
rect 18555 11713 18567 11747
rect 18800 11744 18828 11840
rect 19996 11753 20024 11840
rect 22664 11812 22692 11852
rect 23106 11840 23112 11892
rect 23164 11840 23170 11892
rect 23198 11840 23204 11892
rect 23256 11840 23262 11892
rect 23566 11840 23572 11892
rect 23624 11840 23630 11892
rect 24854 11840 24860 11892
rect 24912 11840 24918 11892
rect 26326 11840 26332 11892
rect 26384 11880 26390 11892
rect 26513 11883 26571 11889
rect 26513 11880 26525 11883
rect 26384 11852 26525 11880
rect 26384 11840 26390 11852
rect 26513 11849 26525 11852
rect 26559 11849 26571 11883
rect 28074 11880 28080 11892
rect 26513 11843 26571 11849
rect 27816 11852 28080 11880
rect 23124 11812 23152 11840
rect 22664 11784 23152 11812
rect 19245 11747 19303 11753
rect 19245 11744 19257 11747
rect 18800 11716 19257 11744
rect 18509 11707 18567 11713
rect 19245 11713 19257 11716
rect 19291 11713 19303 11747
rect 19245 11707 19303 11713
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11744 19487 11747
rect 19981 11747 20039 11753
rect 19981 11744 19993 11747
rect 19475 11716 19993 11744
rect 19475 11713 19487 11716
rect 19429 11707 19487 11713
rect 19981 11713 19993 11716
rect 20027 11744 20039 11747
rect 20441 11747 20499 11753
rect 20441 11744 20453 11747
rect 20027 11716 20453 11744
rect 20027 11713 20039 11716
rect 19981 11707 20039 11713
rect 20441 11713 20453 11716
rect 20487 11713 20499 11747
rect 20441 11707 20499 11713
rect 14277 11679 14335 11685
rect 14277 11645 14289 11679
rect 14323 11676 14335 11679
rect 15102 11676 15108 11688
rect 14323 11648 15108 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 16868 11676 16896 11707
rect 18414 11676 18420 11688
rect 16868 11648 18420 11676
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 18524 11676 18552 11707
rect 21634 11704 21640 11756
rect 21692 11744 21698 11756
rect 22005 11747 22063 11753
rect 22005 11744 22017 11747
rect 21692 11716 22017 11744
rect 21692 11704 21698 11716
rect 22005 11713 22017 11716
rect 22051 11713 22063 11747
rect 22005 11707 22063 11713
rect 22554 11704 22560 11756
rect 22612 11704 22618 11756
rect 22664 11753 22692 11784
rect 23216 11753 23244 11840
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11713 22707 11747
rect 22649 11707 22707 11713
rect 22833 11747 22891 11753
rect 22833 11713 22845 11747
rect 22879 11744 22891 11747
rect 23017 11747 23075 11753
rect 23017 11744 23029 11747
rect 22879 11716 23029 11744
rect 22879 11713 22891 11716
rect 22833 11707 22891 11713
rect 23017 11713 23029 11716
rect 23063 11713 23075 11747
rect 23017 11707 23075 11713
rect 23201 11747 23259 11753
rect 23201 11713 23213 11747
rect 23247 11713 23259 11747
rect 23584 11744 23612 11840
rect 24872 11812 24900 11840
rect 24504 11784 24900 11812
rect 25516 11784 26372 11812
rect 24504 11753 24532 11784
rect 25516 11756 25544 11784
rect 24397 11747 24455 11753
rect 24397 11744 24409 11747
rect 23584 11716 24409 11744
rect 23201 11707 23259 11713
rect 24397 11713 24409 11716
rect 24443 11713 24455 11747
rect 24397 11707 24455 11713
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 18874 11676 18880 11688
rect 18524 11648 18880 11676
rect 18524 11608 18552 11648
rect 18874 11636 18880 11648
rect 18932 11636 18938 11688
rect 19889 11679 19947 11685
rect 19889 11676 19901 11679
rect 19628 11648 19901 11676
rect 14016 11580 18552 11608
rect 19628 11552 19656 11648
rect 19889 11645 19901 11648
rect 19935 11676 19947 11679
rect 20349 11679 20407 11685
rect 20349 11676 20361 11679
rect 19935 11648 20361 11676
rect 19935 11645 19947 11648
rect 19889 11639 19947 11645
rect 20349 11645 20361 11648
rect 20395 11645 20407 11679
rect 20349 11639 20407 11645
rect 21726 11636 21732 11688
rect 21784 11676 21790 11688
rect 21913 11679 21971 11685
rect 21913 11676 21925 11679
rect 21784 11648 21925 11676
rect 21784 11636 21790 11648
rect 21913 11645 21925 11648
rect 21959 11676 21971 11679
rect 24412 11676 24440 11707
rect 24578 11704 24584 11756
rect 24636 11744 24642 11756
rect 24673 11747 24731 11753
rect 24673 11744 24685 11747
rect 24636 11716 24685 11744
rect 24636 11704 24642 11716
rect 24673 11713 24685 11716
rect 24719 11744 24731 11747
rect 25130 11744 25136 11756
rect 24719 11716 25136 11744
rect 24719 11713 24731 11716
rect 24673 11707 24731 11713
rect 25130 11704 25136 11716
rect 25188 11704 25194 11756
rect 25225 11747 25283 11753
rect 25225 11713 25237 11747
rect 25271 11713 25283 11747
rect 25225 11707 25283 11713
rect 25240 11676 25268 11707
rect 25498 11704 25504 11756
rect 25556 11704 25562 11756
rect 25590 11704 25596 11756
rect 25648 11744 25654 11756
rect 26344 11753 26372 11784
rect 27816 11753 27844 11852
rect 28074 11840 28080 11852
rect 28132 11840 28138 11892
rect 28166 11840 28172 11892
rect 28224 11840 28230 11892
rect 28258 11840 28264 11892
rect 28316 11840 28322 11892
rect 28184 11812 28212 11840
rect 28092 11784 28212 11812
rect 26145 11747 26203 11753
rect 26145 11744 26157 11747
rect 25648 11716 26157 11744
rect 25648 11704 25654 11716
rect 26145 11713 26157 11716
rect 26191 11713 26203 11747
rect 26145 11707 26203 11713
rect 26329 11747 26387 11753
rect 26329 11713 26341 11747
rect 26375 11713 26387 11747
rect 26329 11707 26387 11713
rect 27801 11747 27859 11753
rect 27801 11713 27813 11747
rect 27847 11713 27859 11747
rect 27801 11707 27859 11713
rect 27890 11704 27896 11756
rect 27948 11704 27954 11756
rect 28092 11753 28120 11784
rect 28077 11747 28135 11753
rect 28077 11713 28089 11747
rect 28123 11713 28135 11747
rect 28077 11707 28135 11713
rect 28169 11747 28227 11753
rect 28169 11713 28181 11747
rect 28215 11744 28227 11747
rect 28276 11744 28304 11840
rect 28629 11747 28687 11753
rect 28629 11744 28641 11747
rect 28215 11716 28304 11744
rect 28460 11716 28641 11744
rect 28215 11713 28227 11716
rect 28169 11707 28227 11713
rect 21959 11648 22094 11676
rect 24412 11648 25268 11676
rect 21959 11645 21971 11648
rect 21913 11639 21971 11645
rect 22066 11608 22094 11648
rect 25314 11636 25320 11688
rect 25372 11636 25378 11688
rect 26050 11636 26056 11688
rect 26108 11636 26114 11688
rect 27908 11676 27936 11704
rect 28460 11676 28488 11716
rect 28629 11713 28641 11716
rect 28675 11713 28687 11747
rect 28629 11707 28687 11713
rect 27908 11648 28488 11676
rect 24857 11611 24915 11617
rect 22066 11580 22508 11608
rect 22480 11552 22508 11580
rect 24857 11577 24869 11611
rect 24903 11608 24915 11611
rect 27908 11608 27936 11648
rect 28534 11636 28540 11688
rect 28592 11636 28598 11688
rect 24903 11580 27936 11608
rect 24903 11577 24915 11580
rect 24857 11571 24915 11577
rect 28074 11568 28080 11620
rect 28132 11608 28138 11620
rect 28261 11611 28319 11617
rect 28261 11608 28273 11611
rect 28132 11580 28273 11608
rect 28132 11568 28138 11580
rect 28261 11577 28273 11580
rect 28307 11577 28319 11611
rect 28261 11571 28319 11577
rect 14182 11540 14188 11552
rect 13924 11512 14188 11540
rect 14182 11500 14188 11512
rect 14240 11500 14246 11552
rect 14826 11500 14832 11552
rect 14884 11540 14890 11552
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14884 11512 15117 11540
rect 14884 11500 14890 11512
rect 15105 11509 15117 11512
rect 15151 11540 15163 11543
rect 15194 11540 15200 11552
rect 15151 11512 15200 11540
rect 15151 11509 15163 11512
rect 15105 11503 15163 11509
rect 15194 11500 15200 11512
rect 15252 11500 15258 11552
rect 16850 11500 16856 11552
rect 16908 11500 16914 11552
rect 19337 11543 19395 11549
rect 19337 11509 19349 11543
rect 19383 11540 19395 11543
rect 19518 11540 19524 11552
rect 19383 11512 19524 11540
rect 19383 11509 19395 11512
rect 19337 11503 19395 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 19610 11500 19616 11552
rect 19668 11500 19674 11552
rect 19705 11543 19763 11549
rect 19705 11509 19717 11543
rect 19751 11540 19763 11543
rect 20070 11540 20076 11552
rect 19751 11512 20076 11540
rect 19751 11509 19763 11512
rect 19705 11503 19763 11509
rect 20070 11500 20076 11512
rect 20128 11500 20134 11552
rect 20806 11500 20812 11552
rect 20864 11500 20870 11552
rect 22462 11500 22468 11552
rect 22520 11500 22526 11552
rect 23385 11543 23443 11549
rect 23385 11509 23397 11543
rect 23431 11540 23443 11543
rect 23750 11540 23756 11552
rect 23431 11512 23756 11540
rect 23431 11509 23443 11512
rect 23385 11503 23443 11509
rect 23750 11500 23756 11512
rect 23808 11500 23814 11552
rect 27617 11543 27675 11549
rect 27617 11509 27629 11543
rect 27663 11540 27675 11543
rect 27798 11540 27804 11552
rect 27663 11512 27804 11540
rect 27663 11509 27675 11512
rect 27617 11503 27675 11509
rect 27798 11500 27804 11512
rect 27856 11500 27862 11552
rect 1104 11450 35248 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 35248 11450
rect 1104 11376 35248 11398
rect 9122 11296 9128 11348
rect 9180 11296 9186 11348
rect 11054 11296 11060 11348
rect 11112 11336 11118 11348
rect 11241 11339 11299 11345
rect 11241 11336 11253 11339
rect 11112 11308 11253 11336
rect 11112 11296 11118 11308
rect 11241 11305 11253 11308
rect 11287 11305 11299 11339
rect 11241 11299 11299 11305
rect 11698 11296 11704 11348
rect 11756 11296 11762 11348
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12158 11336 12164 11348
rect 12115 11308 12164 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12158 11296 12164 11308
rect 12216 11296 12222 11348
rect 14921 11339 14979 11345
rect 14921 11336 14933 11339
rect 12268 11308 14933 11336
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 12268 11268 12296 11308
rect 14921 11305 14933 11308
rect 14967 11336 14979 11339
rect 15010 11336 15016 11348
rect 14967 11308 15016 11336
rect 14967 11305 14979 11308
rect 14921 11299 14979 11305
rect 15010 11296 15016 11308
rect 15068 11336 15074 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15068 11308 15485 11336
rect 15068 11296 15074 11308
rect 15473 11305 15485 11308
rect 15519 11305 15531 11339
rect 15473 11299 15531 11305
rect 16390 11296 16396 11348
rect 16448 11296 16454 11348
rect 19426 11296 19432 11348
rect 19484 11296 19490 11348
rect 19610 11296 19616 11348
rect 19668 11296 19674 11348
rect 24854 11296 24860 11348
rect 24912 11296 24918 11348
rect 25130 11296 25136 11348
rect 25188 11336 25194 11348
rect 25188 11308 25268 11336
rect 25188 11296 25194 11308
rect 11572 11240 12296 11268
rect 11572 11228 11578 11240
rect 9677 11203 9735 11209
rect 9677 11169 9689 11203
rect 9723 11200 9735 11203
rect 9723 11172 11192 11200
rect 9723 11169 9735 11172
rect 9677 11163 9735 11169
rect 9306 11092 9312 11144
rect 9364 11092 9370 11144
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9416 11008 9444 11095
rect 9766 11092 9772 11144
rect 9824 11092 9830 11144
rect 10045 11135 10103 11141
rect 10045 11101 10057 11135
rect 10091 11101 10103 11135
rect 10045 11095 10103 11101
rect 10060 11064 10088 11095
rect 10226 11092 10232 11144
rect 10284 11092 10290 11144
rect 11164 11141 11192 11172
rect 11606 11160 11612 11212
rect 11664 11200 11670 11212
rect 12066 11200 12072 11212
rect 11664 11172 12072 11200
rect 11664 11160 11670 11172
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 12268 11209 12296 11240
rect 14844 11240 15884 11268
rect 12253 11203 12311 11209
rect 12253 11169 12265 11203
rect 12299 11169 12311 11203
rect 12253 11163 12311 11169
rect 12710 11160 12716 11212
rect 12768 11200 12774 11212
rect 14642 11200 14648 11212
rect 12768 11172 14648 11200
rect 12768 11160 12774 11172
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 14844 11144 14872 11240
rect 15381 11203 15439 11209
rect 15381 11169 15393 11203
rect 15427 11200 15439 11203
rect 15470 11200 15476 11212
rect 15427 11172 15476 11200
rect 15427 11169 15439 11172
rect 15381 11163 15439 11169
rect 15470 11160 15476 11172
rect 15528 11160 15534 11212
rect 15562 11160 15568 11212
rect 15620 11160 15626 11212
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11101 11207 11135
rect 11149 11095 11207 11101
rect 10318 11064 10324 11076
rect 10060 11036 10324 11064
rect 10318 11024 10324 11036
rect 10376 11024 10382 11076
rect 11054 11024 11060 11076
rect 11112 11024 11118 11076
rect 11164 11064 11192 11095
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 13354 11092 13360 11144
rect 13412 11132 13418 11144
rect 13412 11104 14780 11132
rect 13412 11092 13418 11104
rect 12621 11067 12679 11073
rect 12621 11064 12633 11067
rect 11164 11036 12633 11064
rect 12621 11033 12633 11036
rect 12667 11064 12679 11067
rect 14752 11064 14780 11104
rect 14826 11092 14832 11144
rect 14884 11092 14890 11144
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11101 15163 11135
rect 15105 11095 15163 11101
rect 15120 11064 15148 11095
rect 15194 11092 15200 11144
rect 15252 11092 15258 11144
rect 15749 11135 15807 11141
rect 15749 11132 15761 11135
rect 15304 11104 15761 11132
rect 12667 11036 13860 11064
rect 14752 11036 15148 11064
rect 12667 11033 12679 11036
rect 12621 11027 12679 11033
rect 9398 10956 9404 11008
rect 9456 10956 9462 11008
rect 13832 10996 13860 11036
rect 14826 10996 14832 11008
rect 13832 10968 14832 10996
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 15120 10996 15148 11036
rect 15304 10996 15332 11104
rect 15749 11101 15761 11104
rect 15795 11101 15807 11135
rect 15856 11132 15884 11240
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 19444 11200 19472 11296
rect 19518 11228 19524 11280
rect 19576 11268 19582 11280
rect 20438 11268 20444 11280
rect 19576 11240 20444 11268
rect 19576 11228 19582 11240
rect 20438 11228 20444 11240
rect 20496 11228 20502 11280
rect 24872 11209 24900 11296
rect 25240 11277 25268 11308
rect 25314 11296 25320 11348
rect 25372 11296 25378 11348
rect 25501 11339 25559 11345
rect 25501 11305 25513 11339
rect 25547 11336 25559 11339
rect 26142 11336 26148 11348
rect 25547 11308 26148 11336
rect 25547 11305 25559 11308
rect 25501 11299 25559 11305
rect 26142 11296 26148 11308
rect 26200 11296 26206 11348
rect 27430 11296 27436 11348
rect 27488 11296 27494 11348
rect 27706 11296 27712 11348
rect 27764 11296 27770 11348
rect 25225 11271 25283 11277
rect 25225 11237 25237 11271
rect 25271 11237 25283 11271
rect 25225 11231 25283 11237
rect 24857 11203 24915 11209
rect 16172 11172 16528 11200
rect 19444 11172 19748 11200
rect 16172 11160 16178 11172
rect 16298 11132 16304 11144
rect 15856 11104 16304 11132
rect 15749 11095 15807 11101
rect 16298 11092 16304 11104
rect 16356 11132 16362 11144
rect 16500 11141 16528 11172
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 16356 11104 16405 11132
rect 16356 11092 16362 11104
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 18506 11132 18512 11144
rect 16531 11104 18512 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 18506 11092 18512 11104
rect 18564 11092 18570 11144
rect 19518 11092 19524 11144
rect 19576 11092 19582 11144
rect 19720 11141 19748 11172
rect 24857 11169 24869 11203
rect 24903 11169 24915 11203
rect 24857 11163 24915 11169
rect 27617 11203 27675 11209
rect 27617 11169 27629 11203
rect 27663 11200 27675 11203
rect 27724 11200 27752 11296
rect 27663 11172 27752 11200
rect 27663 11169 27675 11172
rect 27617 11163 27675 11169
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11101 19763 11135
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 19705 11095 19763 11101
rect 25332 11104 25421 11132
rect 25332 11076 25360 11104
rect 25409 11101 25421 11104
rect 25455 11132 25467 11135
rect 25498 11132 25504 11144
rect 25455 11104 25504 11132
rect 25455 11101 25467 11104
rect 25409 11095 25467 11101
rect 25498 11092 25504 11104
rect 25556 11092 25562 11144
rect 25590 11092 25596 11144
rect 25648 11092 25654 11144
rect 27709 11135 27767 11141
rect 27709 11101 27721 11135
rect 27755 11132 27767 11135
rect 28353 11135 28411 11141
rect 28353 11132 28365 11135
rect 27755 11104 28365 11132
rect 27755 11101 27767 11104
rect 27709 11095 27767 11101
rect 28353 11101 28365 11104
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 15473 11067 15531 11073
rect 15473 11033 15485 11067
rect 15519 11033 15531 11067
rect 15473 11027 15531 11033
rect 15120 10968 15332 10996
rect 15488 10996 15516 11027
rect 16666 11024 16672 11076
rect 16724 11024 16730 11076
rect 25314 11024 25320 11076
rect 25372 11024 25378 11076
rect 25608 11064 25636 11092
rect 25516 11036 25636 11064
rect 25516 11008 25544 11036
rect 27982 11024 27988 11076
rect 28040 11024 28046 11076
rect 28166 11024 28172 11076
rect 28224 11024 28230 11076
rect 15746 10996 15752 11008
rect 15488 10968 15752 10996
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 15933 10999 15991 11005
rect 15933 10965 15945 10999
rect 15979 10996 15991 10999
rect 16022 10996 16028 11008
rect 15979 10968 16028 10996
rect 15979 10965 15991 10968
rect 15933 10959 15991 10965
rect 16022 10956 16028 10968
rect 16080 10956 16086 11008
rect 16206 10956 16212 11008
rect 16264 10956 16270 11008
rect 25498 10956 25504 11008
rect 25556 10956 25562 11008
rect 1104 10906 35236 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 35236 10906
rect 1104 10832 35236 10854
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 13722 10792 13728 10804
rect 12759 10764 13728 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 13722 10752 13728 10764
rect 13780 10752 13786 10804
rect 16206 10752 16212 10804
rect 16264 10752 16270 10804
rect 21634 10752 21640 10804
rect 21692 10752 21698 10804
rect 21818 10752 21824 10804
rect 21876 10752 21882 10804
rect 23290 10752 23296 10804
rect 23348 10752 23354 10804
rect 24765 10795 24823 10801
rect 24765 10761 24777 10795
rect 24811 10792 24823 10795
rect 25314 10792 25320 10804
rect 24811 10764 25320 10792
rect 24811 10761 24823 10764
rect 24765 10755 24823 10761
rect 25314 10752 25320 10764
rect 25372 10752 25378 10804
rect 14372 10736 14424 10742
rect 11238 10724 11244 10736
rect 10350 10696 11244 10724
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 15013 10727 15071 10733
rect 15013 10724 15025 10727
rect 14372 10678 14424 10684
rect 14476 10696 15025 10724
rect 10410 10616 10416 10668
rect 10468 10616 10474 10668
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10873 10659 10931 10665
rect 10873 10656 10885 10659
rect 10836 10628 10885 10656
rect 10836 10616 10842 10628
rect 10873 10625 10885 10628
rect 10919 10625 10931 10659
rect 10873 10619 10931 10625
rect 12345 10659 12403 10665
rect 12345 10625 12357 10659
rect 12391 10656 12403 10659
rect 12986 10656 12992 10668
rect 12391 10628 12992 10656
rect 12391 10625 12403 10628
rect 12345 10619 12403 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13725 10659 13783 10665
rect 13725 10656 13737 10659
rect 13096 10628 13737 10656
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 13096 10588 13124 10628
rect 13725 10625 13737 10628
rect 13771 10646 13783 10659
rect 13998 10656 14004 10668
rect 13924 10646 14004 10656
rect 13771 10628 14004 10646
rect 13771 10625 13952 10628
rect 13725 10619 13952 10625
rect 13740 10618 13952 10619
rect 13998 10616 14004 10628
rect 14056 10616 14062 10668
rect 12483 10560 13124 10588
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 13446 10480 13452 10532
rect 13504 10520 13510 10532
rect 13906 10520 13912 10532
rect 13504 10492 13912 10520
rect 13504 10480 13510 10492
rect 13906 10480 13912 10492
rect 13964 10520 13970 10532
rect 14476 10520 14504 10696
rect 15013 10693 15025 10696
rect 15059 10693 15071 10727
rect 15013 10687 15071 10693
rect 16022 10684 16028 10736
rect 16080 10684 16086 10736
rect 16117 10727 16175 10733
rect 16117 10693 16129 10727
rect 16163 10724 16175 10727
rect 16224 10724 16252 10752
rect 23308 10724 23336 10752
rect 16163 10696 17264 10724
rect 16163 10693 16175 10696
rect 16117 10687 16175 10693
rect 14826 10616 14832 10668
rect 14884 10616 14890 10668
rect 17236 10665 17264 10696
rect 21192 10696 22416 10724
rect 23308 10696 23520 10724
rect 15105 10659 15163 10665
rect 15105 10656 15117 10659
rect 14936 10628 15117 10656
rect 13964 10492 14504 10520
rect 13964 10480 13970 10492
rect 9309 10455 9367 10461
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9398 10452 9404 10464
rect 9355 10424 9404 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9398 10412 9404 10424
rect 9456 10452 9462 10464
rect 11330 10452 11336 10464
rect 9456 10424 11336 10452
rect 9456 10412 9462 10424
rect 11330 10412 11336 10424
rect 11388 10412 11394 10464
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 14936 10452 14964 10628
rect 15105 10625 15117 10628
rect 15151 10625 15163 10659
rect 15105 10619 15163 10625
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10625 15255 10659
rect 15841 10659 15899 10665
rect 15841 10656 15853 10659
rect 15197 10619 15255 10625
rect 15672 10628 15853 10656
rect 15212 10588 15240 10619
rect 15378 10588 15384 10600
rect 15212 10560 15384 10588
rect 15378 10548 15384 10560
rect 15436 10548 15442 10600
rect 15672 10532 15700 10628
rect 15841 10625 15853 10628
rect 15887 10625 15899 10659
rect 16209 10659 16267 10665
rect 16209 10656 16221 10659
rect 15841 10619 15899 10625
rect 16132 10628 16221 10656
rect 15654 10520 15660 10532
rect 15396 10492 15660 10520
rect 15396 10461 15424 10492
rect 15654 10480 15660 10492
rect 15712 10480 15718 10532
rect 16132 10464 16160 10628
rect 16209 10625 16221 10628
rect 16255 10625 16267 10659
rect 16209 10619 16267 10625
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10625 17279 10659
rect 17221 10619 17279 10625
rect 17310 10548 17316 10600
rect 17368 10548 17374 10600
rect 21192 10597 21220 10696
rect 21358 10616 21364 10668
rect 21416 10616 21422 10668
rect 21450 10616 21456 10668
rect 21508 10656 21514 10668
rect 22005 10659 22063 10665
rect 22005 10656 22017 10659
rect 21508 10628 22017 10656
rect 21508 10616 21514 10628
rect 22005 10625 22017 10628
rect 22051 10625 22063 10659
rect 22005 10619 22063 10625
rect 22094 10616 22100 10668
rect 22152 10616 22158 10668
rect 22388 10665 22416 10696
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 21177 10591 21235 10597
rect 21177 10557 21189 10591
rect 21223 10557 21235 10591
rect 21177 10551 21235 10557
rect 21269 10591 21327 10597
rect 21269 10557 21281 10591
rect 21315 10588 21327 10591
rect 21910 10588 21916 10600
rect 21315 10560 21916 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 17589 10523 17647 10529
rect 17589 10489 17601 10523
rect 17635 10520 17647 10523
rect 17678 10520 17684 10532
rect 17635 10492 17684 10520
rect 17635 10489 17647 10492
rect 17589 10483 17647 10489
rect 17678 10480 17684 10492
rect 17736 10480 17742 10532
rect 21192 10520 21220 10551
rect 21910 10548 21916 10560
rect 21968 10588 21974 10600
rect 22204 10588 22232 10619
rect 22462 10616 22468 10668
rect 22520 10616 22526 10668
rect 22922 10616 22928 10668
rect 22980 10656 22986 10668
rect 23293 10659 23351 10665
rect 23293 10656 23305 10659
rect 22980 10628 23305 10656
rect 22980 10616 22986 10628
rect 23293 10625 23305 10628
rect 23339 10625 23351 10659
rect 23293 10619 23351 10625
rect 23492 10597 23520 10696
rect 23591 10659 23649 10665
rect 23591 10625 23603 10659
rect 23637 10656 23649 10659
rect 24581 10659 24639 10665
rect 24581 10656 24593 10659
rect 23637 10628 24593 10656
rect 23637 10625 23649 10628
rect 23591 10619 23649 10625
rect 24581 10625 24593 10628
rect 24627 10625 24639 10659
rect 24581 10619 24639 10625
rect 26418 10616 26424 10668
rect 26476 10656 26482 10668
rect 26513 10659 26571 10665
rect 26513 10656 26525 10659
rect 26476 10628 26525 10656
rect 26476 10616 26482 10628
rect 26513 10625 26525 10628
rect 26559 10625 26571 10659
rect 26513 10619 26571 10625
rect 26697 10659 26755 10665
rect 26697 10625 26709 10659
rect 26743 10656 26755 10659
rect 26786 10656 26792 10668
rect 26743 10628 26792 10656
rect 26743 10625 26755 10628
rect 26697 10619 26755 10625
rect 26786 10616 26792 10628
rect 26844 10616 26850 10668
rect 21968 10560 22232 10588
rect 23477 10591 23535 10597
rect 21968 10548 21974 10560
rect 23477 10557 23489 10591
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 23842 10548 23848 10600
rect 23900 10588 23906 10600
rect 24397 10591 24455 10597
rect 24397 10588 24409 10591
rect 23900 10560 24409 10588
rect 23900 10548 23906 10560
rect 24397 10557 24409 10560
rect 24443 10588 24455 10591
rect 24670 10588 24676 10600
rect 24443 10560 24676 10588
rect 24443 10557 24455 10560
rect 24397 10551 24455 10557
rect 24670 10548 24676 10560
rect 24728 10548 24734 10600
rect 23661 10523 23719 10529
rect 21192 10492 21312 10520
rect 21284 10464 21312 10492
rect 23661 10489 23673 10523
rect 23707 10520 23719 10523
rect 23934 10520 23940 10532
rect 23707 10492 23940 10520
rect 23707 10489 23719 10492
rect 23661 10483 23719 10489
rect 23934 10480 23940 10492
rect 23992 10480 23998 10532
rect 24026 10480 24032 10532
rect 24084 10480 24090 10532
rect 12216 10424 14964 10452
rect 15381 10455 15439 10461
rect 12216 10412 12222 10424
rect 15381 10421 15393 10455
rect 15427 10421 15439 10455
rect 15381 10415 15439 10421
rect 16114 10412 16120 10464
rect 16172 10412 16178 10464
rect 16390 10412 16396 10464
rect 16448 10412 16454 10464
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 19886 10452 19892 10464
rect 17828 10424 19892 10452
rect 17828 10412 17834 10424
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 23385 10455 23443 10461
rect 23385 10421 23397 10455
rect 23431 10452 23443 10455
rect 23566 10452 23572 10464
rect 23431 10424 23572 10452
rect 23431 10421 23443 10424
rect 23385 10415 23443 10421
rect 23566 10412 23572 10424
rect 23624 10452 23630 10464
rect 24044 10452 24072 10480
rect 23624 10424 24072 10452
rect 23624 10412 23630 10424
rect 26510 10412 26516 10464
rect 26568 10412 26574 10464
rect 1104 10362 35248 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 35248 10362
rect 1104 10288 35248 10310
rect 10870 10208 10876 10260
rect 10928 10208 10934 10260
rect 14550 10248 14556 10260
rect 13648 10220 14556 10248
rect 13648 10180 13676 10220
rect 14550 10208 14556 10220
rect 14608 10248 14614 10260
rect 15378 10248 15384 10260
rect 14608 10220 15384 10248
rect 14608 10208 14614 10220
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 16022 10208 16028 10260
rect 16080 10248 16086 10260
rect 17310 10248 17316 10260
rect 16080 10220 17316 10248
rect 16080 10208 16086 10220
rect 17310 10208 17316 10220
rect 17368 10248 17374 10260
rect 17589 10251 17647 10257
rect 17589 10248 17601 10251
rect 17368 10220 17601 10248
rect 17368 10208 17374 10220
rect 17589 10217 17601 10220
rect 17635 10217 17647 10251
rect 17589 10211 17647 10217
rect 18322 10208 18328 10260
rect 18380 10208 18386 10260
rect 20809 10251 20867 10257
rect 20809 10217 20821 10251
rect 20855 10248 20867 10251
rect 21266 10248 21272 10260
rect 20855 10220 21272 10248
rect 20855 10217 20867 10220
rect 20809 10211 20867 10217
rect 21266 10208 21272 10220
rect 21324 10248 21330 10260
rect 22465 10251 22523 10257
rect 22465 10248 22477 10251
rect 21324 10220 22477 10248
rect 21324 10208 21330 10220
rect 12728 10152 13676 10180
rect 12728 10121 12756 10152
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10081 12771 10115
rect 13538 10112 13544 10124
rect 12713 10075 12771 10081
rect 13372 10084 13544 10112
rect 7285 10047 7343 10053
rect 7285 10013 7297 10047
rect 7331 10044 7343 10047
rect 7331 10016 7604 10044
rect 7331 10013 7343 10016
rect 7285 10007 7343 10013
rect 7576 9908 7604 10016
rect 7742 10004 7748 10056
rect 7800 10044 7806 10056
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 7800 10016 9045 10044
rect 7800 10004 7806 10016
rect 9033 10013 9045 10016
rect 9079 10013 9091 10047
rect 9033 10007 9091 10013
rect 9398 10004 9404 10056
rect 9456 10004 9462 10056
rect 11054 10004 11060 10056
rect 11112 10004 11118 10056
rect 11698 10004 11704 10056
rect 11756 10004 11762 10056
rect 11882 10004 11888 10056
rect 11940 10004 11946 10056
rect 12434 10004 12440 10056
rect 12492 10044 12498 10056
rect 13372 10053 13400 10084
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13648 10053 13676 10152
rect 13722 10140 13728 10192
rect 13780 10140 13786 10192
rect 13909 10183 13967 10189
rect 13909 10149 13921 10183
rect 13955 10180 13967 10183
rect 18141 10183 18199 10189
rect 13955 10152 18092 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 13740 10112 13768 10140
rect 14274 10112 14280 10124
rect 13740 10084 14280 10112
rect 14274 10072 14280 10084
rect 14332 10112 14338 10124
rect 14332 10084 14504 10112
rect 14332 10072 14338 10084
rect 13357 10047 13415 10053
rect 13357 10044 13369 10047
rect 12492 10016 13369 10044
rect 12492 10004 12498 10016
rect 13357 10013 13369 10016
rect 13403 10013 13415 10047
rect 13357 10007 13415 10013
rect 13633 10047 13691 10053
rect 13633 10013 13645 10047
rect 13679 10013 13691 10047
rect 13633 10007 13691 10013
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14182 10044 14188 10056
rect 14139 10016 14188 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 11072 9976 11100 10004
rect 13446 9976 13452 9988
rect 8418 9948 9674 9976
rect 11072 9948 13452 9976
rect 9398 9908 9404 9920
rect 7576 9880 9404 9908
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9646 9908 9674 9948
rect 13446 9936 13452 9948
rect 13504 9976 13510 9988
rect 13541 9979 13599 9985
rect 13541 9976 13553 9979
rect 13504 9948 13553 9976
rect 13504 9936 13510 9948
rect 13541 9945 13553 9948
rect 13587 9945 13599 9979
rect 13541 9939 13599 9945
rect 13740 9976 13768 10007
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14476 10053 14504 10084
rect 15654 10072 15660 10124
rect 15712 10112 15718 10124
rect 17497 10115 17555 10121
rect 17497 10112 17509 10115
rect 15712 10084 15792 10112
rect 15712 10072 15718 10084
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10013 14519 10047
rect 14918 10044 14924 10056
rect 14461 10007 14519 10013
rect 14568 10016 14924 10044
rect 14277 9979 14335 9985
rect 14277 9976 14289 9979
rect 13740 9948 14289 9976
rect 11790 9908 11796 9920
rect 9646 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9908 11854 9920
rect 13740 9908 13768 9948
rect 14277 9945 14289 9948
rect 14323 9945 14335 9979
rect 14277 9939 14335 9945
rect 14366 9936 14372 9988
rect 14424 9976 14430 9988
rect 14568 9976 14596 10016
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15764 10053 15792 10084
rect 16224 10084 17509 10112
rect 16224 10056 16252 10084
rect 15749 10047 15807 10053
rect 15749 10013 15761 10047
rect 15795 10013 15807 10047
rect 15749 10007 15807 10013
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16022 10044 16028 10056
rect 15979 10016 16028 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16022 10004 16028 10016
rect 16080 10004 16086 10056
rect 16114 10004 16120 10056
rect 16172 10004 16178 10056
rect 16206 10004 16212 10056
rect 16264 10004 16270 10056
rect 16298 10004 16304 10056
rect 16356 10004 16362 10056
rect 16500 10053 16528 10084
rect 17497 10081 17509 10084
rect 17543 10081 17555 10115
rect 18064 10112 18092 10152
rect 18141 10149 18153 10183
rect 18187 10180 18199 10183
rect 19334 10180 19340 10192
rect 18187 10152 19340 10180
rect 18187 10149 18199 10152
rect 18141 10143 18199 10149
rect 19334 10140 19340 10152
rect 19392 10140 19398 10192
rect 20165 10183 20223 10189
rect 20165 10149 20177 10183
rect 20211 10180 20223 10183
rect 21450 10180 21456 10192
rect 20211 10152 21456 10180
rect 20211 10149 20223 10152
rect 20165 10143 20223 10149
rect 21450 10140 21456 10152
rect 21508 10140 21514 10192
rect 18064 10084 18184 10112
rect 17497 10075 17555 10081
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10013 16543 10047
rect 16485 10007 16543 10013
rect 17770 10004 17776 10056
rect 17828 10044 17834 10056
rect 17960 10047 18018 10053
rect 17960 10044 17972 10047
rect 17828 10016 17972 10044
rect 17828 10004 17834 10016
rect 17960 10013 17972 10016
rect 18006 10013 18018 10047
rect 18156 10044 18184 10084
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 18288 10084 18337 10112
rect 18288 10072 18294 10084
rect 18325 10081 18337 10084
rect 18371 10081 18383 10115
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 18325 10075 18383 10081
rect 18432 10084 18828 10112
rect 18432 10044 18460 10084
rect 18156 10016 18460 10044
rect 17960 10007 18018 10013
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 18800 10053 18828 10084
rect 18984 10084 19809 10112
rect 18984 10053 19012 10084
rect 19797 10081 19809 10084
rect 19843 10112 19855 10115
rect 20257 10115 20315 10121
rect 20257 10112 20269 10115
rect 19843 10084 20269 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 20257 10081 20269 10084
rect 20303 10081 20315 10115
rect 20257 10075 20315 10081
rect 18785 10047 18843 10053
rect 18785 10013 18797 10047
rect 18831 10013 18843 10047
rect 18785 10007 18843 10013
rect 18969 10047 19027 10053
rect 18969 10013 18981 10047
rect 19015 10013 19027 10047
rect 18969 10007 19027 10013
rect 19705 10047 19763 10053
rect 19705 10013 19717 10047
rect 19751 10013 19763 10047
rect 19705 10007 19763 10013
rect 16132 9976 16160 10004
rect 14424 9948 14596 9976
rect 14660 9948 16160 9976
rect 14424 9936 14430 9948
rect 14660 9917 14688 9948
rect 18046 9936 18052 9988
rect 18104 9976 18110 9988
rect 18233 9979 18291 9985
rect 18233 9976 18245 9979
rect 18104 9948 18245 9976
rect 18104 9936 18110 9948
rect 18233 9945 18245 9948
rect 18279 9945 18291 9979
rect 18984 9976 19012 10007
rect 18233 9939 18291 9945
rect 18708 9948 19012 9976
rect 19720 9976 19748 10007
rect 19886 10004 19892 10056
rect 19944 10004 19950 10056
rect 19981 10047 20039 10053
rect 19981 10013 19993 10047
rect 20027 10044 20039 10047
rect 20530 10044 20536 10056
rect 20027 10016 20536 10044
rect 20027 10013 20039 10016
rect 19981 10007 20039 10013
rect 20530 10004 20536 10016
rect 20588 10004 20594 10056
rect 21468 10053 21496 10140
rect 21744 10053 21772 10220
rect 22465 10217 22477 10220
rect 22511 10217 22523 10251
rect 22465 10211 22523 10217
rect 22922 10208 22928 10260
rect 22980 10248 22986 10260
rect 23385 10251 23443 10257
rect 23385 10248 23397 10251
rect 22980 10220 23397 10248
rect 22980 10208 22986 10220
rect 23385 10217 23397 10220
rect 23431 10217 23443 10251
rect 23385 10211 23443 10217
rect 23842 10208 23848 10260
rect 23900 10208 23906 10260
rect 24118 10208 24124 10260
rect 24176 10208 24182 10260
rect 24765 10251 24823 10257
rect 24765 10217 24777 10251
rect 24811 10248 24823 10251
rect 25498 10248 25504 10260
rect 24811 10220 25504 10248
rect 24811 10217 24823 10220
rect 24765 10211 24823 10217
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 22094 10140 22100 10192
rect 22152 10180 22158 10192
rect 22152 10152 22784 10180
rect 22152 10140 22158 10152
rect 22756 10121 22784 10152
rect 23290 10140 23296 10192
rect 23348 10180 23354 10192
rect 23348 10152 23704 10180
rect 23348 10140 23354 10152
rect 22649 10115 22707 10121
rect 22649 10112 22661 10115
rect 21954 10084 22661 10112
rect 21954 10056 21982 10084
rect 22649 10081 22661 10084
rect 22695 10081 22707 10115
rect 22649 10075 22707 10081
rect 22741 10115 22799 10121
rect 22741 10081 22753 10115
rect 22787 10081 22799 10115
rect 22741 10075 22799 10081
rect 23566 10072 23572 10124
rect 23624 10072 23630 10124
rect 21453 10047 21511 10053
rect 21453 10013 21465 10047
rect 21499 10013 21511 10047
rect 21453 10007 21511 10013
rect 21729 10047 21787 10053
rect 21729 10013 21741 10047
rect 21775 10013 21787 10047
rect 21729 10007 21787 10013
rect 21821 10047 21879 10053
rect 21821 10013 21833 10047
rect 21867 10013 21879 10047
rect 21821 10007 21879 10013
rect 20254 9976 20260 9988
rect 19720 9948 20260 9976
rect 11848 9880 13768 9908
rect 14645 9911 14703 9917
rect 11848 9868 11854 9880
rect 14645 9877 14657 9911
rect 14691 9877 14703 9911
rect 14645 9871 14703 9877
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 18708 9917 18736 9948
rect 20254 9936 20260 9948
rect 20312 9976 20318 9988
rect 20625 9979 20683 9985
rect 20625 9976 20637 9979
rect 20312 9948 20637 9976
rect 20312 9936 20318 9948
rect 20625 9945 20637 9948
rect 20671 9945 20683 9979
rect 20625 9939 20683 9945
rect 21545 9979 21603 9985
rect 21545 9945 21557 9979
rect 21591 9976 21603 9979
rect 21836 9976 21864 10007
rect 21910 10004 21916 10056
rect 21968 10053 21982 10056
rect 21968 10047 21990 10053
rect 21978 10013 21990 10047
rect 21968 10007 21990 10013
rect 21968 10004 21974 10007
rect 22094 10004 22100 10056
rect 22152 10044 22158 10056
rect 23676 10053 23704 10152
rect 26786 10072 26792 10124
rect 26844 10072 26850 10124
rect 22373 10047 22431 10053
rect 22152 10016 22194 10044
rect 22152 10004 22158 10016
rect 22373 10013 22385 10047
rect 22419 10013 22431 10047
rect 22373 10007 22431 10013
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 22388 9976 22416 10007
rect 23934 10004 23940 10056
rect 23992 10004 23998 10056
rect 24486 10004 24492 10056
rect 24544 10004 24550 10056
rect 24578 10004 24584 10056
rect 24636 10004 24642 10056
rect 24854 10004 24860 10056
rect 24912 10004 24918 10056
rect 24946 10004 24952 10056
rect 25004 10004 25010 10056
rect 25133 10047 25191 10053
rect 25133 10013 25145 10047
rect 25179 10013 25191 10047
rect 25133 10007 25191 10013
rect 21591 9948 22416 9976
rect 21591 9945 21603 9948
rect 21545 9939 21603 9945
rect 23290 9936 23296 9988
rect 23348 9976 23354 9988
rect 23385 9979 23443 9985
rect 23385 9976 23397 9979
rect 23348 9948 23397 9976
rect 23348 9936 23354 9948
rect 23385 9945 23397 9948
rect 23431 9976 23443 9979
rect 23952 9976 23980 10004
rect 23431 9948 23980 9976
rect 24872 9976 24900 10004
rect 25148 9976 25176 10007
rect 26418 10004 26424 10056
rect 26476 10044 26482 10056
rect 26973 10047 27031 10053
rect 26973 10044 26985 10047
rect 26476 10016 26985 10044
rect 26476 10004 26482 10016
rect 26973 10013 26985 10016
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 27157 10047 27215 10053
rect 27157 10013 27169 10047
rect 27203 10044 27215 10047
rect 27249 10047 27307 10053
rect 27249 10044 27261 10047
rect 27203 10016 27261 10044
rect 27203 10013 27215 10016
rect 27157 10007 27215 10013
rect 27249 10013 27261 10016
rect 27295 10013 27307 10047
rect 27249 10007 27307 10013
rect 27433 10047 27491 10053
rect 27433 10013 27445 10047
rect 27479 10013 27491 10047
rect 27433 10007 27491 10013
rect 24872 9948 25176 9976
rect 23431 9945 23443 9948
rect 23385 9939 23443 9945
rect 26510 9936 26516 9988
rect 26568 9976 26574 9988
rect 27448 9976 27476 10007
rect 26568 9948 27476 9976
rect 26568 9936 26574 9948
rect 17957 9911 18015 9917
rect 17957 9908 17969 9911
rect 17644 9880 17969 9908
rect 17644 9868 17650 9880
rect 17957 9877 17969 9880
rect 18003 9877 18015 9911
rect 17957 9871 18015 9877
rect 18693 9911 18751 9917
rect 18693 9877 18705 9911
rect 18739 9877 18751 9911
rect 18693 9871 18751 9877
rect 18874 9868 18880 9920
rect 18932 9868 18938 9920
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 20441 9911 20499 9917
rect 20441 9908 20453 9911
rect 19944 9880 20453 9908
rect 19944 9868 19950 9880
rect 20441 9877 20453 9880
rect 20487 9877 20499 9911
rect 20441 9871 20499 9877
rect 21358 9868 21364 9920
rect 21416 9908 21422 9920
rect 22094 9908 22100 9920
rect 21416 9880 22100 9908
rect 21416 9868 21422 9880
rect 22094 9868 22100 9880
rect 22152 9868 22158 9920
rect 22278 9868 22284 9920
rect 22336 9868 22342 9920
rect 22738 9868 22744 9920
rect 22796 9868 22802 9920
rect 25041 9911 25099 9917
rect 25041 9877 25053 9911
rect 25087 9908 25099 9911
rect 25498 9908 25504 9920
rect 25087 9880 25504 9908
rect 25087 9877 25099 9880
rect 25041 9871 25099 9877
rect 25498 9868 25504 9880
rect 25556 9868 25562 9920
rect 27338 9868 27344 9920
rect 27396 9868 27402 9920
rect 1104 9818 35236 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 35236 9818
rect 1104 9744 35236 9766
rect 10870 9664 10876 9716
rect 10928 9704 10934 9716
rect 15838 9704 15844 9716
rect 10928 9676 15844 9704
rect 10928 9664 10934 9676
rect 15838 9664 15844 9676
rect 15896 9664 15902 9716
rect 18322 9704 18328 9716
rect 17420 9676 18328 9704
rect 11698 9636 11704 9648
rect 9890 9608 10916 9636
rect 8754 9528 8760 9580
rect 8812 9528 8818 9580
rect 9214 9528 9220 9580
rect 9272 9528 9278 9580
rect 10888 9432 10916 9608
rect 10980 9608 11704 9636
rect 10980 9580 11008 9608
rect 11698 9596 11704 9608
rect 11756 9636 11762 9648
rect 13541 9639 13599 9645
rect 11756 9608 12112 9636
rect 11756 9596 11762 9608
rect 10962 9528 10968 9580
rect 11020 9528 11026 9580
rect 11882 9528 11888 9580
rect 11940 9528 11946 9580
rect 12084 9577 12112 9608
rect 13541 9605 13553 9639
rect 13587 9636 13599 9639
rect 15562 9636 15568 9648
rect 13587 9608 15568 9636
rect 13587 9605 13599 9608
rect 13541 9599 13599 9605
rect 15562 9596 15568 9608
rect 15620 9636 15626 9648
rect 17420 9636 17448 9676
rect 15620 9608 17448 9636
rect 17497 9639 17555 9645
rect 15620 9596 15626 9608
rect 17497 9605 17509 9639
rect 17543 9636 17555 9639
rect 17586 9636 17592 9648
rect 17543 9608 17592 9636
rect 17543 9605 17555 9608
rect 17497 9599 17555 9605
rect 17586 9596 17592 9608
rect 17644 9596 17650 9648
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 17773 9571 17831 9577
rect 17773 9568 17785 9571
rect 15436 9540 17785 9568
rect 15436 9528 15442 9540
rect 17773 9537 17785 9540
rect 17819 9537 17831 9571
rect 17773 9531 17831 9537
rect 17957 9571 18015 9577
rect 17957 9537 17969 9571
rect 18003 9537 18015 9571
rect 17957 9531 18015 9537
rect 18049 9571 18107 9577
rect 18049 9537 18061 9571
rect 18095 9568 18107 9571
rect 18156 9568 18184 9676
rect 18322 9664 18328 9676
rect 18380 9664 18386 9716
rect 20530 9664 20536 9716
rect 20588 9664 20594 9716
rect 21545 9707 21603 9713
rect 21545 9673 21557 9707
rect 21591 9704 21603 9707
rect 21910 9704 21916 9716
rect 21591 9676 21916 9704
rect 21591 9673 21603 9676
rect 21545 9667 21603 9673
rect 21910 9664 21916 9676
rect 21968 9664 21974 9716
rect 22278 9664 22284 9716
rect 22336 9664 22342 9716
rect 22738 9664 22744 9716
rect 22796 9664 22802 9716
rect 24029 9707 24087 9713
rect 23400 9676 23980 9704
rect 21174 9596 21180 9648
rect 21232 9596 21238 9648
rect 22296 9636 22324 9664
rect 22112 9608 22324 9636
rect 18095 9540 18184 9568
rect 18233 9571 18291 9577
rect 18095 9537 18107 9540
rect 18049 9531 18107 9537
rect 18233 9537 18245 9571
rect 18279 9568 18291 9571
rect 18506 9568 18512 9580
rect 18279 9540 18512 9568
rect 18279 9537 18291 9540
rect 18233 9531 18291 9537
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16666 9500 16672 9512
rect 15896 9472 16672 9500
rect 15896 9460 15902 9472
rect 16666 9460 16672 9472
rect 16724 9500 16730 9512
rect 17589 9503 17647 9509
rect 17589 9500 17601 9503
rect 16724 9472 17601 9500
rect 16724 9460 16730 9472
rect 17589 9469 17601 9472
rect 17635 9500 17647 9503
rect 17862 9500 17868 9512
rect 17635 9472 17868 9500
rect 17635 9469 17647 9472
rect 17589 9463 17647 9469
rect 17862 9460 17868 9472
rect 17920 9460 17926 9512
rect 17972 9500 18000 9531
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19705 9571 19763 9577
rect 19705 9568 19717 9571
rect 19392 9540 19717 9568
rect 19392 9528 19398 9540
rect 19705 9537 19717 9540
rect 19751 9568 19763 9571
rect 20165 9571 20223 9577
rect 20165 9568 20177 9571
rect 19751 9540 20177 9568
rect 19751 9537 19763 9540
rect 19705 9531 19763 9537
rect 20165 9537 20177 9540
rect 20211 9537 20223 9571
rect 20165 9531 20223 9537
rect 20349 9571 20407 9577
rect 20349 9537 20361 9571
rect 20395 9568 20407 9571
rect 20530 9568 20536 9580
rect 20395 9540 20536 9568
rect 20395 9537 20407 9540
rect 20349 9531 20407 9537
rect 20530 9528 20536 9540
rect 20588 9528 20594 9580
rect 22112 9577 22140 9608
rect 21361 9571 21419 9577
rect 21361 9537 21373 9571
rect 21407 9537 21419 9571
rect 21361 9531 21419 9537
rect 22097 9571 22155 9577
rect 22097 9537 22109 9571
rect 22143 9537 22155 9571
rect 22097 9531 22155 9537
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9568 22339 9571
rect 22756 9568 22784 9664
rect 23014 9596 23020 9648
rect 23072 9596 23078 9648
rect 22327 9540 22784 9568
rect 22327 9537 22339 9540
rect 22281 9531 22339 9537
rect 19797 9503 19855 9509
rect 17972 9472 18092 9500
rect 12434 9432 12440 9444
rect 10888 9404 12440 9432
rect 12434 9392 12440 9404
rect 12492 9392 12498 9444
rect 15746 9324 15752 9376
rect 15804 9364 15810 9376
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 15804 9336 17693 9364
rect 15804 9324 15810 9336
rect 17681 9333 17693 9336
rect 17727 9364 17739 9367
rect 17954 9364 17960 9376
rect 17727 9336 17960 9364
rect 17727 9333 17739 9336
rect 17681 9327 17739 9333
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 18064 9373 18092 9472
rect 19797 9469 19809 9503
rect 19843 9500 19855 9503
rect 19978 9500 19984 9512
rect 19843 9472 19984 9500
rect 19843 9469 19855 9472
rect 19797 9463 19855 9469
rect 19978 9460 19984 9472
rect 20036 9460 20042 9512
rect 20073 9503 20131 9509
rect 20073 9469 20085 9503
rect 20119 9500 20131 9503
rect 20990 9500 20996 9512
rect 20119 9472 20996 9500
rect 20119 9469 20131 9472
rect 20073 9463 20131 9469
rect 20990 9460 20996 9472
rect 21048 9500 21054 9512
rect 21376 9500 21404 9531
rect 21048 9472 21404 9500
rect 23032 9500 23060 9596
rect 23400 9509 23428 9676
rect 23952 9580 23980 9676
rect 24029 9673 24041 9707
rect 24075 9704 24087 9707
rect 24578 9704 24584 9716
rect 24075 9676 24584 9704
rect 24075 9673 24087 9676
rect 24029 9667 24087 9673
rect 24578 9664 24584 9676
rect 24636 9664 24642 9716
rect 24765 9707 24823 9713
rect 24765 9673 24777 9707
rect 24811 9673 24823 9707
rect 24765 9667 24823 9673
rect 24486 9596 24492 9648
rect 24544 9636 24550 9648
rect 24780 9636 24808 9667
rect 26053 9639 26111 9645
rect 26053 9636 26065 9639
rect 24544 9608 25084 9636
rect 24544 9596 24550 9608
rect 23753 9571 23811 9577
rect 23753 9537 23765 9571
rect 23799 9537 23811 9571
rect 23753 9531 23811 9537
rect 23385 9503 23443 9509
rect 23385 9500 23397 9503
rect 23032 9472 23397 9500
rect 21048 9460 21054 9472
rect 23385 9469 23397 9472
rect 23431 9469 23443 9503
rect 23385 9463 23443 9469
rect 23474 9460 23480 9512
rect 23532 9460 23538 9512
rect 23768 9500 23796 9531
rect 23842 9528 23848 9580
rect 23900 9528 23906 9580
rect 23934 9528 23940 9580
rect 23992 9568 23998 9580
rect 24121 9571 24179 9577
rect 24121 9568 24133 9571
rect 23992 9540 24133 9568
rect 23992 9528 23998 9540
rect 24121 9537 24133 9540
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 24210 9528 24216 9580
rect 24268 9568 24274 9580
rect 24581 9571 24639 9577
rect 24581 9568 24593 9571
rect 24268 9540 24593 9568
rect 24268 9528 24274 9540
rect 24581 9537 24593 9540
rect 24627 9537 24639 9571
rect 24581 9531 24639 9537
rect 24670 9528 24676 9580
rect 24728 9568 24734 9580
rect 25056 9577 25084 9608
rect 25424 9608 26065 9636
rect 25424 9577 25452 9608
rect 26053 9605 26065 9608
rect 26099 9636 26111 9639
rect 26510 9636 26516 9648
rect 26099 9608 26516 9636
rect 26099 9605 26111 9608
rect 26053 9599 26111 9605
rect 26510 9596 26516 9608
rect 26568 9596 26574 9648
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24728 9540 24869 9568
rect 24728 9528 24734 9540
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 24857 9531 24915 9537
rect 25041 9571 25099 9577
rect 25041 9537 25053 9571
rect 25087 9537 25099 9571
rect 25041 9531 25099 9537
rect 25409 9571 25467 9577
rect 25409 9537 25421 9571
rect 25455 9537 25467 9571
rect 25409 9531 25467 9537
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9568 25835 9571
rect 25823 9540 26004 9568
rect 25823 9537 25835 9540
rect 25777 9531 25835 9537
rect 24397 9503 24455 9509
rect 24397 9500 24409 9503
rect 23768 9472 24409 9500
rect 24136 9444 24164 9472
rect 24397 9469 24409 9472
rect 24443 9469 24455 9503
rect 24397 9463 24455 9469
rect 25498 9460 25504 9512
rect 25556 9500 25562 9512
rect 25685 9503 25743 9509
rect 25685 9500 25697 9503
rect 25556 9472 25697 9500
rect 25556 9460 25562 9472
rect 25685 9469 25697 9472
rect 25731 9500 25743 9503
rect 25869 9503 25927 9509
rect 25869 9500 25881 9503
rect 25731 9472 25881 9500
rect 25731 9469 25743 9472
rect 25685 9463 25743 9469
rect 25869 9469 25881 9472
rect 25915 9469 25927 9503
rect 25869 9463 25927 9469
rect 24118 9392 24124 9444
rect 24176 9392 24182 9444
rect 25406 9392 25412 9444
rect 25464 9432 25470 9444
rect 25593 9435 25651 9441
rect 25593 9432 25605 9435
rect 25464 9404 25605 9432
rect 25464 9392 25470 9404
rect 25593 9401 25605 9404
rect 25639 9432 25651 9435
rect 25976 9432 26004 9540
rect 26970 9528 26976 9580
rect 27028 9568 27034 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 27028 9540 27169 9568
rect 27028 9528 27034 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 27249 9503 27307 9509
rect 27249 9469 27261 9503
rect 27295 9500 27307 9503
rect 27338 9500 27344 9512
rect 27295 9472 27344 9500
rect 27295 9469 27307 9472
rect 27249 9463 27307 9469
rect 27338 9460 27344 9472
rect 27396 9460 27402 9512
rect 27522 9460 27528 9512
rect 27580 9460 27586 9512
rect 25639 9404 26004 9432
rect 25639 9401 25651 9404
rect 25593 9395 25651 9401
rect 18049 9367 18107 9373
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 19426 9364 19432 9376
rect 18095 9336 19432 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 19426 9324 19432 9336
rect 19484 9324 19490 9376
rect 22189 9367 22247 9373
rect 22189 9333 22201 9367
rect 22235 9364 22247 9367
rect 22462 9364 22468 9376
rect 22235 9336 22468 9364
rect 22235 9333 22247 9336
rect 22189 9327 22247 9333
rect 22462 9324 22468 9336
rect 22520 9324 22526 9376
rect 23382 9324 23388 9376
rect 23440 9364 23446 9376
rect 23842 9364 23848 9376
rect 23440 9336 23848 9364
rect 23440 9324 23446 9336
rect 23842 9324 23848 9336
rect 23900 9364 23906 9376
rect 24213 9367 24271 9373
rect 24213 9364 24225 9367
rect 23900 9336 24225 9364
rect 23900 9324 23906 9336
rect 24213 9333 24225 9336
rect 24259 9333 24271 9367
rect 24213 9327 24271 9333
rect 24854 9324 24860 9376
rect 24912 9364 24918 9376
rect 25041 9367 25099 9373
rect 25041 9364 25053 9367
rect 24912 9336 25053 9364
rect 24912 9324 24918 9336
rect 25041 9333 25053 9336
rect 25087 9333 25099 9367
rect 25041 9327 25099 9333
rect 25222 9324 25228 9376
rect 25280 9324 25286 9376
rect 25774 9324 25780 9376
rect 25832 9324 25838 9376
rect 1104 9274 35248 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 35248 9274
rect 1104 9200 35248 9222
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 14829 9163 14887 9169
rect 14829 9160 14841 9163
rect 11931 9132 14841 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 14829 9129 14841 9132
rect 14875 9160 14887 9163
rect 15746 9160 15752 9172
rect 14875 9132 15752 9160
rect 14875 9129 14887 9132
rect 14829 9123 14887 9129
rect 15746 9120 15752 9132
rect 15804 9120 15810 9172
rect 15838 9120 15844 9172
rect 15896 9120 15902 9172
rect 16577 9163 16635 9169
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 16623 9132 17356 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 14274 9052 14280 9104
rect 14332 9052 14338 9104
rect 14369 9095 14427 9101
rect 14369 9061 14381 9095
rect 14415 9092 14427 9095
rect 14734 9092 14740 9104
rect 14415 9064 14740 9092
rect 14415 9061 14427 9064
rect 14369 9055 14427 9061
rect 14734 9052 14740 9064
rect 14792 9052 14798 9104
rect 16209 9095 16267 9101
rect 16209 9061 16221 9095
rect 16255 9092 16267 9095
rect 16255 9064 16896 9092
rect 16255 9061 16267 9064
rect 16209 9055 16267 9061
rect 10226 8916 10232 8968
rect 10284 8916 10290 8968
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 14292 8965 14320 9052
rect 14826 8984 14832 9036
rect 14884 8984 14890 9036
rect 15010 8984 15016 9036
rect 15068 8984 15074 9036
rect 15223 9027 15281 9033
rect 15223 8993 15235 9027
rect 15269 9024 15281 9027
rect 16224 9024 16252 9055
rect 15269 8996 16252 9024
rect 15269 8993 15281 8996
rect 15223 8987 15281 8993
rect 10413 8959 10471 8965
rect 10413 8956 10425 8959
rect 10376 8928 10425 8956
rect 10376 8916 10382 8928
rect 10413 8925 10425 8928
rect 10459 8925 10471 8959
rect 10413 8919 10471 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14182 8848 14188 8900
rect 14240 8888 14246 8900
rect 14476 8888 14504 8919
rect 14550 8916 14556 8968
rect 14608 8916 14614 8968
rect 14737 8959 14795 8965
rect 14737 8925 14749 8959
rect 14783 8956 14795 8959
rect 14844 8956 14872 8984
rect 14783 8928 14872 8956
rect 15381 8959 15439 8965
rect 14783 8925 14795 8928
rect 14737 8919 14795 8925
rect 15381 8925 15393 8959
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15194 8888 15200 8900
rect 14240 8860 14596 8888
rect 14240 8848 14246 8860
rect 14568 8832 14596 8860
rect 14660 8860 15200 8888
rect 14660 8832 14688 8860
rect 15194 8848 15200 8860
rect 15252 8888 15258 8900
rect 15396 8888 15424 8919
rect 15252 8860 15424 8888
rect 15252 8848 15258 8860
rect 14550 8780 14556 8832
rect 14608 8780 14614 8832
rect 14642 8780 14648 8832
rect 14700 8780 14706 8832
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15488 8820 15516 8919
rect 15654 8916 15660 8968
rect 15712 8956 15718 8968
rect 15841 8959 15899 8965
rect 15841 8956 15853 8959
rect 15712 8928 15853 8956
rect 15712 8916 15718 8928
rect 15841 8925 15853 8928
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8925 16175 8959
rect 16117 8919 16175 8925
rect 16132 8888 16160 8919
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 16868 8965 16896 9064
rect 17328 8965 17356 9132
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 21637 9163 21695 9169
rect 21637 9160 21649 9163
rect 21416 9132 21649 9160
rect 21416 9120 21422 9132
rect 21637 9129 21649 9132
rect 21683 9129 21695 9163
rect 21637 9123 21695 9129
rect 23474 9120 23480 9172
rect 23532 9160 23538 9172
rect 23753 9163 23811 9169
rect 23753 9160 23765 9163
rect 23532 9132 23765 9160
rect 23532 9120 23538 9132
rect 23753 9129 23765 9132
rect 23799 9129 23811 9163
rect 23753 9123 23811 9129
rect 24118 9120 24124 9172
rect 24176 9120 24182 9172
rect 24946 9120 24952 9172
rect 25004 9120 25010 9172
rect 25774 9120 25780 9172
rect 25832 9120 25838 9172
rect 27525 9163 27583 9169
rect 27525 9129 27537 9163
rect 27571 9160 27583 9163
rect 27614 9160 27620 9172
rect 27571 9132 27620 9160
rect 27571 9129 27583 9132
rect 27525 9123 27583 9129
rect 27614 9120 27620 9132
rect 27672 9160 27678 9172
rect 27672 9132 28120 9160
rect 27672 9120 27678 9132
rect 21174 9092 21180 9104
rect 20824 9064 21180 9092
rect 16393 8959 16451 8965
rect 16393 8956 16405 8959
rect 16356 8928 16405 8956
rect 16356 8916 16362 8928
rect 16393 8925 16405 8928
rect 16439 8925 16451 8959
rect 16393 8919 16451 8925
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8956 17095 8959
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 17083 8928 17141 8956
rect 17083 8925 17095 8928
rect 17037 8919 17095 8925
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 16776 8888 16804 8919
rect 15672 8860 16804 8888
rect 15672 8829 15700 8860
rect 16776 8832 16804 8860
rect 16868 8832 16896 8919
rect 17678 8916 17684 8968
rect 17736 8916 17742 8968
rect 20824 8965 20852 9064
rect 21174 9052 21180 9064
rect 21232 9052 21238 9104
rect 23293 9095 23351 9101
rect 23293 9061 23305 9095
rect 23339 9092 23351 9095
rect 23658 9092 23664 9104
rect 23339 9064 23664 9092
rect 23339 9061 23351 9064
rect 23293 9055 23351 9061
rect 23658 9052 23664 9064
rect 23716 9092 23722 9104
rect 24136 9092 24164 9120
rect 23716 9064 24164 9092
rect 23716 9052 23722 9064
rect 20901 9027 20959 9033
rect 20901 8993 20913 9027
rect 20947 9024 20959 9027
rect 21821 9027 21879 9033
rect 21821 9024 21833 9027
rect 20947 8996 21833 9024
rect 20947 8993 20959 8996
rect 20901 8987 20959 8993
rect 21821 8993 21833 8996
rect 21867 8993 21879 9027
rect 21821 8987 21879 8993
rect 24581 9027 24639 9033
rect 24581 8993 24593 9027
rect 24627 9024 24639 9027
rect 24670 9024 24676 9036
rect 24627 8996 24676 9024
rect 24627 8993 24639 8996
rect 24581 8987 24639 8993
rect 24670 8984 24676 8996
rect 24728 8984 24734 9036
rect 20809 8959 20867 8965
rect 20809 8925 20821 8959
rect 20855 8925 20867 8959
rect 20809 8919 20867 8925
rect 20990 8916 20996 8968
rect 21048 8916 21054 8968
rect 21085 8959 21143 8965
rect 21085 8925 21097 8959
rect 21131 8956 21143 8959
rect 21174 8956 21180 8968
rect 21131 8928 21180 8956
rect 21131 8925 21143 8928
rect 21085 8919 21143 8925
rect 21174 8916 21180 8928
rect 21232 8916 21238 8968
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 21910 8916 21916 8968
rect 21968 8956 21974 8968
rect 22005 8959 22063 8965
rect 22005 8956 22017 8959
rect 21968 8928 22017 8956
rect 21968 8916 21974 8928
rect 22005 8925 22017 8928
rect 22051 8925 22063 8959
rect 22005 8919 22063 8925
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24210 8956 24216 8968
rect 23891 8928 24216 8956
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 24210 8916 24216 8928
rect 24268 8916 24274 8968
rect 24486 8916 24492 8968
rect 24544 8916 24550 8968
rect 24765 8959 24823 8965
rect 24765 8925 24777 8959
rect 24811 8925 24823 8959
rect 24765 8919 24823 8925
rect 17586 8848 17592 8900
rect 17644 8848 17650 8900
rect 21008 8888 21036 8916
rect 21269 8891 21327 8897
rect 21269 8888 21281 8891
rect 21008 8860 21281 8888
rect 21269 8857 21281 8860
rect 21315 8857 21327 8891
rect 21269 8851 21327 8857
rect 21361 8891 21419 8897
rect 21361 8857 21373 8891
rect 21407 8857 21419 8891
rect 24504 8888 24532 8916
rect 24780 8888 24808 8919
rect 25222 8916 25228 8968
rect 25280 8916 25286 8968
rect 25409 8959 25467 8965
rect 25409 8925 25421 8959
rect 25455 8956 25467 8959
rect 25792 8956 25820 9120
rect 27157 9095 27215 9101
rect 27157 9061 27169 9095
rect 27203 9092 27215 9095
rect 27706 9092 27712 9104
rect 27203 9064 27712 9092
rect 27203 9061 27215 9064
rect 27157 9055 27215 9061
rect 27706 9052 27712 9064
rect 27764 9092 27770 9104
rect 27982 9092 27988 9104
rect 27764 9064 27988 9092
rect 27764 9052 27770 9064
rect 27982 9052 27988 9064
rect 28040 9052 28046 9104
rect 25455 8928 25820 8956
rect 25455 8925 25467 8928
rect 25409 8919 25467 8925
rect 27890 8916 27896 8968
rect 27948 8916 27954 8968
rect 28092 8965 28120 9132
rect 28077 8959 28135 8965
rect 28077 8925 28089 8959
rect 28123 8925 28135 8959
rect 28077 8919 28135 8925
rect 24504 8860 24808 8888
rect 27525 8891 27583 8897
rect 21361 8851 21419 8857
rect 27525 8857 27537 8891
rect 27571 8888 27583 8891
rect 27798 8888 27804 8900
rect 27571 8860 27804 8888
rect 27571 8857 27583 8860
rect 27525 8851 27583 8857
rect 14792 8792 15516 8820
rect 15657 8823 15715 8829
rect 14792 8780 14798 8792
rect 15657 8789 15669 8823
rect 15703 8789 15715 8823
rect 15657 8783 15715 8789
rect 16758 8780 16764 8832
rect 16816 8780 16822 8832
rect 16850 8780 16856 8832
rect 16908 8780 16914 8832
rect 21174 8780 21180 8832
rect 21232 8820 21238 8832
rect 21376 8820 21404 8851
rect 27798 8848 27804 8860
rect 27856 8848 27862 8900
rect 21232 8792 21404 8820
rect 21232 8780 21238 8792
rect 22186 8780 22192 8832
rect 22244 8780 22250 8832
rect 23934 8780 23940 8832
rect 23992 8820 23998 8832
rect 24213 8823 24271 8829
rect 24213 8820 24225 8823
rect 23992 8792 24225 8820
rect 23992 8780 23998 8792
rect 24213 8789 24225 8792
rect 24259 8820 24271 8823
rect 24578 8820 24584 8832
rect 24259 8792 24584 8820
rect 24259 8789 24271 8792
rect 24213 8783 24271 8789
rect 24578 8780 24584 8792
rect 24636 8780 24642 8832
rect 25317 8823 25375 8829
rect 25317 8789 25329 8823
rect 25363 8820 25375 8823
rect 25866 8820 25872 8832
rect 25363 8792 25872 8820
rect 25363 8789 25375 8792
rect 25317 8783 25375 8789
rect 25866 8780 25872 8792
rect 25924 8780 25930 8832
rect 27709 8823 27767 8829
rect 27709 8789 27721 8823
rect 27755 8820 27767 8823
rect 27982 8820 27988 8832
rect 27755 8792 27988 8820
rect 27755 8789 27767 8792
rect 27709 8783 27767 8789
rect 27982 8780 27988 8792
rect 28040 8780 28046 8832
rect 28902 8780 28908 8832
rect 28960 8780 28966 8832
rect 1104 8730 35236 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 35236 8730
rect 1104 8656 35236 8678
rect 10226 8576 10232 8628
rect 10284 8616 10290 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 10284 8588 10517 8616
rect 10284 8576 10290 8588
rect 10505 8585 10517 8588
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 10704 8588 11836 8616
rect 6825 8551 6883 8557
rect 6825 8517 6837 8551
rect 6871 8548 6883 8551
rect 7742 8548 7748 8560
rect 6871 8520 7748 8548
rect 6871 8517 6883 8520
rect 6825 8511 6883 8517
rect 7742 8508 7748 8520
rect 7800 8508 7806 8560
rect 7852 8520 8800 8548
rect 7282 8440 7288 8492
rect 7340 8440 7346 8492
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 7852 8489 7880 8520
rect 8772 8492 8800 8520
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9272 8520 9444 8548
rect 9272 8508 9278 8520
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 7837 8443 7895 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8480 8079 8483
rect 8067 8452 8156 8480
rect 8067 8449 8079 8452
rect 8021 8443 8079 8449
rect 8128 8344 8156 8452
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9416 8489 9444 8520
rect 10704 8489 10732 8588
rect 11808 8548 11836 8588
rect 11974 8576 11980 8628
rect 12032 8616 12038 8628
rect 12032 8588 13124 8616
rect 12032 8576 12038 8588
rect 11164 8520 11744 8548
rect 11808 8520 11928 8548
rect 9401 8483 9459 8489
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 9401 8443 9459 8449
rect 9600 8452 10701 8480
rect 9600 8356 9628 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 10689 8443 10747 8449
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8449 11023 8483
rect 10965 8443 11023 8449
rect 10134 8372 10140 8424
rect 10192 8372 10198 8424
rect 10870 8412 10876 8424
rect 10244 8384 10876 8412
rect 10244 8356 10272 8384
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 10980 8412 11008 8443
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11164 8489 11192 8520
rect 11149 8483 11207 8489
rect 11149 8480 11161 8483
rect 11112 8452 11161 8480
rect 11112 8440 11118 8452
rect 11149 8449 11161 8452
rect 11195 8449 11207 8483
rect 11149 8443 11207 8449
rect 11514 8440 11520 8492
rect 11572 8440 11578 8492
rect 11716 8489 11744 8520
rect 11900 8489 11928 8520
rect 12066 8508 12072 8560
rect 12124 8548 12130 8560
rect 12161 8551 12219 8557
rect 12161 8548 12173 8551
rect 12124 8520 12173 8548
rect 12124 8508 12130 8520
rect 12161 8517 12173 8520
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 13096 8492 13124 8588
rect 14642 8576 14648 8628
rect 14700 8576 14706 8628
rect 14734 8576 14740 8628
rect 14792 8576 14798 8628
rect 15378 8576 15384 8628
rect 15436 8616 15442 8628
rect 15562 8616 15568 8628
rect 15436 8588 15568 8616
rect 15436 8576 15442 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 18874 8576 18880 8628
rect 18932 8576 18938 8628
rect 19889 8619 19947 8625
rect 19889 8585 19901 8619
rect 19935 8616 19947 8619
rect 19978 8616 19984 8628
rect 19935 8588 19984 8616
rect 19935 8585 19947 8588
rect 19889 8579 19947 8585
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 23658 8576 23664 8628
rect 23716 8576 23722 8628
rect 27173 8619 27231 8625
rect 27173 8616 27185 8619
rect 26528 8588 27185 8616
rect 11701 8483 11759 8489
rect 11701 8449 11713 8483
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8449 11851 8483
rect 11793 8443 11851 8449
rect 11886 8483 11944 8489
rect 11886 8449 11898 8483
rect 11932 8480 11944 8483
rect 11932 8452 12434 8480
rect 11932 8449 11944 8452
rect 11886 8443 11944 8449
rect 11532 8412 11560 8440
rect 10980 8384 11560 8412
rect 8128 8316 8340 8344
rect 8312 8276 8340 8316
rect 9122 8304 9128 8356
rect 9180 8344 9186 8356
rect 9180 8316 9536 8344
rect 9180 8304 9186 8316
rect 8846 8276 8852 8288
rect 8312 8248 8852 8276
rect 8846 8236 8852 8248
rect 8904 8236 8910 8288
rect 9508 8276 9536 8316
rect 9582 8304 9588 8356
rect 9640 8304 9646 8356
rect 10226 8304 10232 8356
rect 10284 8304 10290 8356
rect 10781 8347 10839 8353
rect 10781 8344 10793 8347
rect 10336 8316 10793 8344
rect 10336 8276 10364 8316
rect 10781 8313 10793 8316
rect 10827 8344 10839 8347
rect 11808 8344 11836 8443
rect 12406 8356 12434 8452
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12584 8452 12725 8480
rect 12584 8440 12590 8452
rect 12713 8449 12725 8452
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14660 8489 14688 8576
rect 17494 8508 17500 8560
rect 17552 8508 17558 8560
rect 18892 8548 18920 8576
rect 18708 8520 18920 8548
rect 23676 8548 23704 8576
rect 26528 8560 26556 8588
rect 27173 8585 27185 8588
rect 27219 8585 27231 8619
rect 27173 8579 27231 8585
rect 27341 8619 27399 8625
rect 27341 8585 27353 8619
rect 27387 8585 27399 8619
rect 27341 8579 27399 8585
rect 27525 8619 27583 8625
rect 27525 8585 27537 8619
rect 27571 8616 27583 8619
rect 27614 8616 27620 8628
rect 27571 8588 27620 8616
rect 27571 8585 27583 8588
rect 27525 8579 27583 8585
rect 23676 8520 24072 8548
rect 16856 8492 16908 8498
rect 18708 8492 18736 8520
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8449 14703 8483
rect 14645 8443 14703 8449
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 16758 8440 16764 8492
rect 16816 8440 16822 8492
rect 18690 8440 18696 8492
rect 18748 8440 18754 8492
rect 18874 8440 18880 8492
rect 18932 8440 18938 8492
rect 18966 8440 18972 8492
rect 19024 8440 19030 8492
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 20530 8480 20536 8492
rect 19383 8452 20536 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 23566 8440 23572 8492
rect 23624 8480 23630 8492
rect 23845 8483 23903 8489
rect 23845 8480 23857 8483
rect 23624 8452 23857 8480
rect 23624 8440 23630 8452
rect 23845 8449 23857 8452
rect 23891 8480 23903 8483
rect 23934 8480 23940 8492
rect 23891 8452 23940 8480
rect 23891 8449 23903 8452
rect 23845 8443 23903 8449
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 24044 8489 24072 8520
rect 26510 8508 26516 8560
rect 26568 8508 26574 8560
rect 26697 8551 26755 8557
rect 26697 8517 26709 8551
rect 26743 8548 26755 8551
rect 26970 8548 26976 8560
rect 26743 8520 26976 8548
rect 26743 8517 26755 8520
rect 26697 8511 26755 8517
rect 24029 8483 24087 8489
rect 24029 8449 24041 8483
rect 24075 8449 24087 8483
rect 24029 8443 24087 8449
rect 24854 8440 24860 8492
rect 24912 8480 24918 8492
rect 25041 8483 25099 8489
rect 25041 8480 25053 8483
rect 24912 8452 25053 8480
rect 24912 8440 24918 8452
rect 25041 8449 25053 8452
rect 25087 8449 25099 8483
rect 25041 8443 25099 8449
rect 25222 8440 25228 8492
rect 25280 8440 25286 8492
rect 25774 8440 25780 8492
rect 25832 8480 25838 8492
rect 26712 8480 26740 8511
rect 26970 8508 26976 8520
rect 27028 8508 27034 8560
rect 27062 8508 27068 8560
rect 27120 8548 27126 8560
rect 27356 8548 27384 8579
rect 27614 8576 27620 8588
rect 27672 8576 27678 8628
rect 27890 8576 27896 8628
rect 27948 8616 27954 8628
rect 28077 8619 28135 8625
rect 28077 8616 28089 8619
rect 27948 8588 28089 8616
rect 27948 8576 27954 8588
rect 28077 8585 28089 8588
rect 28123 8585 28135 8619
rect 28077 8579 28135 8585
rect 27120 8520 27476 8548
rect 27120 8508 27126 8520
rect 25832 8452 26740 8480
rect 26789 8483 26847 8489
rect 25832 8440 25838 8452
rect 26789 8449 26801 8483
rect 26835 8480 26847 8483
rect 27338 8480 27344 8492
rect 26835 8452 27344 8480
rect 26835 8449 26847 8452
rect 26789 8443 26847 8449
rect 27338 8440 27344 8452
rect 27396 8440 27402 8492
rect 27448 8489 27476 8520
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 27617 8483 27675 8489
rect 27617 8449 27629 8483
rect 27663 8449 27675 8483
rect 27617 8443 27675 8449
rect 11974 8344 11980 8356
rect 10827 8316 11980 8344
rect 10827 8313 10839 8316
rect 10781 8307 10839 8313
rect 11974 8304 11980 8316
rect 12032 8304 12038 8356
rect 12342 8304 12348 8356
rect 12400 8344 12434 8356
rect 14200 8344 14228 8440
rect 16856 8434 16908 8440
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8412 14611 8415
rect 15102 8412 15108 8424
rect 14599 8384 15108 8412
rect 14599 8381 14611 8384
rect 14553 8375 14611 8381
rect 15102 8372 15108 8384
rect 15160 8412 15166 8424
rect 15654 8412 15660 8424
rect 15160 8384 15660 8412
rect 15160 8372 15166 8384
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 19978 8372 19984 8424
rect 20036 8412 20042 8424
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 20036 8384 20085 8412
rect 20036 8372 20042 8384
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 20162 8372 20168 8424
rect 20220 8372 20226 8424
rect 24213 8415 24271 8421
rect 24213 8381 24225 8415
rect 24259 8412 24271 8415
rect 24946 8412 24952 8424
rect 24259 8384 24952 8412
rect 24259 8381 24271 8384
rect 24213 8375 24271 8381
rect 24946 8372 24952 8384
rect 25004 8412 25010 8424
rect 25792 8412 25820 8440
rect 27632 8412 27660 8443
rect 27706 8440 27712 8492
rect 27764 8440 27770 8492
rect 27798 8440 27804 8492
rect 27856 8480 27862 8492
rect 27856 8452 27901 8480
rect 27856 8440 27862 8452
rect 25004 8384 25820 8412
rect 26528 8384 27660 8412
rect 25004 8372 25010 8384
rect 12400 8316 14228 8344
rect 14921 8347 14979 8353
rect 12400 8304 12406 8316
rect 14921 8313 14933 8347
rect 14967 8344 14979 8347
rect 15286 8344 15292 8356
rect 14967 8316 15292 8344
rect 14967 8313 14979 8316
rect 14921 8307 14979 8313
rect 15286 8304 15292 8316
rect 15344 8304 15350 8356
rect 25314 8344 25320 8356
rect 16592 8316 16988 8344
rect 9508 8248 10364 8276
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 16592 8276 16620 8316
rect 12676 8248 16620 8276
rect 16960 8276 16988 8316
rect 24596 8316 25320 8344
rect 24596 8288 24624 8316
rect 25314 8304 25320 8316
rect 25372 8344 25378 8356
rect 26528 8353 26556 8384
rect 25501 8347 25559 8353
rect 25501 8344 25513 8347
rect 25372 8316 25513 8344
rect 25372 8304 25378 8316
rect 25501 8313 25513 8316
rect 25547 8313 25559 8347
rect 25501 8307 25559 8313
rect 26513 8347 26571 8353
rect 26513 8313 26525 8347
rect 26559 8313 26571 8347
rect 26513 8307 26571 8313
rect 23014 8276 23020 8288
rect 16960 8248 23020 8276
rect 12676 8236 12682 8248
rect 23014 8236 23020 8248
rect 23072 8276 23078 8288
rect 24489 8279 24547 8285
rect 24489 8276 24501 8279
rect 23072 8248 24501 8276
rect 23072 8236 23078 8248
rect 24489 8245 24501 8248
rect 24535 8276 24547 8279
rect 24578 8276 24584 8288
rect 24535 8248 24584 8276
rect 24535 8245 24547 8248
rect 24489 8239 24547 8245
rect 24578 8236 24584 8248
rect 24636 8236 24642 8288
rect 25222 8236 25228 8288
rect 25280 8236 25286 8288
rect 27157 8279 27215 8285
rect 27157 8245 27169 8279
rect 27203 8276 27215 8279
rect 27246 8276 27252 8288
rect 27203 8248 27252 8276
rect 27203 8245 27215 8248
rect 27157 8239 27215 8245
rect 27246 8236 27252 8248
rect 27304 8236 27310 8288
rect 1104 8186 35248 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 35248 8186
rect 1104 8112 35248 8134
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 12250 8072 12256 8084
rect 11572 8044 12256 8072
rect 11572 8032 11578 8044
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12437 8075 12495 8081
rect 12437 8041 12449 8075
rect 12483 8072 12495 8075
rect 12526 8072 12532 8084
rect 12483 8044 12532 8072
rect 12483 8041 12495 8044
rect 12437 8035 12495 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 19061 8075 19119 8081
rect 19061 8041 19073 8075
rect 19107 8072 19119 8075
rect 19978 8072 19984 8084
rect 19107 8044 19984 8072
rect 19107 8041 19119 8044
rect 19061 8035 19119 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20088 8044 23152 8072
rect 11054 8004 11060 8016
rect 7300 7976 11060 8004
rect 7300 7948 7328 7976
rect 7282 7896 7288 7948
rect 7340 7896 7346 7948
rect 9214 7896 9220 7948
rect 9272 7896 9278 7948
rect 9508 7945 9536 7976
rect 11054 7964 11060 7976
rect 11112 8004 11118 8016
rect 11112 7976 11284 8004
rect 11112 7964 11118 7976
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 11146 7936 11152 7948
rect 9493 7899 9551 7905
rect 9600 7908 11152 7936
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 9600 7877 9628 7908
rect 11146 7896 11152 7908
rect 11204 7896 11210 7948
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 7616 7840 9597 7868
rect 7616 7828 7622 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 9953 7831 10011 7837
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7837 10195 7871
rect 10137 7831 10195 7837
rect 10413 7871 10471 7877
rect 10413 7837 10425 7871
rect 10459 7868 10471 7871
rect 10502 7868 10508 7880
rect 10459 7840 10508 7868
rect 10459 7837 10471 7840
rect 10413 7831 10471 7837
rect 8846 7760 8852 7812
rect 8904 7800 8910 7812
rect 9968 7800 9996 7831
rect 8904 7772 9996 7800
rect 8904 7760 8910 7772
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10152 7732 10180 7831
rect 10502 7828 10508 7840
rect 10560 7828 10566 7880
rect 10594 7828 10600 7880
rect 10652 7828 10658 7880
rect 10686 7760 10692 7812
rect 10744 7760 10750 7812
rect 11256 7800 11284 7976
rect 12544 7936 12572 8032
rect 20088 8004 20116 8044
rect 13648 7976 20116 8004
rect 12897 7939 12955 7945
rect 12544 7908 12848 7936
rect 12342 7868 12348 7880
rect 12268 7840 12348 7868
rect 12066 7800 12072 7812
rect 11256 7772 12072 7800
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 12268 7809 12296 7840
rect 12342 7828 12348 7840
rect 12400 7828 12406 7880
rect 12820 7854 12848 7908
rect 12897 7905 12909 7939
rect 12943 7936 12955 7939
rect 13078 7936 13084 7948
rect 12943 7908 13084 7936
rect 12943 7905 12955 7908
rect 12897 7899 12955 7905
rect 13078 7896 13084 7908
rect 13136 7896 13142 7948
rect 12253 7803 12311 7809
rect 12253 7769 12265 7803
rect 12299 7769 12311 7803
rect 13648 7800 13676 7976
rect 20162 7964 20168 8016
rect 20220 8004 20226 8016
rect 20220 7976 20760 8004
rect 20220 7964 20226 7976
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7936 13783 7939
rect 14366 7936 14372 7948
rect 13771 7908 14372 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 15102 7936 15108 7948
rect 14424 7908 15108 7936
rect 14424 7896 14430 7908
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7936 18383 7939
rect 18874 7936 18880 7948
rect 18371 7908 18880 7936
rect 18371 7905 18383 7908
rect 18325 7899 18383 7905
rect 18874 7896 18880 7908
rect 18932 7896 18938 7948
rect 18966 7896 18972 7948
rect 19024 7896 19030 7948
rect 20438 7936 20444 7948
rect 20088 7908 20444 7936
rect 14734 7828 14740 7880
rect 14792 7868 14798 7880
rect 15013 7871 15071 7877
rect 15013 7868 15025 7871
rect 14792 7840 15025 7868
rect 14792 7828 14798 7840
rect 15013 7837 15025 7840
rect 15059 7837 15071 7871
rect 15013 7831 15071 7837
rect 12253 7763 12311 7769
rect 12406 7772 13676 7800
rect 15028 7800 15056 7831
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 15289 7871 15347 7877
rect 15289 7868 15301 7871
rect 15252 7840 15301 7868
rect 15252 7828 15258 7840
rect 15289 7837 15301 7840
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 15473 7871 15531 7877
rect 15473 7837 15485 7871
rect 15519 7837 15531 7871
rect 15473 7831 15531 7837
rect 15488 7800 15516 7831
rect 17586 7828 17592 7880
rect 17644 7828 17650 7880
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7868 17923 7871
rect 17954 7868 17960 7880
rect 17911 7840 17960 7868
rect 17911 7837 17923 7840
rect 17865 7831 17923 7837
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 18690 7868 18696 7880
rect 18463 7840 18696 7868
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 15028 7772 15516 7800
rect 17604 7800 17632 7828
rect 18156 7800 18184 7831
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7868 18843 7871
rect 18984 7868 19012 7896
rect 18831 7840 19012 7868
rect 19797 7871 19855 7877
rect 18831 7837 18843 7840
rect 18785 7831 18843 7837
rect 19797 7837 19809 7871
rect 19843 7868 19855 7871
rect 19886 7868 19892 7880
rect 19843 7840 19892 7868
rect 19843 7837 19855 7840
rect 19797 7831 19855 7837
rect 19886 7828 19892 7840
rect 19944 7828 19950 7880
rect 20088 7877 20116 7908
rect 20438 7896 20444 7908
rect 20496 7896 20502 7948
rect 20533 7939 20591 7945
rect 20533 7905 20545 7939
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20162 7828 20168 7880
rect 20220 7828 20226 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20346 7868 20352 7880
rect 20303 7840 20352 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 20346 7828 20352 7840
rect 20404 7828 20410 7880
rect 17604 7772 18184 7800
rect 20548 7800 20576 7899
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 20732 7868 20760 7976
rect 21450 7936 21456 7948
rect 21100 7908 21456 7936
rect 20898 7868 20904 7880
rect 20732 7840 20904 7868
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 21100 7800 21128 7908
rect 21450 7896 21456 7908
rect 21508 7936 21514 7948
rect 21508 7908 21680 7936
rect 21508 7896 21514 7908
rect 21174 7828 21180 7880
rect 21232 7868 21238 7880
rect 21232 7840 21312 7868
rect 21232 7828 21238 7840
rect 20548 7772 21128 7800
rect 21284 7800 21312 7840
rect 21358 7828 21364 7880
rect 21416 7828 21422 7880
rect 21652 7877 21680 7908
rect 23124 7877 23152 8044
rect 23290 8032 23296 8084
rect 23348 8032 23354 8084
rect 25130 8072 25136 8084
rect 24780 8044 25136 8072
rect 24780 8013 24808 8044
rect 25130 8032 25136 8044
rect 25188 8032 25194 8084
rect 25409 8075 25467 8081
rect 25409 8041 25421 8075
rect 25455 8072 25467 8075
rect 25682 8072 25688 8084
rect 25455 8044 25688 8072
rect 25455 8041 25467 8044
rect 25409 8035 25467 8041
rect 25682 8032 25688 8044
rect 25740 8032 25746 8084
rect 25869 8075 25927 8081
rect 25869 8041 25881 8075
rect 25915 8041 25927 8075
rect 25869 8035 25927 8041
rect 23385 8007 23443 8013
rect 23385 7973 23397 8007
rect 23431 8004 23443 8007
rect 24765 8007 24823 8013
rect 23431 7976 24716 8004
rect 23431 7973 23443 7976
rect 23385 7967 23443 7973
rect 23477 7939 23535 7945
rect 23477 7905 23489 7939
rect 23523 7936 23535 7939
rect 23569 7939 23627 7945
rect 23569 7936 23581 7939
rect 23523 7908 23581 7936
rect 23523 7905 23535 7908
rect 23477 7899 23535 7905
rect 23569 7905 23581 7908
rect 23615 7905 23627 7939
rect 23569 7899 23627 7905
rect 23658 7896 23664 7948
rect 23716 7896 23722 7948
rect 24688 7936 24716 7976
rect 24765 7973 24777 8007
rect 24811 7973 24823 8007
rect 24765 7967 24823 7973
rect 24854 7964 24860 8016
rect 24912 7964 24918 8016
rect 25884 8004 25912 8035
rect 25958 8032 25964 8084
rect 26016 8072 26022 8084
rect 26016 8044 26280 8072
rect 26016 8032 26022 8044
rect 25056 7976 26188 8004
rect 25056 7936 25084 7976
rect 23859 7908 24624 7936
rect 24688 7908 25084 7936
rect 25133 7939 25191 7945
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7837 21695 7871
rect 21637 7831 21695 7837
rect 21821 7871 21879 7877
rect 21821 7837 21833 7871
rect 21867 7837 21879 7871
rect 21821 7831 21879 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 23155 7840 23213 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23201 7837 23213 7840
rect 23247 7868 23259 7871
rect 23676 7868 23704 7896
rect 23859 7877 23887 7908
rect 24596 7880 24624 7908
rect 25133 7905 25145 7939
rect 25179 7936 25191 7939
rect 25958 7936 25964 7948
rect 25179 7908 25964 7936
rect 25179 7905 25191 7908
rect 25133 7899 25191 7905
rect 25958 7896 25964 7908
rect 26016 7896 26022 7948
rect 23247 7840 23704 7868
rect 23844 7871 23902 7877
rect 23247 7837 23259 7840
rect 23201 7831 23259 7837
rect 23844 7837 23856 7871
rect 23890 7837 23902 7871
rect 23844 7831 23902 7837
rect 21836 7800 21864 7831
rect 23934 7828 23940 7880
rect 23992 7828 23998 7880
rect 24489 7871 24547 7877
rect 24489 7837 24501 7871
rect 24535 7837 24547 7871
rect 24489 7831 24547 7837
rect 24504 7800 24532 7831
rect 24578 7828 24584 7880
rect 24636 7868 24642 7880
rect 24673 7871 24731 7877
rect 24673 7868 24685 7871
rect 24636 7840 24685 7868
rect 24636 7828 24642 7840
rect 24673 7837 24685 7840
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 24946 7828 24952 7880
rect 25004 7828 25010 7880
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7837 25283 7871
rect 25225 7831 25283 7837
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7868 25559 7871
rect 25774 7868 25780 7880
rect 25547 7840 25780 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 21284 7772 21864 7800
rect 23860 7772 24532 7800
rect 9824 7704 10180 7732
rect 9824 7692 9830 7704
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 12406 7732 12434 7772
rect 23860 7744 23888 7772
rect 11388 7704 12434 7732
rect 11388 7692 11394 7704
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 15013 7735 15071 7741
rect 15013 7732 15025 7735
rect 14792 7704 15025 7732
rect 14792 7692 14798 7704
rect 15013 7701 15025 7704
rect 15059 7701 15071 7735
rect 15013 7695 15071 7701
rect 15378 7692 15384 7744
rect 15436 7692 15442 7744
rect 17957 7735 18015 7741
rect 17957 7701 17969 7735
rect 18003 7732 18015 7735
rect 18322 7732 18328 7744
rect 18003 7704 18328 7732
rect 18003 7701 18015 7704
rect 17957 7695 18015 7701
rect 18322 7692 18328 7704
rect 18380 7692 18386 7744
rect 19889 7735 19947 7741
rect 19889 7701 19901 7735
rect 19935 7732 19947 7735
rect 20254 7732 20260 7744
rect 19935 7704 20260 7732
rect 19935 7701 19947 7704
rect 19889 7695 19947 7701
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 20530 7692 20536 7744
rect 20588 7732 20594 7744
rect 20717 7735 20775 7741
rect 20717 7732 20729 7735
rect 20588 7704 20729 7732
rect 20588 7692 20594 7704
rect 20717 7701 20729 7704
rect 20763 7701 20775 7735
rect 20717 7695 20775 7701
rect 21082 7692 21088 7744
rect 21140 7692 21146 7744
rect 21266 7692 21272 7744
rect 21324 7692 21330 7744
rect 21818 7692 21824 7744
rect 21876 7692 21882 7744
rect 23842 7692 23848 7744
rect 23900 7692 23906 7744
rect 24504 7732 24532 7772
rect 25242 7732 25270 7831
rect 25774 7828 25780 7840
rect 25832 7828 25838 7880
rect 26160 7877 26188 7976
rect 26145 7871 26203 7877
rect 26145 7837 26157 7871
rect 26191 7837 26203 7871
rect 26252 7868 26280 8044
rect 26510 8032 26516 8084
rect 26568 8032 26574 8084
rect 26421 8007 26479 8013
rect 26421 7973 26433 8007
rect 26467 7973 26479 8007
rect 26421 7967 26479 7973
rect 26436 7868 26464 7967
rect 26513 7871 26571 7877
rect 26513 7868 26525 7871
rect 26252 7840 26372 7868
rect 26436 7840 26525 7868
rect 26145 7831 26203 7837
rect 25314 7760 25320 7812
rect 25372 7760 25378 7812
rect 25682 7760 25688 7812
rect 25740 7800 25746 7812
rect 26237 7803 26295 7809
rect 26237 7800 26249 7803
rect 25740 7772 26249 7800
rect 25740 7760 25746 7772
rect 26237 7769 26249 7772
rect 26283 7769 26295 7803
rect 26344 7800 26372 7840
rect 26513 7837 26525 7840
rect 26559 7837 26571 7871
rect 26513 7831 26571 7837
rect 26697 7871 26755 7877
rect 26697 7837 26709 7871
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 26421 7803 26479 7809
rect 26421 7800 26433 7803
rect 26344 7772 26433 7800
rect 26237 7763 26295 7769
rect 26421 7769 26433 7772
rect 26467 7769 26479 7803
rect 26712 7800 26740 7831
rect 26421 7763 26479 7769
rect 26528 7772 26740 7800
rect 26528 7744 26556 7772
rect 24504 7704 25270 7732
rect 25866 7692 25872 7744
rect 25924 7741 25930 7744
rect 25924 7735 25943 7741
rect 25931 7701 25943 7735
rect 25924 7695 25943 7701
rect 26053 7735 26111 7741
rect 26053 7701 26065 7735
rect 26099 7732 26111 7735
rect 26510 7732 26516 7744
rect 26099 7704 26516 7732
rect 26099 7701 26111 7704
rect 26053 7695 26111 7701
rect 25924 7692 25930 7695
rect 26510 7692 26516 7704
rect 26568 7692 26574 7744
rect 1104 7642 35236 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 35236 7642
rect 1104 7568 35236 7590
rect 16022 7488 16028 7540
rect 16080 7528 16086 7540
rect 16117 7531 16175 7537
rect 16117 7528 16129 7531
rect 16080 7500 16129 7528
rect 16080 7488 16086 7500
rect 16117 7497 16129 7500
rect 16163 7528 16175 7531
rect 16390 7528 16396 7540
rect 16163 7500 16396 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 18509 7531 18567 7537
rect 18509 7497 18521 7531
rect 18555 7528 18567 7531
rect 18966 7528 18972 7540
rect 18555 7500 18972 7528
rect 18555 7497 18567 7500
rect 18509 7491 18567 7497
rect 18966 7488 18972 7500
rect 19024 7488 19030 7540
rect 20254 7488 20260 7540
rect 20312 7488 20318 7540
rect 20530 7528 20536 7540
rect 20364 7500 20536 7528
rect 10594 7460 10600 7472
rect 10336 7432 10600 7460
rect 8478 7352 8484 7404
rect 8536 7392 8542 7404
rect 8846 7392 8852 7404
rect 8536 7364 8852 7392
rect 8536 7352 8542 7364
rect 8846 7352 8852 7364
rect 8904 7352 8910 7404
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 10336 7401 10364 7432
rect 10594 7420 10600 7432
rect 10652 7460 10658 7472
rect 10652 7432 11008 7460
rect 10652 7420 10658 7432
rect 10980 7404 11008 7432
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 14366 7460 14372 7472
rect 12124 7432 13584 7460
rect 12124 7420 12130 7432
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10502 7352 10508 7404
rect 10560 7392 10566 7404
rect 10689 7395 10747 7401
rect 10689 7392 10701 7395
rect 10560 7364 10701 7392
rect 10560 7352 10566 7364
rect 10689 7361 10701 7364
rect 10735 7361 10747 7395
rect 10689 7355 10747 7361
rect 10962 7352 10968 7404
rect 11020 7352 11026 7404
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7392 12679 7395
rect 12802 7392 12808 7404
rect 12667 7364 12808 7392
rect 12667 7361 12679 7364
rect 12621 7355 12679 7361
rect 12802 7352 12808 7364
rect 12860 7352 12866 7404
rect 12897 7395 12955 7401
rect 12897 7361 12909 7395
rect 12943 7392 12955 7395
rect 12986 7392 12992 7404
rect 12943 7364 12992 7392
rect 12943 7361 12955 7364
rect 12897 7355 12955 7361
rect 12986 7352 12992 7364
rect 13044 7392 13050 7404
rect 13446 7392 13452 7404
rect 13044 7364 13452 7392
rect 13044 7352 13050 7364
rect 13446 7352 13452 7364
rect 13504 7352 13510 7404
rect 13556 7401 13584 7432
rect 14200 7432 14372 7460
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7361 13599 7395
rect 13541 7355 13599 7361
rect 10410 7284 10416 7336
rect 10468 7284 10474 7336
rect 10594 7284 10600 7336
rect 10652 7324 10658 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10652 7296 11069 7324
rect 10652 7284 10658 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 12434 7284 12440 7336
rect 12492 7324 12498 7336
rect 12713 7327 12771 7333
rect 12713 7324 12725 7327
rect 12492 7296 12725 7324
rect 12492 7284 12498 7296
rect 12713 7293 12725 7296
rect 12759 7293 12771 7327
rect 12713 7287 12771 7293
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7293 13323 7327
rect 13265 7287 13323 7293
rect 9306 7216 9312 7268
rect 9364 7216 9370 7268
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 12342 7256 12348 7268
rect 11204 7228 12348 7256
rect 11204 7216 11210 7228
rect 12342 7216 12348 7228
rect 12400 7256 12406 7268
rect 13081 7259 13139 7265
rect 12400 7228 12848 7256
rect 12400 7216 12406 7228
rect 12710 7148 12716 7200
rect 12768 7148 12774 7200
rect 12820 7188 12848 7228
rect 13081 7225 13093 7259
rect 13127 7256 13139 7259
rect 13280 7256 13308 7287
rect 14200 7265 14228 7432
rect 14366 7420 14372 7432
rect 14424 7460 14430 7472
rect 14424 7432 15240 7460
rect 14424 7420 14430 7432
rect 14734 7352 14740 7404
rect 14792 7392 14798 7404
rect 14829 7395 14887 7401
rect 14829 7392 14841 7395
rect 14792 7364 14841 7392
rect 14792 7352 14798 7364
rect 14829 7361 14841 7364
rect 14875 7361 14887 7395
rect 14829 7355 14887 7361
rect 15102 7352 15108 7404
rect 15160 7352 15166 7404
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 13127 7228 13308 7256
rect 14185 7259 14243 7265
rect 13127 7225 13139 7228
rect 13081 7219 13139 7225
rect 14185 7225 14197 7259
rect 14231 7225 14243 7259
rect 14185 7219 14243 7225
rect 14476 7188 14504 7287
rect 14918 7284 14924 7336
rect 14976 7284 14982 7336
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7293 15071 7327
rect 15212 7324 15240 7432
rect 15378 7420 15384 7472
rect 15436 7460 15442 7472
rect 15436 7432 16068 7460
rect 15436 7420 15442 7432
rect 16040 7401 16068 7432
rect 17586 7420 17592 7472
rect 17644 7460 17650 7472
rect 18233 7463 18291 7469
rect 18233 7460 18245 7463
rect 17644 7432 18245 7460
rect 17644 7420 17650 7432
rect 18233 7429 18245 7432
rect 18279 7429 18291 7463
rect 18233 7423 18291 7429
rect 18322 7420 18328 7472
rect 18380 7460 18386 7472
rect 18380 7432 18552 7460
rect 18380 7420 18386 7432
rect 16025 7395 16083 7401
rect 16025 7361 16037 7395
rect 16071 7392 16083 7395
rect 16114 7392 16120 7404
rect 16071 7364 16120 7392
rect 16071 7361 16083 7364
rect 16025 7355 16083 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7392 16359 7395
rect 16761 7395 16819 7401
rect 16761 7392 16773 7395
rect 16347 7364 16773 7392
rect 16347 7361 16359 7364
rect 16301 7355 16359 7361
rect 16761 7361 16773 7364
rect 16807 7361 16819 7395
rect 16761 7355 16819 7361
rect 17129 7395 17187 7401
rect 17129 7361 17141 7395
rect 17175 7392 17187 7395
rect 17494 7392 17500 7404
rect 17175 7364 17500 7392
rect 17175 7361 17187 7364
rect 17129 7355 17187 7361
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 18414 7352 18420 7404
rect 18472 7352 18478 7404
rect 18524 7401 18552 7432
rect 18509 7395 18567 7401
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 20257 7395 20315 7401
rect 20257 7361 20269 7395
rect 20303 7392 20315 7395
rect 20364 7392 20392 7500
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20864 7500 21220 7528
rect 20864 7488 20870 7500
rect 20622 7460 20628 7472
rect 20456 7432 20628 7460
rect 20456 7401 20484 7432
rect 20622 7420 20628 7432
rect 20680 7420 20686 7472
rect 20898 7420 20904 7472
rect 20956 7420 20962 7472
rect 20899 7417 20957 7420
rect 20303 7364 20392 7392
rect 20441 7395 20499 7401
rect 20303 7361 20315 7364
rect 20257 7355 20315 7361
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7361 20867 7395
rect 20899 7383 20911 7417
rect 20945 7383 20957 7417
rect 20899 7377 20957 7383
rect 20809 7355 20867 7361
rect 16485 7327 16543 7333
rect 15212 7296 16252 7324
rect 15013 7287 15071 7293
rect 15028 7256 15056 7287
rect 14844 7228 15056 7256
rect 14844 7200 14872 7228
rect 12820 7160 14504 7188
rect 14826 7148 14832 7200
rect 14884 7148 14890 7200
rect 15286 7148 15292 7200
rect 15344 7148 15350 7200
rect 16224 7188 16252 7296
rect 16485 7293 16497 7327
rect 16531 7293 16543 7327
rect 16485 7287 16543 7293
rect 17773 7327 17831 7333
rect 17773 7293 17785 7327
rect 17819 7324 17831 7327
rect 17954 7324 17960 7336
rect 17819 7296 17960 7324
rect 17819 7293 17831 7296
rect 17773 7287 17831 7293
rect 16298 7216 16304 7268
rect 16356 7256 16362 7268
rect 16500 7256 16528 7287
rect 17954 7284 17960 7296
rect 18012 7324 18018 7336
rect 18432 7324 18460 7352
rect 18012 7296 18460 7324
rect 18012 7284 18018 7296
rect 19978 7284 19984 7336
rect 20036 7324 20042 7336
rect 20456 7324 20484 7355
rect 20036 7296 20484 7324
rect 20036 7284 20042 7296
rect 16356 7228 16528 7256
rect 16592 7228 17448 7256
rect 16356 7216 16362 7228
rect 16592 7188 16620 7228
rect 16224 7160 16620 7188
rect 17420 7188 17448 7228
rect 20530 7216 20536 7268
rect 20588 7256 20594 7268
rect 20824 7256 20852 7355
rect 20990 7352 20996 7404
rect 21048 7352 21054 7404
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7361 21143 7395
rect 21192 7392 21220 7500
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 21416 7500 21465 7528
rect 21416 7488 21422 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 21818 7488 21824 7540
rect 21876 7528 21882 7540
rect 21876 7500 22094 7528
rect 21876 7488 21882 7500
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 21192 7364 21281 7392
rect 21085 7355 21143 7361
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 22066 7392 22094 7500
rect 23014 7488 23020 7540
rect 23072 7528 23078 7540
rect 23385 7531 23443 7537
rect 23385 7528 23397 7531
rect 23072 7500 23397 7528
rect 23072 7488 23078 7500
rect 23385 7497 23397 7500
rect 23431 7497 23443 7531
rect 23385 7491 23443 7497
rect 22175 7395 22233 7401
rect 22175 7392 22187 7395
rect 22066 7364 22187 7392
rect 21269 7355 21327 7361
rect 22175 7361 22187 7364
rect 22221 7361 22233 7395
rect 23400 7392 23428 7491
rect 23934 7488 23940 7540
rect 23992 7488 23998 7540
rect 25409 7531 25467 7537
rect 25409 7497 25421 7531
rect 25455 7497 25467 7531
rect 25409 7491 25467 7497
rect 23952 7460 23980 7488
rect 23952 7432 24072 7460
rect 23661 7395 23719 7401
rect 23661 7392 23673 7395
rect 23400 7364 23673 7392
rect 22175 7355 22233 7361
rect 23661 7361 23673 7364
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 21100 7324 21128 7355
rect 23842 7352 23848 7404
rect 23900 7352 23906 7404
rect 24044 7401 24072 7432
rect 23937 7395 23995 7401
rect 23937 7361 23949 7395
rect 23983 7361 23995 7395
rect 23937 7355 23995 7361
rect 24029 7395 24087 7401
rect 24029 7361 24041 7395
rect 24075 7361 24087 7395
rect 24029 7355 24087 7361
rect 25041 7395 25099 7401
rect 25041 7361 25053 7395
rect 25087 7392 25099 7395
rect 25222 7392 25228 7404
rect 25087 7364 25228 7392
rect 25087 7361 25099 7364
rect 25041 7355 25099 7361
rect 21358 7324 21364 7336
rect 20916 7296 21364 7324
rect 20916 7265 20944 7296
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 22097 7327 22155 7333
rect 22097 7293 22109 7327
rect 22143 7293 22155 7327
rect 23860 7324 23888 7352
rect 22097 7287 22155 7293
rect 22296 7296 23888 7324
rect 20588 7228 20852 7256
rect 20901 7259 20959 7265
rect 20588 7216 20594 7228
rect 20901 7225 20913 7259
rect 20947 7225 20959 7259
rect 22112 7256 22140 7287
rect 22186 7256 22192 7268
rect 22112 7228 22192 7256
rect 20901 7219 20959 7225
rect 22186 7216 22192 7228
rect 22244 7216 22250 7268
rect 22296 7188 22324 7296
rect 23658 7216 23664 7268
rect 23716 7256 23722 7268
rect 23952 7256 23980 7355
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 25424 7392 25452 7491
rect 25958 7488 25964 7540
rect 26016 7488 26022 7540
rect 26789 7531 26847 7537
rect 26789 7497 26801 7531
rect 26835 7528 26847 7531
rect 26835 7500 28396 7528
rect 26835 7497 26847 7500
rect 26789 7491 26847 7497
rect 25976 7460 26004 7488
rect 25976 7432 27844 7460
rect 27816 7401 27844 7432
rect 26789 7395 26847 7401
rect 26789 7392 26801 7395
rect 25424 7364 26801 7392
rect 26789 7361 26801 7364
rect 26835 7392 26847 7395
rect 27249 7395 27307 7401
rect 27249 7392 27261 7395
rect 26835 7364 27261 7392
rect 26835 7361 26847 7364
rect 26789 7355 26847 7361
rect 27249 7361 27261 7364
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 27709 7395 27767 7401
rect 27709 7361 27721 7395
rect 27755 7361 27767 7395
rect 27709 7355 27767 7361
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 24305 7327 24363 7333
rect 24305 7293 24317 7327
rect 24351 7324 24363 7327
rect 24949 7327 25007 7333
rect 24949 7324 24961 7327
rect 24351 7296 24961 7324
rect 24351 7293 24363 7296
rect 24305 7287 24363 7293
rect 24949 7293 24961 7296
rect 24995 7293 25007 7327
rect 24949 7287 25007 7293
rect 26510 7284 26516 7336
rect 26568 7324 26574 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26568 7296 26985 7324
rect 26568 7284 26574 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 26973 7287 27031 7293
rect 27062 7284 27068 7336
rect 27120 7284 27126 7336
rect 23716 7228 23980 7256
rect 26697 7259 26755 7265
rect 23716 7216 23722 7228
rect 26697 7225 26709 7259
rect 26743 7256 26755 7259
rect 27080 7256 27108 7284
rect 26743 7228 27108 7256
rect 27433 7259 27491 7265
rect 26743 7225 26755 7228
rect 26697 7219 26755 7225
rect 27433 7225 27445 7259
rect 27479 7256 27491 7259
rect 27724 7256 27752 7355
rect 27982 7352 27988 7404
rect 28040 7352 28046 7404
rect 28368 7401 28396 7500
rect 28077 7395 28135 7401
rect 28077 7361 28089 7395
rect 28123 7361 28135 7395
rect 28077 7355 28135 7361
rect 28353 7395 28411 7401
rect 28353 7361 28365 7395
rect 28399 7361 28411 7395
rect 28353 7355 28411 7361
rect 28537 7395 28595 7401
rect 28537 7361 28549 7395
rect 28583 7361 28595 7395
rect 28537 7355 28595 7361
rect 28092 7324 28120 7355
rect 28166 7324 28172 7336
rect 28092 7296 28172 7324
rect 28166 7284 28172 7296
rect 28224 7324 28230 7336
rect 28445 7327 28503 7333
rect 28445 7324 28457 7327
rect 28224 7296 28457 7324
rect 28224 7284 28230 7296
rect 28445 7293 28457 7296
rect 28491 7293 28503 7327
rect 28445 7287 28503 7293
rect 28552 7256 28580 7355
rect 27479 7228 28580 7256
rect 27479 7225 27491 7228
rect 27433 7219 27491 7225
rect 17420 7160 22324 7188
rect 22370 7148 22376 7200
rect 22428 7148 22434 7200
rect 28258 7148 28264 7200
rect 28316 7148 28322 7200
rect 1104 7098 35248 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 35248 7098
rect 1104 7024 35248 7046
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8938 6984 8944 6996
rect 8352 6956 8944 6984
rect 8352 6944 8358 6956
rect 8938 6944 8944 6956
rect 8996 6944 9002 6996
rect 9263 6987 9321 6993
rect 9263 6984 9275 6987
rect 9048 6956 9275 6984
rect 9048 6916 9076 6956
rect 9263 6953 9275 6956
rect 9309 6984 9321 6987
rect 10226 6984 10232 6996
rect 9309 6956 10232 6984
rect 9309 6953 9321 6956
rect 9263 6947 9321 6953
rect 10226 6944 10232 6956
rect 10284 6944 10290 6996
rect 12452 6956 13584 6984
rect 12452 6928 12480 6956
rect 7208 6888 9076 6916
rect 9401 6919 9459 6925
rect 7208 6792 7236 6888
rect 9401 6885 9413 6919
rect 9447 6885 9459 6919
rect 9401 6879 9459 6885
rect 7282 6808 7288 6860
rect 7340 6848 7346 6860
rect 7837 6851 7895 6857
rect 7837 6848 7849 6851
rect 7340 6820 7849 6848
rect 7340 6808 7346 6820
rect 7837 6817 7849 6820
rect 7883 6817 7895 6851
rect 9122 6848 9128 6860
rect 7837 6811 7895 6817
rect 8588 6820 9128 6848
rect 8588 6792 8616 6820
rect 9122 6808 9128 6820
rect 9180 6848 9186 6860
rect 9416 6848 9444 6879
rect 12434 6876 12440 6928
rect 12492 6876 12498 6928
rect 12710 6876 12716 6928
rect 12768 6916 12774 6928
rect 13078 6916 13084 6928
rect 12768 6888 13084 6916
rect 12768 6876 12774 6888
rect 13078 6876 13084 6888
rect 13136 6876 13142 6928
rect 9180 6820 9444 6848
rect 9493 6851 9551 6857
rect 9180 6808 9186 6820
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9582 6848 9588 6860
rect 9539 6820 9588 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 7190 6740 7196 6792
rect 7248 6740 7254 6792
rect 7558 6740 7564 6792
rect 7616 6740 7622 6792
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 8202 6780 8208 6792
rect 8159 6752 8208 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 8202 6740 8208 6752
rect 8260 6740 8266 6792
rect 8570 6740 8576 6792
rect 8628 6740 8634 6792
rect 8662 6740 8668 6792
rect 8720 6780 8726 6792
rect 9508 6780 9536 6811
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 8720 6752 9536 6780
rect 10413 6783 10471 6789
rect 8720 6740 8726 6752
rect 10413 6749 10425 6783
rect 10459 6780 10471 6783
rect 10594 6780 10600 6792
rect 10459 6752 10600 6780
rect 10459 6749 10471 6752
rect 10413 6743 10471 6749
rect 10594 6740 10600 6752
rect 10652 6740 10658 6792
rect 10686 6740 10692 6792
rect 10744 6740 10750 6792
rect 12618 6740 12624 6792
rect 12676 6740 12682 6792
rect 13078 6740 13084 6792
rect 13136 6780 13142 6792
rect 13173 6783 13231 6789
rect 13173 6780 13185 6783
rect 13136 6752 13185 6780
rect 13136 6740 13142 6752
rect 13173 6749 13185 6752
rect 13219 6749 13231 6783
rect 13556 6780 13584 6956
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 16025 6987 16083 6993
rect 16025 6984 16037 6987
rect 15988 6956 16037 6984
rect 15988 6944 15994 6956
rect 16025 6953 16037 6956
rect 16071 6953 16083 6987
rect 16025 6947 16083 6953
rect 16040 6916 16068 6947
rect 17770 6944 17776 6996
rect 17828 6944 17834 6996
rect 21174 6944 21180 6996
rect 21232 6944 21238 6996
rect 23569 6987 23627 6993
rect 23569 6953 23581 6987
rect 23615 6984 23627 6987
rect 23658 6984 23664 6996
rect 23615 6956 23664 6984
rect 23615 6953 23627 6956
rect 23569 6947 23627 6953
rect 23658 6944 23664 6956
rect 23716 6944 23722 6996
rect 23934 6916 23940 6928
rect 16040 6888 23940 6916
rect 23934 6876 23940 6888
rect 23992 6876 23998 6928
rect 16022 6808 16028 6860
rect 16080 6848 16086 6860
rect 16080 6820 16160 6848
rect 16080 6808 16086 6820
rect 13556 6752 14136 6780
rect 13173 6743 13231 6749
rect 7576 6712 7604 6740
rect 8021 6715 8079 6721
rect 8021 6712 8033 6715
rect 7576 6684 8033 6712
rect 8021 6681 8033 6684
rect 8067 6681 8079 6715
rect 8021 6675 8079 6681
rect 9030 6672 9036 6724
rect 9088 6712 9094 6724
rect 9125 6715 9183 6721
rect 9125 6712 9137 6715
rect 9088 6684 9137 6712
rect 9088 6672 9094 6684
rect 9125 6681 9137 6684
rect 9171 6712 9183 6715
rect 10318 6712 10324 6724
rect 9171 6684 10324 6712
rect 9171 6681 9183 6684
rect 9125 6675 9183 6681
rect 10318 6672 10324 6684
rect 10376 6672 10382 6724
rect 11606 6712 11612 6724
rect 11546 6684 11612 6712
rect 11606 6672 11612 6684
rect 11664 6672 11670 6724
rect 14108 6712 14136 6752
rect 14182 6740 14188 6792
rect 14240 6740 14246 6792
rect 16132 6789 16160 6820
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 18509 6851 18567 6857
rect 18509 6848 18521 6851
rect 18472 6820 18521 6848
rect 18472 6808 18478 6820
rect 18509 6817 18521 6820
rect 18555 6817 18567 6851
rect 18509 6811 18567 6817
rect 18969 6851 19027 6857
rect 18969 6817 18981 6851
rect 19015 6848 19027 6851
rect 19334 6848 19340 6860
rect 19015 6820 19340 6848
rect 19015 6817 19027 6820
rect 18969 6811 19027 6817
rect 19334 6808 19340 6820
rect 19392 6848 19398 6860
rect 19392 6820 19656 6848
rect 19392 6808 19398 6820
rect 14553 6783 14611 6789
rect 14553 6749 14565 6783
rect 14599 6749 14611 6783
rect 14553 6743 14611 6749
rect 16117 6783 16175 6789
rect 16117 6749 16129 6783
rect 16163 6749 16175 6783
rect 16117 6743 16175 6749
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16298 6780 16304 6792
rect 16255 6752 16304 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 14568 6712 14596 6743
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 17497 6783 17555 6789
rect 17497 6749 17509 6783
rect 17543 6780 17555 6783
rect 17586 6780 17592 6792
rect 17543 6752 17592 6780
rect 17543 6749 17555 6752
rect 17497 6743 17555 6749
rect 16408 6712 16436 6743
rect 17586 6740 17592 6752
rect 17644 6740 17650 6792
rect 17773 6783 17831 6789
rect 17773 6749 17785 6783
rect 17819 6749 17831 6783
rect 17773 6743 17831 6749
rect 13570 6684 14044 6712
rect 14108 6684 14596 6712
rect 16132 6684 16436 6712
rect 9769 6647 9827 6653
rect 9769 6613 9781 6647
rect 9815 6644 9827 6647
rect 10502 6644 10508 6656
rect 9815 6616 10508 6644
rect 9815 6613 9827 6616
rect 9769 6607 9827 6613
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 10686 6604 10692 6656
rect 10744 6644 10750 6656
rect 12158 6644 12164 6656
rect 10744 6616 12164 6644
rect 10744 6604 10750 6616
rect 12158 6604 12164 6616
rect 12216 6644 12222 6656
rect 13906 6644 13912 6656
rect 12216 6616 13912 6644
rect 12216 6604 12222 6616
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14016 6644 14044 6684
rect 16132 6656 16160 6684
rect 16482 6672 16488 6724
rect 16540 6712 16546 6724
rect 17678 6712 17684 6724
rect 16540 6684 17684 6712
rect 16540 6672 16546 6684
rect 17678 6672 17684 6684
rect 17736 6672 17742 6724
rect 17788 6656 17816 6743
rect 18322 6740 18328 6792
rect 18380 6780 18386 6792
rect 18601 6783 18659 6789
rect 18601 6780 18613 6783
rect 18380 6752 18613 6780
rect 18380 6740 18386 6752
rect 18601 6749 18613 6752
rect 18647 6749 18659 6783
rect 18601 6743 18659 6749
rect 19426 6740 19432 6792
rect 19484 6740 19490 6792
rect 19628 6789 19656 6820
rect 21082 6808 21088 6860
rect 21140 6808 21146 6860
rect 28166 6808 28172 6860
rect 28224 6808 28230 6860
rect 28442 6808 28448 6860
rect 28500 6808 28506 6860
rect 19613 6783 19671 6789
rect 19613 6749 19625 6783
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 19797 6783 19855 6789
rect 19797 6749 19809 6783
rect 19843 6780 19855 6783
rect 20162 6780 20168 6792
rect 19843 6752 20168 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 20162 6740 20168 6752
rect 20220 6740 20226 6792
rect 20346 6740 20352 6792
rect 20404 6740 20410 6792
rect 20806 6740 20812 6792
rect 20864 6740 20870 6792
rect 21100 6780 21128 6808
rect 21269 6783 21327 6789
rect 21269 6780 21281 6783
rect 21100 6752 21281 6780
rect 21269 6749 21281 6752
rect 21315 6749 21327 6783
rect 21269 6743 21327 6749
rect 21358 6740 21364 6792
rect 21416 6740 21422 6792
rect 27982 6740 27988 6792
rect 28040 6780 28046 6792
rect 28077 6783 28135 6789
rect 28077 6780 28089 6783
rect 28040 6752 28089 6780
rect 28040 6740 28046 6752
rect 28077 6749 28089 6752
rect 28123 6749 28135 6783
rect 28077 6743 28135 6749
rect 20824 6712 20852 6740
rect 21085 6715 21143 6721
rect 21085 6712 21097 6715
rect 20824 6684 21097 6712
rect 21085 6681 21097 6684
rect 21131 6681 21143 6715
rect 21085 6675 21143 6681
rect 14458 6644 14464 6656
rect 14016 6616 14464 6644
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 16114 6604 16120 6656
rect 16172 6604 16178 6656
rect 16574 6604 16580 6656
rect 16632 6604 16638 6656
rect 17770 6604 17776 6656
rect 17828 6604 17834 6656
rect 19978 6604 19984 6656
rect 20036 6604 20042 6656
rect 1104 6554 35236 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 35236 6554
rect 1104 6480 35236 6502
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 9824 6412 12940 6440
rect 9824 6400 9830 6412
rect 9950 6372 9956 6384
rect 8970 6344 9956 6372
rect 9950 6332 9956 6344
rect 10008 6372 10014 6384
rect 10686 6372 10692 6384
rect 10008 6344 10692 6372
rect 10008 6332 10014 6344
rect 10686 6332 10692 6344
rect 10744 6332 10750 6384
rect 11330 6332 11336 6384
rect 11388 6332 11394 6384
rect 12802 6332 12808 6384
rect 12860 6332 12866 6384
rect 12912 6372 12940 6412
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 14826 6440 14832 6452
rect 13964 6412 14832 6440
rect 13964 6400 13970 6412
rect 14826 6400 14832 6412
rect 14884 6400 14890 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6440 14979 6443
rect 15102 6440 15108 6452
rect 14967 6412 15108 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 15286 6400 15292 6452
rect 15344 6400 15350 6452
rect 15562 6400 15568 6452
rect 15620 6400 15626 6452
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 16317 6443 16375 6449
rect 16317 6440 16329 6443
rect 16080 6412 16329 6440
rect 16080 6400 16086 6412
rect 16317 6409 16329 6412
rect 16363 6409 16375 6443
rect 16317 6403 16375 6409
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6409 17279 6443
rect 17221 6403 17279 6409
rect 17865 6443 17923 6449
rect 17865 6409 17877 6443
rect 17911 6440 17923 6443
rect 18322 6440 18328 6452
rect 17911 6412 18328 6440
rect 17911 6409 17923 6412
rect 17865 6403 17923 6409
rect 12912 6344 13860 6372
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 8478 6264 8484 6316
rect 8536 6304 8542 6316
rect 8573 6307 8631 6313
rect 8573 6304 8585 6307
rect 8536 6276 8585 6304
rect 8536 6264 8542 6276
rect 8573 6273 8585 6276
rect 8619 6273 8631 6307
rect 8573 6267 8631 6273
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 10226 6264 10232 6316
rect 10284 6264 10290 6316
rect 12066 6264 12072 6316
rect 12124 6264 12130 6316
rect 12820 6304 12848 6332
rect 13265 6307 13323 6313
rect 13265 6304 13277 6307
rect 12820 6276 13277 6304
rect 11606 6196 11612 6248
rect 11664 6196 11670 6248
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 12250 6236 12256 6248
rect 11756 6208 12256 6236
rect 11756 6196 11762 6208
rect 12250 6196 12256 6208
rect 12308 6236 12314 6248
rect 12805 6239 12863 6245
rect 12805 6236 12817 6239
rect 12308 6208 12817 6236
rect 12308 6196 12314 6208
rect 12805 6205 12817 6208
rect 12851 6205 12863 6239
rect 12805 6199 12863 6205
rect 12526 6128 12532 6180
rect 12584 6128 12590 6180
rect 11054 6060 11060 6112
rect 11112 6100 11118 6112
rect 12912 6100 12940 6276
rect 13265 6273 13277 6276
rect 13311 6273 13323 6307
rect 13265 6267 13323 6273
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 13832 6304 13860 6344
rect 13998 6332 14004 6384
rect 14056 6332 14062 6384
rect 14734 6332 14740 6384
rect 14792 6332 14798 6384
rect 14752 6304 14780 6332
rect 15304 6313 15332 6400
rect 13832 6276 14780 6304
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15289 6267 15347 6273
rect 15473 6307 15531 6313
rect 15473 6273 15485 6307
rect 15519 6304 15531 6307
rect 15580 6304 15608 6400
rect 16117 6375 16175 6381
rect 16117 6341 16129 6375
rect 16163 6372 16175 6375
rect 16206 6372 16212 6384
rect 16163 6344 16212 6372
rect 16163 6341 16175 6344
rect 16117 6335 16175 6341
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 16482 6304 16488 6316
rect 15519 6276 15608 6304
rect 15948 6276 16488 6304
rect 15519 6273 15531 6276
rect 15473 6267 15531 6273
rect 12986 6196 12992 6248
rect 13044 6196 13050 6248
rect 15948 6180 15976 6276
rect 16482 6264 16488 6276
rect 16540 6264 16546 6316
rect 17236 6304 17264 6403
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 19334 6400 19340 6452
rect 19392 6400 19398 6452
rect 19521 6443 19579 6449
rect 19521 6409 19533 6443
rect 19567 6440 19579 6443
rect 20346 6440 20352 6452
rect 19567 6412 20352 6440
rect 19567 6409 19579 6412
rect 19521 6403 19579 6409
rect 20346 6400 20352 6412
rect 20404 6400 20410 6452
rect 17402 6332 17408 6384
rect 17460 6372 17466 6384
rect 17681 6375 17739 6381
rect 17681 6372 17693 6375
rect 17460 6344 17693 6372
rect 17460 6332 17466 6344
rect 17681 6341 17693 6344
rect 17727 6372 17739 6375
rect 19352 6372 19380 6400
rect 17727 6344 18184 6372
rect 19352 6344 19564 6372
rect 17727 6341 17739 6344
rect 17681 6335 17739 6341
rect 17770 6304 17776 6316
rect 17236 6276 17776 6304
rect 17770 6264 17776 6276
rect 17828 6304 17834 6316
rect 18156 6313 18184 6344
rect 17957 6307 18015 6313
rect 17957 6304 17969 6307
rect 17828 6276 17969 6304
rect 17828 6264 17834 6276
rect 17957 6273 17969 6276
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6273 18199 6307
rect 18141 6267 18199 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 16761 6239 16819 6245
rect 16761 6236 16773 6239
rect 16500 6208 16773 6236
rect 14550 6128 14556 6180
rect 14608 6168 14614 6180
rect 14826 6168 14832 6180
rect 14608 6140 14832 6168
rect 14608 6128 14614 6140
rect 14826 6128 14832 6140
rect 14884 6128 14890 6180
rect 15105 6171 15163 6177
rect 15105 6137 15117 6171
rect 15151 6168 15163 6171
rect 15930 6168 15936 6180
rect 15151 6140 15936 6168
rect 15151 6137 15163 6140
rect 15105 6131 15163 6137
rect 15930 6128 15936 6140
rect 15988 6128 15994 6180
rect 16500 6177 16528 6208
rect 16761 6205 16773 6208
rect 16807 6236 16819 6239
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16807 6208 17325 6236
rect 16807 6205 16819 6208
rect 16761 6199 16819 6205
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 17678 6196 17684 6248
rect 17736 6236 17742 6248
rect 18248 6236 18276 6267
rect 19426 6264 19432 6316
rect 19484 6264 19490 6316
rect 19536 6304 19564 6344
rect 19613 6307 19671 6313
rect 19613 6304 19625 6307
rect 19536 6276 19625 6304
rect 19613 6273 19625 6276
rect 19659 6273 19671 6307
rect 19613 6267 19671 6273
rect 17736 6208 18276 6236
rect 17736 6196 17742 6208
rect 16485 6171 16543 6177
rect 16485 6137 16497 6171
rect 16531 6137 16543 6171
rect 16485 6131 16543 6137
rect 16574 6128 16580 6180
rect 16632 6168 16638 6180
rect 17037 6171 17095 6177
rect 17037 6168 17049 6171
rect 16632 6140 17049 6168
rect 16632 6128 16638 6140
rect 17037 6137 17049 6140
rect 17083 6168 17095 6171
rect 17083 6140 17724 6168
rect 17083 6137 17095 6140
rect 17037 6131 17095 6137
rect 11112 6072 12940 6100
rect 15381 6103 15439 6109
rect 11112 6060 11118 6072
rect 15381 6069 15393 6103
rect 15427 6100 15439 6103
rect 16206 6100 16212 6112
rect 15427 6072 16212 6100
rect 15427 6069 15439 6072
rect 15381 6063 15439 6069
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16301 6103 16359 6109
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 16390 6100 16396 6112
rect 16347 6072 16396 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 17696 6109 17724 6140
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18325 6171 18383 6177
rect 18325 6168 18337 6171
rect 18012 6140 18337 6168
rect 18012 6128 18018 6140
rect 18325 6137 18337 6140
rect 18371 6137 18383 6171
rect 18325 6131 18383 6137
rect 17681 6103 17739 6109
rect 17681 6069 17693 6103
rect 17727 6069 17739 6103
rect 17681 6063 17739 6069
rect 18138 6060 18144 6112
rect 18196 6060 18202 6112
rect 1104 6010 35248 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 35248 6010
rect 1104 5936 35248 5958
rect 8478 5856 8484 5908
rect 8536 5856 8542 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9079 5899 9137 5905
rect 9079 5896 9091 5899
rect 8812 5868 9091 5896
rect 8812 5856 8818 5868
rect 9079 5865 9091 5868
rect 9125 5865 9137 5899
rect 9079 5859 9137 5865
rect 9674 5856 9680 5908
rect 9732 5896 9738 5908
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 9732 5868 10149 5896
rect 9732 5856 9738 5868
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 10137 5859 10195 5865
rect 10410 5856 10416 5908
rect 10468 5896 10474 5908
rect 10594 5896 10600 5908
rect 10468 5868 10600 5896
rect 10468 5856 10474 5868
rect 10594 5856 10600 5868
rect 10652 5896 10658 5908
rect 10781 5899 10839 5905
rect 10781 5896 10793 5899
rect 10652 5868 10793 5896
rect 10652 5856 10658 5868
rect 10781 5865 10793 5868
rect 10827 5865 10839 5899
rect 10781 5859 10839 5865
rect 11054 5856 11060 5908
rect 11112 5856 11118 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11606 5896 11612 5908
rect 11287 5868 11612 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 13173 5899 13231 5905
rect 13173 5865 13185 5899
rect 13219 5896 13231 5899
rect 14182 5896 14188 5908
rect 13219 5868 14188 5896
rect 13219 5865 13231 5868
rect 13173 5859 13231 5865
rect 14182 5856 14188 5868
rect 14240 5856 14246 5908
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 14918 5896 14924 5908
rect 14875 5868 14924 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15289 5899 15347 5905
rect 15289 5865 15301 5899
rect 15335 5896 15347 5899
rect 15378 5896 15384 5908
rect 15335 5868 15384 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 17402 5856 17408 5908
rect 17460 5856 17466 5908
rect 17954 5856 17960 5908
rect 18012 5856 18018 5908
rect 18138 5856 18144 5908
rect 18196 5856 18202 5908
rect 21266 5896 21272 5908
rect 20548 5868 21272 5896
rect 8496 5828 8524 5856
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 8496 5800 9229 5828
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 8496 5760 8524 5800
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9217 5791 9275 5797
rect 9585 5831 9643 5837
rect 9585 5797 9597 5831
rect 9631 5828 9643 5831
rect 11072 5828 11100 5856
rect 12802 5828 12808 5840
rect 9631 5800 11100 5828
rect 12406 5800 12808 5828
rect 9631 5797 9643 5800
rect 9585 5791 9643 5797
rect 7239 5732 8524 5760
rect 9309 5763 9367 5769
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 9309 5729 9321 5763
rect 9355 5760 9367 5763
rect 9766 5760 9772 5772
rect 9355 5732 9772 5760
rect 9355 5729 9367 5732
rect 9309 5723 9367 5729
rect 5166 5652 5172 5704
rect 5224 5652 5230 5704
rect 6546 5652 6552 5704
rect 6604 5652 6610 5704
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 9324 5692 9352 5723
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 10873 5763 10931 5769
rect 10873 5760 10885 5763
rect 10244 5732 10885 5760
rect 10244 5704 10272 5732
rect 10873 5729 10885 5732
rect 10919 5729 10931 5763
rect 12406 5760 12434 5800
rect 12802 5788 12808 5800
rect 12860 5788 12866 5840
rect 10873 5723 10931 5729
rect 12268 5732 12434 5760
rect 12529 5763 12587 5769
rect 8260 5664 9352 5692
rect 8260 5652 8266 5664
rect 10226 5652 10232 5704
rect 10284 5652 10290 5704
rect 10318 5652 10324 5704
rect 10376 5652 10382 5704
rect 10410 5652 10416 5704
rect 10468 5652 10474 5704
rect 10502 5652 10508 5704
rect 10560 5652 10566 5704
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5661 10655 5695
rect 10597 5655 10655 5661
rect 4798 5584 4804 5636
rect 4856 5624 4862 5636
rect 5445 5627 5503 5633
rect 5445 5624 5457 5627
rect 4856 5596 5457 5624
rect 4856 5584 4862 5596
rect 5445 5593 5457 5596
rect 5491 5593 5503 5627
rect 5445 5587 5503 5593
rect 8938 5584 8944 5636
rect 8996 5624 9002 5636
rect 9398 5624 9404 5636
rect 8996 5596 9404 5624
rect 8996 5584 9002 5596
rect 9398 5584 9404 5596
rect 9456 5584 9462 5636
rect 10336 5556 10364 5652
rect 10612 5624 10640 5655
rect 10686 5652 10692 5704
rect 10744 5692 10750 5704
rect 10781 5695 10839 5701
rect 10781 5692 10793 5695
rect 10744 5664 10793 5692
rect 10744 5652 10750 5664
rect 10781 5661 10793 5664
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 12268 5701 12296 5732
rect 12529 5729 12541 5763
rect 12575 5760 12587 5763
rect 12618 5760 12624 5772
rect 12575 5732 12624 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 14936 5760 14964 5856
rect 14936 5732 15240 5760
rect 15212 5704 15240 5732
rect 11057 5695 11115 5701
rect 11057 5661 11069 5695
rect 11103 5661 11115 5695
rect 11057 5655 11115 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5661 12311 5695
rect 12253 5655 12311 5661
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5692 12495 5695
rect 12713 5695 12771 5701
rect 12713 5692 12725 5695
rect 12483 5664 12725 5692
rect 12483 5661 12495 5664
rect 12437 5655 12495 5661
rect 12713 5661 12725 5664
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 10980 5624 11008 5652
rect 10612 5596 11008 5624
rect 10778 5556 10784 5568
rect 10336 5528 10784 5556
rect 10778 5516 10784 5528
rect 10836 5556 10842 5568
rect 11072 5556 11100 5655
rect 12728 5624 12756 5655
rect 12894 5652 12900 5704
rect 12952 5652 12958 5704
rect 12989 5695 13047 5701
rect 12989 5661 13001 5695
rect 13035 5692 13047 5695
rect 13446 5692 13452 5704
rect 13035 5664 13452 5692
rect 13035 5661 13047 5664
rect 12989 5655 13047 5661
rect 13446 5652 13452 5664
rect 13504 5652 13510 5704
rect 14734 5652 14740 5704
rect 14792 5652 14798 5704
rect 14826 5652 14832 5704
rect 14884 5692 14890 5704
rect 14921 5695 14979 5701
rect 14921 5692 14933 5695
rect 14884 5664 14933 5692
rect 14884 5652 14890 5664
rect 14921 5661 14933 5664
rect 14967 5661 14979 5695
rect 14921 5655 14979 5661
rect 15194 5652 15200 5704
rect 15252 5652 15258 5704
rect 15562 5652 15568 5704
rect 15620 5692 15626 5704
rect 17313 5695 17371 5701
rect 17313 5692 17325 5695
rect 15620 5664 17325 5692
rect 15620 5652 15626 5664
rect 17313 5661 17325 5664
rect 17359 5661 17371 5695
rect 17313 5655 17371 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5692 17555 5695
rect 17972 5692 18000 5856
rect 18156 5701 18184 5856
rect 20349 5763 20407 5769
rect 20349 5760 20361 5763
rect 19720 5732 20361 5760
rect 17543 5664 18000 5692
rect 18141 5695 18199 5701
rect 17543 5661 17555 5664
rect 17497 5655 17555 5661
rect 18141 5661 18153 5695
rect 18187 5661 18199 5695
rect 18141 5655 18199 5661
rect 18322 5652 18328 5704
rect 18380 5652 18386 5704
rect 19720 5701 19748 5732
rect 20349 5729 20361 5732
rect 20395 5760 20407 5763
rect 20438 5760 20444 5772
rect 20395 5732 20444 5760
rect 20395 5729 20407 5732
rect 20349 5723 20407 5729
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 20548 5769 20576 5868
rect 21266 5856 21272 5868
rect 21324 5856 21330 5908
rect 22925 5899 22983 5905
rect 22925 5865 22937 5899
rect 22971 5896 22983 5899
rect 23474 5896 23480 5908
rect 22971 5868 23480 5896
rect 22971 5865 22983 5868
rect 22925 5859 22983 5865
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 23750 5856 23756 5908
rect 23808 5856 23814 5908
rect 27430 5856 27436 5908
rect 27488 5856 27494 5908
rect 23109 5831 23167 5837
rect 23109 5828 23121 5831
rect 22480 5800 23121 5828
rect 22480 5772 22508 5800
rect 23109 5797 23121 5800
rect 23155 5797 23167 5831
rect 23109 5791 23167 5797
rect 26697 5831 26755 5837
rect 26697 5797 26709 5831
rect 26743 5828 26755 5831
rect 27154 5828 27160 5840
rect 26743 5800 27160 5828
rect 26743 5797 26755 5800
rect 26697 5791 26755 5797
rect 27154 5788 27160 5800
rect 27212 5788 27218 5840
rect 20533 5763 20591 5769
rect 20533 5729 20545 5763
rect 20579 5729 20591 5763
rect 20533 5723 20591 5729
rect 20993 5763 21051 5769
rect 20993 5729 21005 5763
rect 21039 5760 21051 5763
rect 21358 5760 21364 5772
rect 21039 5732 21364 5760
rect 21039 5729 21051 5732
rect 20993 5723 21051 5729
rect 21358 5720 21364 5732
rect 21416 5720 21422 5772
rect 22462 5720 22468 5772
rect 22520 5720 22526 5772
rect 23014 5720 23020 5772
rect 23072 5760 23078 5772
rect 23477 5763 23535 5769
rect 23072 5732 23428 5760
rect 23072 5720 23078 5732
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5692 19947 5695
rect 19978 5692 19984 5704
rect 19935 5664 19984 5692
rect 19935 5661 19947 5664
rect 19889 5655 19947 5661
rect 19978 5652 19984 5664
rect 20036 5692 20042 5704
rect 20165 5695 20223 5701
rect 20165 5692 20177 5695
rect 20036 5664 20177 5692
rect 20036 5652 20042 5664
rect 20165 5661 20177 5664
rect 20211 5661 20223 5695
rect 20165 5655 20223 5661
rect 20625 5695 20683 5701
rect 20625 5661 20637 5695
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 22557 5695 22615 5701
rect 22557 5661 22569 5695
rect 22603 5661 22615 5695
rect 22557 5655 22615 5661
rect 23293 5695 23351 5701
rect 23293 5661 23305 5695
rect 23339 5661 23351 5695
rect 23400 5692 23428 5732
rect 23477 5729 23489 5763
rect 23523 5760 23535 5763
rect 23566 5760 23572 5772
rect 23523 5732 23572 5760
rect 23523 5729 23535 5732
rect 23477 5723 23535 5729
rect 23566 5720 23572 5732
rect 23624 5720 23630 5772
rect 27341 5763 27399 5769
rect 24504 5732 26464 5760
rect 24504 5701 24532 5732
rect 26436 5704 26464 5732
rect 26712 5732 27292 5760
rect 23845 5695 23903 5701
rect 23845 5692 23857 5695
rect 23400 5664 23857 5692
rect 23293 5655 23351 5661
rect 23845 5661 23857 5664
rect 23891 5692 23903 5695
rect 24489 5695 24547 5701
rect 24489 5692 24501 5695
rect 23891 5664 24501 5692
rect 23891 5661 23903 5664
rect 23845 5655 23903 5661
rect 24489 5661 24501 5664
rect 24535 5661 24547 5695
rect 24489 5655 24547 5661
rect 19797 5627 19855 5633
rect 12728 5596 12848 5624
rect 12820 5568 12848 5596
rect 19797 5593 19809 5627
rect 19843 5624 19855 5627
rect 20070 5624 20076 5636
rect 19843 5596 20076 5624
rect 19843 5593 19855 5596
rect 19797 5587 19855 5593
rect 20070 5584 20076 5596
rect 20128 5624 20134 5636
rect 20640 5624 20668 5655
rect 20128 5596 20668 5624
rect 22572 5624 22600 5655
rect 22922 5624 22928 5636
rect 22572 5596 22928 5624
rect 20128 5584 20134 5596
rect 22922 5584 22928 5596
rect 22980 5624 22986 5636
rect 23308 5624 23336 5655
rect 24578 5652 24584 5704
rect 24636 5692 24642 5704
rect 24673 5695 24731 5701
rect 24673 5692 24685 5695
rect 24636 5664 24685 5692
rect 24636 5652 24642 5664
rect 24673 5661 24685 5664
rect 24719 5661 24731 5695
rect 24673 5655 24731 5661
rect 24949 5695 25007 5701
rect 24949 5661 24961 5695
rect 24995 5661 25007 5695
rect 24949 5655 25007 5661
rect 24964 5624 24992 5655
rect 26418 5652 26424 5704
rect 26476 5692 26482 5704
rect 26712 5701 26740 5732
rect 26513 5695 26571 5701
rect 26513 5692 26525 5695
rect 26476 5664 26525 5692
rect 26476 5652 26482 5664
rect 26513 5661 26525 5664
rect 26559 5661 26571 5695
rect 26513 5655 26571 5661
rect 26697 5695 26755 5701
rect 26697 5661 26709 5695
rect 26743 5661 26755 5695
rect 26697 5655 26755 5661
rect 27065 5695 27123 5701
rect 27065 5661 27077 5695
rect 27111 5661 27123 5695
rect 27264 5692 27292 5732
rect 27341 5729 27353 5763
rect 27387 5760 27399 5763
rect 27448 5760 27476 5856
rect 27387 5732 27476 5760
rect 27387 5729 27399 5732
rect 27341 5723 27399 5729
rect 27522 5692 27528 5704
rect 27264 5664 27528 5692
rect 27065 5655 27123 5661
rect 22980 5596 23336 5624
rect 24136 5596 24992 5624
rect 22980 5584 22986 5596
rect 24136 5568 24164 5596
rect 10836 5528 11100 5556
rect 10836 5516 10842 5528
rect 12802 5516 12808 5568
rect 12860 5516 12866 5568
rect 18230 5516 18236 5568
rect 18288 5516 18294 5568
rect 19978 5516 19984 5568
rect 20036 5516 20042 5568
rect 23569 5559 23627 5565
rect 23569 5525 23581 5559
rect 23615 5556 23627 5559
rect 24118 5556 24124 5568
rect 23615 5528 24124 5556
rect 23615 5525 23627 5528
rect 23569 5519 23627 5525
rect 24118 5516 24124 5528
rect 24176 5516 24182 5568
rect 25130 5516 25136 5568
rect 25188 5516 25194 5568
rect 27080 5556 27108 5655
rect 27522 5652 27528 5664
rect 27580 5692 27586 5704
rect 28074 5692 28080 5704
rect 27580 5664 28080 5692
rect 27580 5652 27586 5664
rect 28074 5652 28080 5664
rect 28132 5652 28138 5704
rect 28169 5695 28227 5701
rect 28169 5661 28181 5695
rect 28215 5661 28227 5695
rect 28169 5655 28227 5661
rect 28184 5568 28212 5655
rect 28258 5652 28264 5704
rect 28316 5652 28322 5704
rect 28445 5695 28503 5701
rect 28445 5661 28457 5695
rect 28491 5661 28503 5695
rect 28445 5655 28503 5661
rect 28537 5695 28595 5701
rect 28537 5661 28549 5695
rect 28583 5692 28595 5695
rect 28902 5692 28908 5704
rect 28583 5664 28908 5692
rect 28583 5661 28595 5664
rect 28537 5655 28595 5661
rect 28460 5624 28488 5655
rect 28902 5652 28908 5664
rect 28960 5652 28966 5704
rect 28460 5596 28580 5624
rect 28552 5568 28580 5596
rect 27246 5556 27252 5568
rect 27080 5528 27252 5556
rect 27246 5516 27252 5528
rect 27304 5516 27310 5568
rect 27341 5559 27399 5565
rect 27341 5525 27353 5559
rect 27387 5556 27399 5559
rect 27706 5556 27712 5568
rect 27387 5528 27712 5556
rect 27387 5525 27399 5528
rect 27341 5519 27399 5525
rect 27706 5516 27712 5528
rect 27764 5516 27770 5568
rect 28166 5516 28172 5568
rect 28224 5516 28230 5568
rect 28534 5516 28540 5568
rect 28592 5516 28598 5568
rect 28721 5559 28779 5565
rect 28721 5525 28733 5559
rect 28767 5556 28779 5559
rect 29546 5556 29552 5568
rect 28767 5528 29552 5556
rect 28767 5525 28779 5528
rect 28721 5519 28779 5525
rect 29546 5516 29552 5528
rect 29604 5516 29610 5568
rect 1104 5466 35236 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 35236 5466
rect 1104 5392 35236 5414
rect 12066 5312 12072 5364
rect 12124 5312 12130 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15381 5355 15439 5361
rect 15381 5352 15393 5355
rect 15252 5324 15393 5352
rect 15252 5312 15258 5324
rect 15381 5321 15393 5324
rect 15427 5321 15439 5355
rect 15381 5315 15439 5321
rect 15470 5312 15476 5364
rect 15528 5312 15534 5364
rect 22922 5312 22928 5364
rect 22980 5312 22986 5364
rect 26050 5312 26056 5364
rect 26108 5312 26114 5364
rect 26878 5312 26884 5364
rect 26936 5352 26942 5364
rect 26973 5355 27031 5361
rect 26973 5352 26985 5355
rect 26936 5324 26985 5352
rect 26936 5312 26942 5324
rect 26973 5321 26985 5324
rect 27019 5321 27031 5355
rect 26973 5315 27031 5321
rect 27430 5312 27436 5364
rect 27488 5352 27494 5364
rect 27488 5324 28028 5352
rect 27488 5312 27494 5324
rect 8481 5287 8539 5293
rect 8481 5253 8493 5287
rect 8527 5284 8539 5287
rect 8754 5284 8760 5296
rect 8527 5256 8760 5284
rect 8527 5253 8539 5256
rect 8481 5247 8539 5253
rect 8754 5244 8760 5256
rect 8812 5244 8818 5296
rect 8294 5216 8300 5228
rect 7866 5188 8300 5216
rect 8294 5176 8300 5188
rect 8352 5176 8358 5228
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11609 5219 11667 5225
rect 11609 5216 11621 5219
rect 11204 5188 11621 5216
rect 11204 5176 11210 5188
rect 11609 5185 11621 5188
rect 11655 5216 11667 5219
rect 11698 5216 11704 5228
rect 11655 5188 11704 5216
rect 11655 5185 11667 5188
rect 11609 5179 11667 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 12084 5216 12112 5312
rect 12802 5244 12808 5296
rect 12860 5284 12866 5296
rect 15488 5284 15516 5312
rect 15749 5287 15807 5293
rect 12860 5256 13768 5284
rect 12860 5244 12866 5256
rect 13740 5228 13768 5256
rect 15488 5256 15700 5284
rect 12342 5216 12348 5228
rect 11808 5188 12204 5216
rect 12303 5188 12348 5216
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 6420 5120 6469 5148
rect 6420 5108 6426 5120
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6457 5111 6515 5117
rect 6730 5108 6736 5160
rect 6788 5108 6794 5160
rect 11517 5151 11575 5157
rect 11517 5117 11529 5151
rect 11563 5148 11575 5151
rect 11808 5148 11836 5188
rect 11563 5120 11836 5148
rect 12069 5151 12127 5157
rect 11563 5117 11575 5120
rect 11517 5111 11575 5117
rect 12069 5117 12081 5151
rect 12115 5117 12127 5151
rect 12176 5148 12204 5188
rect 12342 5176 12348 5188
rect 12400 5216 12406 5228
rect 13538 5216 13544 5228
rect 12400 5188 13544 5216
rect 12400 5176 12406 5188
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 14645 5219 14703 5225
rect 14645 5185 14657 5219
rect 14691 5216 14703 5219
rect 15289 5219 15347 5225
rect 14691 5188 14780 5216
rect 14691 5185 14703 5188
rect 14645 5179 14703 5185
rect 12253 5151 12311 5157
rect 12253 5148 12265 5151
rect 12176 5120 12265 5148
rect 12069 5111 12127 5117
rect 12253 5117 12265 5120
rect 12299 5117 12311 5151
rect 12253 5111 12311 5117
rect 10962 5040 10968 5092
rect 11020 5080 11026 5092
rect 12084 5080 12112 5111
rect 14752 5080 14780 5188
rect 15289 5185 15301 5219
rect 15335 5216 15347 5219
rect 15488 5216 15516 5256
rect 15335 5188 15516 5216
rect 15565 5219 15623 5225
rect 15335 5185 15347 5188
rect 15289 5179 15347 5185
rect 15565 5185 15577 5219
rect 15611 5185 15623 5219
rect 15672 5216 15700 5256
rect 15749 5253 15761 5287
rect 15795 5284 15807 5287
rect 16574 5284 16580 5296
rect 15795 5256 16580 5284
rect 15795 5253 15807 5256
rect 15749 5247 15807 5253
rect 16574 5244 16580 5256
rect 16632 5284 16638 5296
rect 16632 5256 16988 5284
rect 16632 5244 16638 5256
rect 15841 5219 15899 5225
rect 15841 5216 15853 5219
rect 15672 5188 15853 5216
rect 15565 5179 15623 5185
rect 15841 5185 15853 5188
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15580 5148 15608 5179
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 16025 5219 16083 5225
rect 16025 5216 16037 5219
rect 15988 5188 16037 5216
rect 15988 5176 15994 5188
rect 16025 5185 16037 5188
rect 16071 5185 16083 5219
rect 16025 5179 16083 5185
rect 16206 5176 16212 5228
rect 16264 5176 16270 5228
rect 16298 5176 16304 5228
rect 16356 5176 16362 5228
rect 16960 5225 16988 5256
rect 22296 5256 23060 5284
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5216 16543 5219
rect 16761 5219 16819 5225
rect 16761 5216 16773 5219
rect 16531 5188 16773 5216
rect 16531 5185 16543 5188
rect 16485 5179 16543 5185
rect 16761 5185 16773 5188
rect 16807 5185 16819 5219
rect 16761 5179 16819 5185
rect 16945 5219 17003 5225
rect 16945 5185 16957 5219
rect 16991 5185 17003 5219
rect 16945 5179 17003 5185
rect 16224 5148 16252 5176
rect 16500 5148 16528 5179
rect 19978 5176 19984 5228
rect 20036 5176 20042 5228
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 22296 5225 22324 5256
rect 23032 5228 23060 5256
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 20128 5188 20177 5216
rect 20128 5176 20134 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 21453 5219 21511 5225
rect 21453 5216 21465 5219
rect 20165 5179 20223 5185
rect 20272 5188 21465 5216
rect 15243 5120 15700 5148
rect 16224 5120 16528 5148
rect 16669 5151 16727 5157
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 11020 5052 14780 5080
rect 15672 5080 15700 5120
rect 16669 5117 16681 5151
rect 16715 5148 16727 5151
rect 20272 5148 20300 5188
rect 21453 5185 21465 5188
rect 21499 5216 21511 5219
rect 22281 5219 22339 5225
rect 22281 5216 22293 5219
rect 21499 5188 22293 5216
rect 21499 5185 21511 5188
rect 21453 5179 21511 5185
rect 22281 5185 22293 5188
rect 22327 5185 22339 5219
rect 22281 5179 22339 5185
rect 22370 5176 22376 5228
rect 22428 5216 22434 5228
rect 22465 5219 22523 5225
rect 22465 5216 22477 5219
rect 22428 5188 22477 5216
rect 22428 5176 22434 5188
rect 22465 5185 22477 5188
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5185 22799 5219
rect 22741 5179 22799 5185
rect 21177 5151 21235 5157
rect 21177 5148 21189 5151
rect 16715 5120 20300 5148
rect 20824 5120 21189 5148
rect 16715 5117 16727 5120
rect 16669 5111 16727 5117
rect 16684 5080 16712 5111
rect 15672 5052 16712 5080
rect 11020 5040 11026 5052
rect 14752 5024 14780 5052
rect 20824 5024 20852 5120
rect 21177 5117 21189 5120
rect 21223 5117 21235 5151
rect 21177 5111 21235 5117
rect 22756 5080 22784 5179
rect 23014 5176 23020 5228
rect 23072 5176 23078 5228
rect 23566 5176 23572 5228
rect 23624 5176 23630 5228
rect 24118 5176 24124 5228
rect 24176 5216 24182 5228
rect 24305 5219 24363 5225
rect 24305 5216 24317 5219
rect 24176 5188 24317 5216
rect 24176 5176 24182 5188
rect 24305 5185 24317 5188
rect 24351 5185 24363 5219
rect 24305 5179 24363 5185
rect 25130 5176 25136 5228
rect 25188 5216 25194 5228
rect 25409 5219 25467 5225
rect 25409 5216 25421 5219
rect 25188 5188 25421 5216
rect 25188 5176 25194 5188
rect 25409 5185 25421 5188
rect 25455 5216 25467 5219
rect 25869 5219 25927 5225
rect 25869 5216 25881 5219
rect 25455 5188 25881 5216
rect 25455 5185 25467 5188
rect 25409 5179 25467 5185
rect 25869 5185 25881 5188
rect 25915 5185 25927 5219
rect 26068 5216 26096 5312
rect 27172 5256 27752 5284
rect 27172 5228 27200 5256
rect 26237 5219 26295 5225
rect 26237 5216 26249 5219
rect 25869 5179 25927 5185
rect 25976 5188 26249 5216
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 23750 5148 23756 5160
rect 23707 5120 23756 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 23750 5108 23756 5120
rect 23808 5108 23814 5160
rect 24394 5108 24400 5160
rect 24452 5108 24458 5160
rect 25501 5151 25559 5157
rect 25501 5117 25513 5151
rect 25547 5148 25559 5151
rect 25976 5148 26004 5188
rect 26237 5185 26249 5188
rect 26283 5185 26295 5219
rect 26237 5179 26295 5185
rect 26418 5176 26424 5228
rect 26476 5176 26482 5228
rect 27154 5176 27160 5228
rect 27212 5176 27218 5228
rect 27724 5225 27752 5256
rect 27341 5219 27399 5225
rect 27341 5185 27353 5219
rect 27387 5216 27399 5219
rect 27617 5219 27675 5225
rect 27617 5216 27629 5219
rect 27387 5188 27629 5216
rect 27387 5185 27399 5188
rect 27341 5179 27399 5185
rect 27617 5185 27629 5188
rect 27663 5185 27675 5219
rect 27617 5179 27675 5185
rect 27709 5219 27767 5225
rect 27709 5185 27721 5219
rect 27755 5185 27767 5219
rect 27709 5179 27767 5185
rect 27246 5148 27252 5160
rect 25547 5120 26004 5148
rect 26988 5120 27252 5148
rect 25547 5117 25559 5120
rect 25501 5111 25559 5117
rect 21284 5052 22784 5080
rect 24673 5083 24731 5089
rect 14734 4972 14740 5024
rect 14792 4972 14798 5024
rect 16022 4972 16028 5024
rect 16080 4972 16086 5024
rect 16298 4972 16304 5024
rect 16356 4972 16362 5024
rect 17126 4972 17132 5024
rect 17184 4972 17190 5024
rect 19978 4972 19984 5024
rect 20036 4972 20042 5024
rect 20806 4972 20812 5024
rect 20864 4972 20870 5024
rect 21284 5021 21312 5052
rect 22066 5024 22094 5052
rect 24673 5049 24685 5083
rect 24719 5080 24731 5083
rect 24946 5080 24952 5092
rect 24719 5052 24952 5080
rect 24719 5049 24731 5052
rect 24673 5043 24731 5049
rect 24946 5040 24952 5052
rect 25004 5040 25010 5092
rect 25777 5083 25835 5089
rect 25777 5049 25789 5083
rect 25823 5080 25835 5083
rect 26234 5080 26240 5092
rect 25823 5052 26240 5080
rect 25823 5049 25835 5052
rect 25777 5043 25835 5049
rect 26234 5040 26240 5052
rect 26292 5040 26298 5092
rect 21269 5015 21327 5021
rect 21269 4981 21281 5015
rect 21315 4981 21327 5015
rect 21269 4975 21327 4981
rect 21358 4972 21364 5024
rect 21416 4972 21422 5024
rect 22002 4972 22008 5024
rect 22060 4984 22094 5024
rect 23937 5015 23995 5021
rect 22060 4972 22066 4984
rect 23937 4981 23949 5015
rect 23983 5012 23995 5015
rect 24302 5012 24308 5024
rect 23983 4984 24308 5012
rect 23983 4981 23995 4984
rect 23937 4975 23995 4981
rect 24302 4972 24308 4984
rect 24360 4972 24366 5024
rect 25961 5015 26019 5021
rect 25961 4981 25973 5015
rect 26007 5012 26019 5015
rect 26988 5012 27016 5120
rect 27246 5108 27252 5120
rect 27304 5148 27310 5160
rect 27356 5148 27384 5179
rect 27798 5176 27804 5228
rect 27856 5216 27862 5228
rect 28000 5225 28028 5324
rect 28166 5244 28172 5296
rect 28224 5284 28230 5296
rect 28224 5256 29040 5284
rect 28224 5244 28230 5256
rect 28368 5225 28396 5256
rect 27893 5219 27951 5225
rect 27893 5216 27905 5219
rect 27856 5188 27905 5216
rect 27856 5176 27862 5188
rect 27893 5185 27905 5188
rect 27939 5185 27951 5219
rect 27893 5179 27951 5185
rect 27985 5219 28043 5225
rect 27985 5185 27997 5219
rect 28031 5185 28043 5219
rect 27985 5179 28043 5185
rect 28353 5219 28411 5225
rect 28353 5185 28365 5219
rect 28399 5185 28411 5219
rect 28353 5179 28411 5185
rect 27304 5120 27384 5148
rect 27433 5151 27491 5157
rect 27304 5108 27310 5120
rect 27433 5117 27445 5151
rect 27479 5148 27491 5151
rect 27522 5148 27528 5160
rect 27479 5120 27528 5148
rect 27479 5117 27491 5120
rect 27433 5111 27491 5117
rect 27522 5108 27528 5120
rect 27580 5108 27586 5160
rect 27908 5148 27936 5179
rect 28442 5176 28448 5228
rect 28500 5176 28506 5228
rect 28629 5219 28687 5225
rect 28629 5185 28641 5219
rect 28675 5185 28687 5219
rect 28629 5179 28687 5185
rect 28721 5219 28779 5225
rect 28721 5185 28733 5219
rect 28767 5216 28779 5219
rect 28902 5216 28908 5228
rect 28767 5188 28908 5216
rect 28767 5185 28779 5188
rect 28721 5179 28779 5185
rect 28534 5148 28540 5160
rect 27908 5120 28540 5148
rect 28534 5108 28540 5120
rect 28592 5148 28598 5160
rect 28644 5148 28672 5179
rect 28902 5176 28908 5188
rect 28960 5176 28966 5228
rect 29012 5216 29040 5256
rect 29546 5244 29552 5296
rect 29604 5284 29610 5296
rect 30377 5287 30435 5293
rect 30377 5284 30389 5287
rect 29604 5256 30389 5284
rect 29604 5244 29610 5256
rect 30377 5253 30389 5256
rect 30423 5253 30435 5287
rect 30377 5247 30435 5253
rect 30834 5244 30840 5296
rect 30892 5244 30898 5296
rect 29365 5219 29423 5225
rect 29365 5216 29377 5219
rect 29012 5188 29377 5216
rect 29365 5185 29377 5188
rect 29411 5185 29423 5219
rect 29365 5179 29423 5185
rect 28592 5120 28672 5148
rect 28920 5148 28948 5176
rect 29273 5151 29331 5157
rect 29273 5148 29285 5151
rect 28920 5120 29285 5148
rect 28592 5108 28598 5120
rect 29273 5117 29285 5120
rect 29319 5117 29331 5151
rect 29273 5111 29331 5117
rect 30098 5108 30104 5160
rect 30156 5108 30162 5160
rect 28905 5083 28963 5089
rect 28905 5049 28917 5083
rect 28951 5080 28963 5083
rect 29086 5080 29092 5092
rect 28951 5052 29092 5080
rect 28951 5049 28963 5052
rect 28905 5043 28963 5049
rect 29086 5040 29092 5052
rect 29144 5040 29150 5092
rect 26007 4984 27016 5012
rect 26007 4981 26019 4984
rect 25961 4975 26019 4981
rect 28994 4972 29000 5024
rect 29052 4972 29058 5024
rect 31846 4972 31852 5024
rect 31904 4972 31910 5024
rect 1104 4922 35248 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 35248 4922
rect 1104 4848 35248 4870
rect 11146 4768 11152 4820
rect 11204 4768 11210 4820
rect 16298 4768 16304 4820
rect 16356 4768 16362 4820
rect 16574 4768 16580 4820
rect 16632 4768 16638 4820
rect 17126 4768 17132 4820
rect 17184 4768 17190 4820
rect 18230 4768 18236 4820
rect 18288 4768 18294 4820
rect 19978 4768 19984 4820
rect 20036 4768 20042 4820
rect 27154 4768 27160 4820
rect 27212 4768 27218 4820
rect 7190 4632 7196 4684
rect 7248 4632 7254 4684
rect 8941 4675 8999 4681
rect 8941 4641 8953 4675
rect 8987 4672 8999 4675
rect 9306 4672 9312 4684
rect 8987 4644 9312 4672
rect 8987 4641 8999 4644
rect 8941 4635 8999 4641
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10468 4644 10977 4672
rect 10468 4632 10474 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 12250 4632 12256 4684
rect 12308 4672 12314 4684
rect 12897 4675 12955 4681
rect 12897 4672 12909 4675
rect 12308 4644 12909 4672
rect 12308 4632 12314 4644
rect 12897 4641 12909 4644
rect 12943 4641 12955 4675
rect 16316 4672 16344 4768
rect 16393 4675 16451 4681
rect 16393 4672 16405 4675
rect 16316 4644 16405 4672
rect 12897 4635 12955 4641
rect 16393 4641 16405 4644
rect 16439 4641 16451 4675
rect 16393 4635 16451 4641
rect 5166 4564 5172 4616
rect 5224 4564 5230 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6604 4576 8340 4604
rect 10350 4590 11546 4604
rect 10350 4576 11560 4590
rect 6604 4564 6610 4576
rect 5184 4468 5212 4564
rect 8312 4548 8340 4576
rect 5442 4496 5448 4548
rect 5500 4496 5506 4548
rect 8294 4496 8300 4548
rect 8352 4496 8358 4548
rect 9214 4496 9220 4548
rect 9272 4496 9278 4548
rect 6362 4468 6368 4480
rect 5184 4440 6368 4468
rect 6362 4428 6368 4440
rect 6420 4428 6426 4480
rect 11532 4468 11560 4576
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14185 4607 14243 4613
rect 14185 4604 14197 4607
rect 13780 4576 14197 4604
rect 13780 4564 13786 4576
rect 14185 4573 14197 4576
rect 14231 4573 14243 4607
rect 14185 4567 14243 4573
rect 14734 4564 14740 4616
rect 14792 4564 14798 4616
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4604 16543 4607
rect 16592 4604 16620 4768
rect 16531 4576 16620 4604
rect 17144 4604 17172 4768
rect 17865 4675 17923 4681
rect 17865 4641 17877 4675
rect 17911 4672 17923 4675
rect 18248 4672 18276 4768
rect 19426 4700 19432 4752
rect 19484 4740 19490 4752
rect 19889 4743 19947 4749
rect 19889 4740 19901 4743
rect 19484 4712 19901 4740
rect 19484 4700 19490 4712
rect 19889 4709 19901 4712
rect 19935 4709 19947 4743
rect 19889 4703 19947 4709
rect 18693 4675 18751 4681
rect 18693 4672 18705 4675
rect 17911 4644 18705 4672
rect 17911 4641 17923 4644
rect 17865 4635 17923 4641
rect 18693 4641 18705 4644
rect 18739 4641 18751 4675
rect 18693 4635 18751 4641
rect 19613 4675 19671 4681
rect 19613 4641 19625 4675
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 17773 4607 17831 4613
rect 17773 4604 17785 4607
rect 17144 4576 17785 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 17773 4573 17785 4576
rect 17819 4604 17831 4607
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 17819 4576 18245 4604
rect 17819 4573 17831 4576
rect 17773 4567 17831 4573
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18601 4607 18659 4613
rect 18601 4573 18613 4607
rect 18647 4604 18659 4607
rect 18877 4607 18935 4613
rect 18647 4576 18736 4604
rect 18647 4573 18659 4576
rect 18601 4567 18659 4573
rect 12621 4539 12679 4545
rect 12621 4505 12633 4539
rect 12667 4536 12679 4539
rect 14458 4536 14464 4548
rect 12667 4508 14464 4536
rect 12667 4505 12679 4508
rect 12621 4499 12679 4505
rect 14458 4496 14464 4508
rect 14516 4496 14522 4548
rect 15930 4536 15936 4548
rect 15686 4508 15936 4536
rect 15930 4496 15936 4508
rect 15988 4536 15994 4548
rect 18708 4536 18736 4576
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19521 4607 19579 4613
rect 19521 4604 19533 4607
rect 18923 4576 19533 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19521 4573 19533 4576
rect 19567 4573 19579 4607
rect 19628 4604 19656 4635
rect 19996 4613 20024 4768
rect 20257 4743 20315 4749
rect 20257 4709 20269 4743
rect 20303 4709 20315 4743
rect 20257 4703 20315 4709
rect 21177 4743 21235 4749
rect 21177 4709 21189 4743
rect 21223 4740 21235 4743
rect 22094 4740 22100 4752
rect 21223 4712 22100 4740
rect 21223 4709 21235 4712
rect 21177 4703 21235 4709
rect 19981 4607 20039 4613
rect 19981 4604 19993 4607
rect 19628 4576 19993 4604
rect 19521 4567 19579 4573
rect 19981 4573 19993 4576
rect 20027 4573 20039 4607
rect 20272 4604 20300 4703
rect 22094 4700 22100 4712
rect 22152 4700 22158 4752
rect 27525 4743 27583 4749
rect 27525 4709 27537 4743
rect 27571 4709 27583 4743
rect 27525 4703 27583 4709
rect 20901 4675 20959 4681
rect 20901 4641 20913 4675
rect 20947 4672 20959 4675
rect 21358 4672 21364 4684
rect 20947 4644 21364 4672
rect 20947 4641 20959 4644
rect 20901 4635 20959 4641
rect 21358 4632 21364 4644
rect 21416 4632 21422 4684
rect 22002 4632 22008 4684
rect 22060 4672 22066 4684
rect 22189 4675 22247 4681
rect 22060 4644 22140 4672
rect 22060 4632 22066 4644
rect 20806 4604 20812 4616
rect 20272 4576 20812 4604
rect 19981 4567 20039 4573
rect 15988 4508 18736 4536
rect 19536 4536 19564 4567
rect 20806 4564 20812 4576
rect 20864 4564 20870 4616
rect 22112 4613 22140 4644
rect 22189 4641 22201 4675
rect 22235 4672 22247 4675
rect 22370 4672 22376 4684
rect 22235 4644 22376 4672
rect 22235 4641 22247 4644
rect 22189 4635 22247 4641
rect 22370 4632 22376 4644
rect 22428 4632 22434 4684
rect 27246 4632 27252 4684
rect 27304 4632 27310 4684
rect 27540 4672 27568 4703
rect 27617 4675 27675 4681
rect 27617 4672 27629 4675
rect 27540 4644 27629 4672
rect 27617 4641 27629 4644
rect 27663 4641 27675 4675
rect 27617 4635 27675 4641
rect 22097 4607 22155 4613
rect 22097 4573 22109 4607
rect 22143 4573 22155 4607
rect 22097 4567 22155 4573
rect 25590 4564 25596 4616
rect 25648 4564 25654 4616
rect 27157 4607 27215 4613
rect 27157 4573 27169 4607
rect 27203 4604 27215 4607
rect 27430 4604 27436 4616
rect 27203 4576 27436 4604
rect 27203 4573 27215 4576
rect 27157 4567 27215 4573
rect 27430 4564 27436 4576
rect 27488 4564 27494 4616
rect 27706 4564 27712 4616
rect 27764 4604 27770 4616
rect 27801 4607 27859 4613
rect 27801 4604 27813 4607
rect 27764 4576 27813 4604
rect 27764 4564 27770 4576
rect 27801 4573 27813 4576
rect 27847 4573 27859 4607
rect 27801 4567 27859 4573
rect 20257 4539 20315 4545
rect 20257 4536 20269 4539
rect 19536 4508 20269 4536
rect 15988 4496 15994 4508
rect 13262 4468 13268 4480
rect 11532 4440 13268 4468
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 16850 4428 16856 4480
rect 16908 4428 16914 4480
rect 18138 4428 18144 4480
rect 18196 4428 18202 4480
rect 18708 4468 18736 4508
rect 20257 4505 20269 4508
rect 20303 4505 20315 4539
rect 20257 4499 20315 4505
rect 22066 4508 24808 4536
rect 20073 4471 20131 4477
rect 20073 4468 20085 4471
rect 18708 4440 20085 4468
rect 20073 4437 20085 4440
rect 20119 4468 20131 4471
rect 22066 4468 22094 4508
rect 20119 4440 22094 4468
rect 20119 4437 20131 4440
rect 20073 4431 20131 4437
rect 22462 4428 22468 4480
rect 22520 4428 22526 4480
rect 24780 4468 24808 4508
rect 24854 4496 24860 4548
rect 24912 4496 24918 4548
rect 27798 4468 27804 4480
rect 24780 4440 27804 4468
rect 27798 4428 27804 4440
rect 27856 4428 27862 4480
rect 27982 4428 27988 4480
rect 28040 4428 28046 4480
rect 1104 4378 35236 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 35236 4378
rect 1104 4304 35236 4326
rect 15930 4224 15936 4276
rect 15988 4224 15994 4276
rect 29178 4264 29184 4276
rect 29012 4236 29184 4264
rect 8202 4156 8208 4208
rect 8260 4196 8266 4208
rect 8389 4199 8447 4205
rect 8389 4196 8401 4199
rect 8260 4168 8401 4196
rect 8260 4156 8266 4168
rect 8389 4165 8401 4168
rect 8435 4165 8447 4199
rect 8389 4159 8447 4165
rect 11977 4199 12035 4205
rect 11977 4165 11989 4199
rect 12023 4196 12035 4199
rect 12066 4196 12072 4208
rect 12023 4168 12072 4196
rect 12023 4165 12035 4168
rect 11977 4159 12035 4165
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 13262 4156 13268 4208
rect 13320 4156 13326 4208
rect 8294 4128 8300 4140
rect 7774 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 10502 4128 10508 4140
rect 9890 4100 10508 4128
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 15381 4131 15439 4137
rect 15381 4097 15393 4131
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 6362 4020 6368 4072
rect 6420 4020 6426 4072
rect 6638 4020 6644 4072
rect 6696 4020 6702 4072
rect 8481 4063 8539 4069
rect 8481 4029 8493 4063
rect 8527 4029 8539 4063
rect 8481 4023 8539 4029
rect 6380 3924 6408 4020
rect 8496 3936 8524 4023
rect 8754 4020 8760 4072
rect 8812 4020 8818 4072
rect 10226 4020 10232 4072
rect 10284 4020 10290 4072
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4060 13783 4063
rect 14001 4063 14059 4069
rect 13771 4032 13952 4060
rect 13771 4029 13783 4032
rect 13725 4023 13783 4029
rect 13924 3992 13952 4032
rect 14001 4029 14013 4063
rect 14047 4060 14059 4063
rect 14090 4060 14096 4072
rect 14047 4032 14096 4060
rect 14047 4029 14059 4032
rect 14001 4023 14059 4029
rect 14090 4020 14096 4032
rect 14148 4020 14154 4072
rect 15289 4063 15347 4069
rect 15289 4029 15301 4063
rect 15335 4029 15347 4063
rect 15396 4060 15424 4091
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15528 4100 15853 4128
rect 15528 4088 15534 4100
rect 15841 4097 15853 4100
rect 15887 4097 15899 4131
rect 15948 4128 15976 4224
rect 29012 4196 29040 4236
rect 29178 4224 29184 4236
rect 29236 4264 29242 4276
rect 30098 4264 30104 4276
rect 29236 4236 30104 4264
rect 29236 4224 29242 4236
rect 30098 4224 30104 4236
rect 30156 4224 30162 4276
rect 30374 4196 30380 4208
rect 28828 4168 29040 4196
rect 30314 4182 30380 4196
rect 30300 4168 30380 4182
rect 16025 4131 16083 4137
rect 16025 4128 16037 4131
rect 15948 4100 16037 4128
rect 15841 4091 15899 4097
rect 16025 4097 16037 4100
rect 16071 4097 16083 4131
rect 16025 4091 16083 4097
rect 16758 4088 16764 4140
rect 16816 4088 16822 4140
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 23566 4088 23572 4140
rect 23624 4088 23630 4140
rect 23934 4088 23940 4140
rect 23992 4088 23998 4140
rect 26510 4088 26516 4140
rect 26568 4088 26574 4140
rect 26694 4088 26700 4140
rect 26752 4128 26758 4140
rect 28828 4137 28856 4168
rect 26973 4131 27031 4137
rect 26973 4128 26985 4131
rect 26752 4100 26985 4128
rect 26752 4088 26758 4100
rect 26973 4097 26985 4100
rect 27019 4097 27031 4131
rect 26973 4091 27031 4097
rect 28813 4131 28871 4137
rect 28813 4097 28825 4131
rect 28859 4097 28871 4131
rect 28813 4091 28871 4097
rect 15933 4063 15991 4069
rect 15933 4060 15945 4063
rect 15396 4032 15945 4060
rect 15289 4023 15347 4029
rect 15933 4029 15945 4032
rect 15979 4029 15991 4063
rect 15933 4023 15991 4029
rect 15304 3992 15332 4023
rect 17218 4020 17224 4072
rect 17276 4020 17282 4072
rect 18414 4020 18420 4072
rect 18472 4060 18478 4072
rect 18693 4063 18751 4069
rect 18693 4060 18705 4063
rect 18472 4032 18705 4060
rect 18472 4020 18478 4032
rect 18693 4029 18705 4032
rect 18739 4029 18751 4063
rect 18693 4023 18751 4029
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 22465 4063 22523 4069
rect 22465 4060 22477 4063
rect 22244 4032 22477 4060
rect 22244 4020 22250 4032
rect 22465 4029 22477 4032
rect 22511 4029 22523 4063
rect 22465 4023 22523 4029
rect 23290 4020 23296 4072
rect 23348 4060 23354 4072
rect 24213 4063 24271 4069
rect 24213 4060 24225 4063
rect 23348 4032 24225 4060
rect 23348 4020 23354 4032
rect 24213 4029 24225 4032
rect 24259 4029 24271 4063
rect 24213 4023 24271 4029
rect 25222 4020 25228 4072
rect 25280 4060 25286 4072
rect 25501 4063 25559 4069
rect 25501 4060 25513 4063
rect 25280 4032 25513 4060
rect 25280 4020 25286 4032
rect 25501 4029 25513 4032
rect 25547 4029 25559 4063
rect 25501 4023 25559 4029
rect 26418 4020 26424 4072
rect 26476 4060 26482 4072
rect 27433 4063 27491 4069
rect 27433 4060 27445 4063
rect 26476 4032 27445 4060
rect 26476 4020 26482 4032
rect 27433 4029 27445 4032
rect 27479 4029 27491 4063
rect 27433 4023 27491 4029
rect 29086 4020 29092 4072
rect 29144 4020 29150 4072
rect 16022 3992 16028 4004
rect 13924 3964 14412 3992
rect 15304 3964 16028 3992
rect 14384 3936 14412 3964
rect 16022 3952 16028 3964
rect 16080 3952 16086 4004
rect 6822 3924 6828 3936
rect 6380 3896 6828 3924
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 9306 3924 9312 3936
rect 8536 3896 9312 3924
rect 8536 3884 8542 3896
rect 9306 3884 9312 3896
rect 9364 3884 9370 3936
rect 14366 3884 14372 3936
rect 14424 3884 14430 3936
rect 15654 3884 15660 3936
rect 15712 3884 15718 3936
rect 27706 3884 27712 3936
rect 27764 3924 27770 3936
rect 30300 3924 30328 4168
rect 30374 4156 30380 4168
rect 30432 4196 30438 4208
rect 30834 4196 30840 4208
rect 30432 4168 30840 4196
rect 30432 4156 30438 4168
rect 30834 4156 30840 4168
rect 30892 4156 30898 4208
rect 27764 3896 30328 3924
rect 27764 3884 27770 3896
rect 30558 3884 30564 3936
rect 30616 3884 30622 3936
rect 1104 3834 35248 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 35248 3834
rect 1104 3760 35248 3782
rect 5074 3720 5080 3732
rect 4632 3692 5080 3720
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4632 3593 4660 3692
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 8662 3720 8668 3732
rect 6656 3692 8668 3720
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4212 3556 4629 3584
rect 4212 3544 4218 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 6546 3516 6552 3528
rect 6052 3488 6552 3516
rect 6052 3476 6058 3488
rect 6546 3476 6552 3488
rect 6604 3476 6610 3528
rect 6656 3525 6684 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 13262 3720 13268 3732
rect 11164 3692 13268 3720
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3584 8815 3587
rect 9030 3584 9036 3596
rect 8803 3556 9036 3584
rect 8803 3553 8815 3556
rect 8757 3547 8815 3553
rect 9030 3544 9036 3556
rect 9088 3544 9094 3596
rect 10502 3584 10508 3596
rect 9140 3556 10508 3584
rect 6641 3519 6699 3525
rect 6641 3485 6653 3519
rect 6687 3485 6699 3519
rect 6641 3479 6699 3485
rect 6733 3519 6791 3525
rect 6733 3485 6745 3519
rect 6779 3485 6791 3519
rect 8294 3516 8300 3528
rect 8142 3488 8300 3516
rect 6733 3479 6791 3485
rect 4890 3408 4896 3460
rect 4948 3408 4954 3460
rect 6748 3448 6776 3479
rect 8294 3476 8300 3488
rect 8352 3516 8358 3528
rect 9140 3516 9168 3556
rect 10502 3544 10508 3556
rect 10560 3584 10566 3596
rect 11164 3584 11192 3692
rect 13262 3680 13268 3692
rect 13320 3680 13326 3732
rect 15654 3680 15660 3732
rect 15712 3680 15718 3732
rect 18049 3723 18107 3729
rect 18049 3689 18061 3723
rect 18095 3720 18107 3723
rect 18230 3720 18236 3732
rect 18095 3692 18236 3720
rect 18095 3689 18107 3692
rect 18049 3683 18107 3689
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 23658 3720 23664 3732
rect 22204 3692 23664 3720
rect 10560 3556 11192 3584
rect 10560 3544 10566 3556
rect 8352 3488 9168 3516
rect 8352 3476 8358 3488
rect 9306 3476 9312 3528
rect 9364 3516 9370 3528
rect 9769 3519 9827 3525
rect 9769 3516 9781 3519
rect 9364 3488 9781 3516
rect 9364 3476 9370 3488
rect 9769 3485 9781 3488
rect 9815 3485 9827 3519
rect 11164 3502 11192 3556
rect 11793 3587 11851 3593
rect 11793 3553 11805 3587
rect 11839 3584 11851 3587
rect 12894 3584 12900 3596
rect 11839 3556 12900 3584
rect 11839 3553 11851 3556
rect 11793 3547 11851 3553
rect 12894 3544 12900 3556
rect 12952 3544 12958 3596
rect 15672 3584 15700 3680
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 15672 3556 16589 3584
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 18690 3584 18696 3596
rect 16577 3547 16635 3553
rect 17696 3556 18696 3584
rect 11885 3519 11943 3525
rect 9769 3479 9827 3485
rect 11885 3485 11897 3519
rect 11931 3516 11943 3519
rect 12342 3516 12348 3528
rect 11931 3488 12348 3516
rect 11931 3485 11943 3488
rect 11885 3479 11943 3485
rect 6748 3420 6868 3448
rect 6840 3392 6868 3420
rect 7006 3408 7012 3460
rect 7064 3408 7070 3460
rect 6822 3340 6828 3392
rect 6880 3340 6886 3392
rect 9784 3380 9812 3479
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3516 13967 3519
rect 14090 3516 14096 3528
rect 13955 3488 14096 3516
rect 13955 3485 13967 3488
rect 13909 3479 13967 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 16301 3519 16359 3525
rect 16301 3485 16313 3519
rect 16347 3485 16359 3519
rect 16301 3479 16359 3485
rect 10042 3408 10048 3460
rect 10100 3408 10106 3460
rect 12894 3408 12900 3460
rect 12952 3408 12958 3460
rect 13633 3451 13691 3457
rect 13633 3417 13645 3451
rect 13679 3448 13691 3451
rect 13998 3448 14004 3460
rect 13679 3420 14004 3448
rect 13679 3417 13691 3420
rect 13633 3411 13691 3417
rect 13998 3408 14004 3420
rect 14056 3408 14062 3460
rect 11054 3380 11060 3392
rect 9784 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 12250 3340 12256 3392
rect 12308 3380 12314 3392
rect 14108 3380 14136 3476
rect 16316 3448 16344 3479
rect 16574 3448 16580 3460
rect 16316 3420 16580 3448
rect 16574 3408 16580 3420
rect 16632 3408 16638 3460
rect 12308 3352 14136 3380
rect 12308 3340 12314 3352
rect 16482 3340 16488 3392
rect 16540 3380 16546 3392
rect 17696 3380 17724 3556
rect 18690 3544 18696 3556
rect 18748 3584 18754 3596
rect 22204 3593 22232 3692
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 23934 3680 23940 3732
rect 23992 3680 23998 3732
rect 24302 3680 24308 3732
rect 24360 3680 24366 3732
rect 24394 3680 24400 3732
rect 24452 3720 24458 3732
rect 26145 3723 26203 3729
rect 24452 3692 25728 3720
rect 24452 3680 24458 3692
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 18748 3556 19349 3584
rect 18748 3544 18754 3556
rect 19337 3553 19349 3556
rect 19383 3553 19395 3587
rect 22189 3587 22247 3593
rect 22189 3584 22201 3587
rect 19337 3547 19395 3553
rect 21836 3556 22201 3584
rect 21836 3528 21864 3556
rect 22189 3553 22201 3556
rect 22235 3553 22247 3587
rect 22189 3547 22247 3553
rect 22462 3544 22468 3596
rect 22520 3544 22526 3596
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 17862 3408 17868 3460
rect 17920 3448 17926 3460
rect 18325 3451 18383 3457
rect 18325 3448 18337 3451
rect 17920 3420 18337 3448
rect 17920 3408 17926 3420
rect 18325 3417 18337 3420
rect 18371 3417 18383 3451
rect 18325 3411 18383 3417
rect 16540 3352 17724 3380
rect 18616 3380 18644 3479
rect 19886 3476 19892 3528
rect 19944 3476 19950 3528
rect 21818 3476 21824 3528
rect 21876 3476 21882 3528
rect 21910 3476 21916 3528
rect 21968 3476 21974 3528
rect 23676 3516 23704 3680
rect 24320 3584 24348 3680
rect 24673 3587 24731 3593
rect 24673 3584 24685 3587
rect 24320 3556 24685 3584
rect 24673 3553 24685 3556
rect 24719 3553 24731 3587
rect 25700 3584 25728 3692
rect 26145 3689 26157 3723
rect 26191 3720 26203 3723
rect 26510 3720 26516 3732
rect 26191 3692 26516 3720
rect 26191 3689 26203 3692
rect 26145 3683 26203 3689
rect 26510 3680 26516 3692
rect 26568 3680 26574 3732
rect 28810 3680 28816 3732
rect 28868 3720 28874 3732
rect 29178 3720 29184 3732
rect 28868 3692 29184 3720
rect 28868 3680 28874 3692
rect 29178 3680 29184 3692
rect 29236 3680 29242 3732
rect 26234 3612 26240 3664
rect 26292 3612 26298 3664
rect 28718 3612 28724 3664
rect 28776 3652 28782 3664
rect 28776 3624 29224 3652
rect 28776 3612 28782 3624
rect 26252 3584 26280 3612
rect 26513 3587 26571 3593
rect 26513 3584 26525 3587
rect 25700 3556 25912 3584
rect 26252 3556 26525 3584
rect 24673 3547 24731 3553
rect 24394 3516 24400 3528
rect 23676 3488 24400 3516
rect 24394 3476 24400 3488
rect 24452 3476 24458 3528
rect 25884 3516 25912 3556
rect 26513 3553 26525 3556
rect 26559 3553 26571 3587
rect 26513 3547 26571 3553
rect 27985 3587 28043 3593
rect 27985 3553 27997 3587
rect 28031 3584 28043 3587
rect 29086 3584 29092 3596
rect 28031 3556 29092 3584
rect 28031 3553 28043 3556
rect 27985 3547 28043 3553
rect 29086 3544 29092 3556
rect 29144 3544 29150 3596
rect 29196 3584 29224 3624
rect 29270 3612 29276 3664
rect 29328 3652 29334 3664
rect 29328 3624 31524 3652
rect 29328 3612 29334 3624
rect 31496 3593 31524 3624
rect 30009 3587 30067 3593
rect 30009 3584 30021 3587
rect 29196 3556 30021 3584
rect 30009 3553 30021 3556
rect 30055 3553 30067 3587
rect 30009 3547 30067 3553
rect 31481 3587 31539 3593
rect 31481 3553 31493 3587
rect 31527 3553 31539 3587
rect 31481 3547 31539 3553
rect 32306 3544 32312 3596
rect 32364 3584 32370 3596
rect 32953 3587 33011 3593
rect 32953 3584 32965 3587
rect 32364 3556 32965 3584
rect 32364 3544 32370 3556
rect 32953 3553 32965 3556
rect 32999 3553 33011 3587
rect 32953 3547 33011 3553
rect 26234 3516 26240 3528
rect 25884 3488 26240 3516
rect 26234 3476 26240 3488
rect 26292 3476 26298 3528
rect 28721 3519 28779 3525
rect 28721 3516 28733 3519
rect 27816 3488 28733 3516
rect 21082 3408 21088 3460
rect 21140 3408 21146 3460
rect 22922 3408 22928 3460
rect 22980 3408 22986 3460
rect 25314 3408 25320 3460
rect 25372 3408 25378 3460
rect 26970 3408 26976 3460
rect 27028 3408 27034 3460
rect 27816 3380 27844 3488
rect 28721 3485 28733 3488
rect 28767 3516 28779 3519
rect 28767 3488 29040 3516
rect 28767 3485 28779 3488
rect 28721 3479 28779 3485
rect 18616 3352 27844 3380
rect 16540 3340 16546 3352
rect 28810 3340 28816 3392
rect 28868 3380 28874 3392
rect 28905 3383 28963 3389
rect 28905 3380 28917 3383
rect 28868 3352 28917 3380
rect 28868 3340 28874 3352
rect 28905 3349 28917 3352
rect 28951 3349 28963 3383
rect 29012 3380 29040 3488
rect 29178 3476 29184 3528
rect 29236 3516 29242 3528
rect 29549 3519 29607 3525
rect 29549 3516 29561 3519
rect 29236 3488 29561 3516
rect 29236 3476 29242 3488
rect 29549 3485 29561 3488
rect 29595 3485 29607 3519
rect 29549 3479 29607 3485
rect 31018 3476 31024 3528
rect 31076 3476 31082 3528
rect 31846 3476 31852 3528
rect 31904 3516 31910 3528
rect 32493 3519 32551 3525
rect 32493 3516 32505 3519
rect 31904 3488 32505 3516
rect 31904 3476 31910 3488
rect 32493 3485 32505 3488
rect 32539 3485 32551 3519
rect 32493 3479 32551 3485
rect 33594 3380 33600 3392
rect 29012 3352 33600 3380
rect 28905 3343 28963 3349
rect 33594 3340 33600 3352
rect 33652 3340 33658 3392
rect 1104 3290 35236 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 35236 3290
rect 1104 3216 35236 3238
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 8478 3176 8484 3188
rect 6880 3148 8484 3176
rect 6880 3136 6886 3148
rect 5994 3108 6000 3120
rect 5658 3080 6000 3108
rect 5994 3068 6000 3080
rect 6052 3068 6058 3120
rect 6932 3049 6960 3148
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8754 3136 8760 3188
rect 8812 3176 8818 3188
rect 13173 3179 13231 3185
rect 13173 3176 13185 3179
rect 8812 3148 13185 3176
rect 8812 3136 8818 3148
rect 13173 3145 13185 3148
rect 13219 3145 13231 3179
rect 13173 3139 13231 3145
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 15562 3176 15568 3188
rect 13320 3148 15568 3176
rect 13320 3136 13326 3148
rect 8938 3068 8944 3120
rect 8996 3068 9002 3120
rect 10502 3108 10508 3120
rect 10350 3080 10508 3108
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 10781 3111 10839 3117
rect 10781 3077 10793 3111
rect 10827 3108 10839 3111
rect 11146 3108 11152 3120
rect 10827 3080 11152 3108
rect 10827 3077 10839 3080
rect 10781 3071 10839 3077
rect 11146 3068 11152 3080
rect 11204 3068 11210 3120
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 13280 3108 13308 3136
rect 12952 3080 13308 3108
rect 12952 3068 12958 3080
rect 13538 3068 13544 3120
rect 13596 3068 13602 3120
rect 14936 3108 14964 3148
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 16574 3136 16580 3188
rect 16632 3176 16638 3188
rect 17862 3176 17868 3188
rect 16632 3148 17868 3176
rect 16632 3136 16638 3148
rect 14858 3080 14964 3108
rect 15289 3111 15347 3117
rect 15289 3077 15301 3111
rect 15335 3108 15347 3111
rect 16666 3108 16672 3120
rect 15335 3080 16672 3108
rect 15335 3077 15347 3080
rect 15289 3071 15347 3077
rect 16666 3068 16672 3080
rect 16724 3068 16730 3120
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 11974 3000 11980 3052
rect 12032 3000 12038 3052
rect 12250 3000 12256 3052
rect 12308 3000 12314 3052
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13357 3043 13415 3049
rect 13357 3040 13369 3043
rect 13136 3012 13369 3040
rect 13136 3000 13142 3012
rect 13357 3009 13369 3012
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 15565 3043 15623 3049
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 16776 3040 16804 3148
rect 17862 3136 17868 3148
rect 17920 3136 17926 3188
rect 21545 3179 21603 3185
rect 19996 3148 21496 3176
rect 18138 3068 18144 3120
rect 18196 3108 18202 3120
rect 18233 3111 18291 3117
rect 18233 3108 18245 3111
rect 18196 3080 18245 3108
rect 18196 3068 18202 3080
rect 18233 3077 18245 3080
rect 18279 3077 18291 3111
rect 19996 3108 20024 3148
rect 19458 3080 20024 3108
rect 20456 3108 20484 3148
rect 21468 3108 21496 3148
rect 21545 3145 21557 3179
rect 21591 3176 21603 3179
rect 21910 3176 21916 3188
rect 21591 3148 21916 3176
rect 21591 3145 21603 3148
rect 21545 3139 21603 3145
rect 21910 3136 21916 3148
rect 21968 3136 21974 3188
rect 22922 3176 22928 3188
rect 22020 3148 22928 3176
rect 22020 3108 22048 3148
rect 20456 3080 20562 3108
rect 21468 3080 22048 3108
rect 18233 3071 18291 3077
rect 22094 3068 22100 3120
rect 22152 3068 22158 3120
rect 22480 3108 22508 3148
rect 22922 3136 22928 3148
rect 22980 3176 22986 3188
rect 25314 3176 25320 3188
rect 22980 3148 25320 3176
rect 22980 3136 22986 3148
rect 22480 3080 22586 3108
rect 23474 3068 23480 3120
rect 23532 3108 23538 3120
rect 23937 3111 23995 3117
rect 23937 3108 23949 3111
rect 23532 3080 23949 3108
rect 23532 3068 23538 3080
rect 23937 3077 23949 3080
rect 23983 3077 23995 3111
rect 24320 3108 24348 3148
rect 25314 3136 25320 3148
rect 25372 3136 25378 3188
rect 25409 3179 25467 3185
rect 25409 3145 25421 3179
rect 25455 3176 25467 3179
rect 25590 3176 25596 3188
rect 25455 3148 25596 3176
rect 25455 3145 25467 3148
rect 25409 3139 25467 3145
rect 25590 3136 25596 3148
rect 25648 3136 25654 3188
rect 27522 3136 27528 3188
rect 27580 3176 27586 3188
rect 28721 3179 28779 3185
rect 27580 3148 28580 3176
rect 27580 3136 27586 3148
rect 25332 3108 25360 3136
rect 26970 3108 26976 3120
rect 24320 3080 24426 3108
rect 25332 3080 26976 3108
rect 23937 3071 23995 3077
rect 26970 3068 26976 3080
rect 27028 3108 27034 3120
rect 27706 3108 27712 3120
rect 27028 3080 27712 3108
rect 27028 3068 27034 3080
rect 27706 3068 27712 3080
rect 27764 3068 27770 3120
rect 15611 3012 16804 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 4154 2932 4160 2984
rect 4212 2932 4218 2984
rect 4430 2932 4436 2984
rect 4488 2932 4494 2984
rect 6181 2975 6239 2981
rect 6181 2941 6193 2975
rect 6227 2941 6239 2975
rect 6181 2935 6239 2941
rect 6196 2836 6224 2935
rect 7190 2932 7196 2984
rect 7248 2932 7254 2984
rect 9033 2975 9091 2981
rect 9033 2941 9045 2975
rect 9079 2972 9091 2975
rect 10318 2972 10324 2984
rect 9079 2944 10324 2972
rect 9079 2941 9091 2944
rect 9033 2935 9091 2941
rect 10318 2932 10324 2944
rect 10376 2932 10382 2984
rect 11054 2932 11060 2984
rect 11112 2972 11118 2984
rect 12268 2972 12296 3000
rect 11112 2944 12296 2972
rect 11112 2932 11118 2944
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 15580 2972 15608 3003
rect 23566 3000 23572 3052
rect 23624 3000 23630 3052
rect 23658 3000 23664 3052
rect 23716 3000 23722 3052
rect 26234 3000 26240 3052
rect 26292 3040 26298 3052
rect 28552 3040 28580 3148
rect 28721 3145 28733 3179
rect 28767 3176 28779 3179
rect 29178 3176 29184 3188
rect 28767 3148 29184 3176
rect 28767 3145 28779 3148
rect 28721 3139 28779 3145
rect 29178 3136 29184 3148
rect 29236 3136 29242 3188
rect 30558 3136 30564 3188
rect 30616 3176 30622 3188
rect 30616 3148 32168 3176
rect 30616 3136 30622 3148
rect 28994 3068 29000 3120
rect 29052 3108 29058 3120
rect 29089 3111 29147 3117
rect 29089 3108 29101 3111
rect 29052 3080 29101 3108
rect 29052 3068 29058 3080
rect 29089 3077 29101 3080
rect 29135 3077 29147 3111
rect 30374 3108 30380 3120
rect 30314 3080 30380 3108
rect 29089 3071 29147 3077
rect 30374 3068 30380 3080
rect 30432 3108 30438 3120
rect 30929 3111 30987 3117
rect 30929 3108 30941 3111
rect 30432 3080 30941 3108
rect 30432 3068 30438 3080
rect 30929 3077 30941 3080
rect 30975 3077 30987 3111
rect 30929 3071 30987 3077
rect 28810 3040 28816 3052
rect 26292 3012 27016 3040
rect 28552 3012 28816 3040
rect 26292 3000 26298 3012
rect 14148 2944 15608 2972
rect 17957 2975 18015 2981
rect 14148 2932 14154 2944
rect 17957 2941 17969 2975
rect 18003 2972 18015 2975
rect 19794 2972 19800 2984
rect 18003 2944 19800 2972
rect 18003 2941 18015 2944
rect 17957 2935 18015 2941
rect 19794 2932 19800 2944
rect 19852 2932 19858 2984
rect 20073 2975 20131 2981
rect 20073 2972 20085 2975
rect 19904 2944 20085 2972
rect 19426 2864 19432 2916
rect 19484 2904 19490 2916
rect 19904 2904 19932 2944
rect 20073 2941 20085 2944
rect 20119 2941 20131 2975
rect 20073 2935 20131 2941
rect 20162 2932 20168 2984
rect 20220 2972 20226 2984
rect 21818 2972 21824 2984
rect 20220 2944 21824 2972
rect 20220 2932 20226 2944
rect 21818 2932 21824 2944
rect 21876 2932 21882 2984
rect 23584 2913 23612 3000
rect 26988 2984 27016 3012
rect 28810 3000 28816 3012
rect 28868 3000 28874 3052
rect 32140 3049 32168 3148
rect 33594 3136 33600 3188
rect 33652 3136 33658 3188
rect 30653 3043 30711 3049
rect 30653 3009 30665 3043
rect 30699 3009 30711 3043
rect 30653 3003 30711 3009
rect 32125 3043 32183 3049
rect 32125 3009 32137 3043
rect 32171 3009 32183 3043
rect 32125 3003 32183 3009
rect 26878 2932 26884 2984
rect 26936 2932 26942 2984
rect 26970 2932 26976 2984
rect 27028 2932 27034 2984
rect 27798 2932 27804 2984
rect 27856 2972 27862 2984
rect 30668 2972 30696 3003
rect 33318 3000 33324 3052
rect 33376 3040 33382 3052
rect 33781 3043 33839 3049
rect 33781 3040 33793 3043
rect 33376 3012 33793 3040
rect 33376 3000 33382 3012
rect 33781 3009 33793 3012
rect 33827 3009 33839 3043
rect 33781 3003 33839 3009
rect 27856 2944 30696 2972
rect 27856 2932 27862 2944
rect 19484 2876 19932 2904
rect 23569 2907 23627 2913
rect 19484 2864 19490 2876
rect 23569 2873 23581 2907
rect 23615 2873 23627 2907
rect 26896 2904 26924 2932
rect 30668 2904 30696 2944
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 32585 2975 32643 2981
rect 32585 2972 32597 2975
rect 31352 2944 32597 2972
rect 31352 2932 31358 2944
rect 32585 2941 32597 2944
rect 32631 2941 32643 2975
rect 32585 2935 32643 2941
rect 26896 2876 27108 2904
rect 30668 2876 34284 2904
rect 23569 2867 23627 2873
rect 8570 2836 8576 2848
rect 6196 2808 8576 2836
rect 8570 2796 8576 2808
rect 8628 2796 8634 2848
rect 11790 2796 11796 2848
rect 11848 2796 11854 2848
rect 19705 2839 19763 2845
rect 19705 2805 19717 2839
rect 19751 2836 19763 2839
rect 21818 2836 21824 2848
rect 19751 2808 21824 2836
rect 19751 2805 19763 2808
rect 19705 2799 19763 2805
rect 21818 2796 21824 2808
rect 21876 2796 21882 2848
rect 27080 2836 27108 2876
rect 34256 2848 34284 2876
rect 27230 2839 27288 2845
rect 27230 2836 27242 2839
rect 27080 2808 27242 2836
rect 27230 2805 27242 2808
rect 27276 2805 27288 2839
rect 27230 2799 27288 2805
rect 27430 2796 27436 2848
rect 27488 2836 27494 2848
rect 30374 2836 30380 2848
rect 27488 2808 30380 2836
rect 27488 2796 27494 2808
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 30561 2839 30619 2845
rect 30561 2805 30573 2839
rect 30607 2836 30619 2839
rect 32122 2836 32128 2848
rect 30607 2808 32128 2836
rect 30607 2805 30619 2808
rect 30561 2799 30619 2805
rect 32122 2796 32128 2808
rect 32180 2796 32186 2848
rect 34238 2796 34244 2848
rect 34296 2796 34302 2848
rect 1104 2746 35248 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 35248 2746
rect 1104 2672 35248 2694
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 4614 2632 4620 2644
rect 3283 2604 4620 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 4614 2592 4620 2604
rect 4672 2592 4678 2644
rect 4890 2592 4896 2644
rect 4948 2592 4954 2644
rect 5261 2635 5319 2641
rect 5261 2601 5273 2635
rect 5307 2632 5319 2635
rect 5442 2632 5448 2644
rect 5307 2604 5448 2632
rect 5307 2601 5319 2604
rect 5261 2595 5319 2601
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 6549 2635 6607 2641
rect 6549 2601 6561 2635
rect 6595 2632 6607 2635
rect 6730 2632 6736 2644
rect 6595 2604 6736 2632
rect 6595 2601 6607 2604
rect 6549 2595 6607 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 7006 2592 7012 2644
rect 7064 2632 7070 2644
rect 7101 2635 7159 2641
rect 7101 2632 7113 2635
rect 7064 2604 7113 2632
rect 7064 2592 7070 2604
rect 7101 2601 7113 2604
rect 7147 2601 7159 2635
rect 7101 2595 7159 2601
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 8113 2635 8171 2641
rect 8113 2632 8125 2635
rect 7248 2604 8125 2632
rect 7248 2592 7254 2604
rect 8113 2601 8125 2604
rect 8159 2601 8171 2635
rect 8113 2595 8171 2601
rect 9214 2592 9220 2644
rect 9272 2632 9278 2644
rect 9309 2635 9367 2641
rect 9309 2632 9321 2635
rect 9272 2604 9321 2632
rect 9272 2592 9278 2604
rect 9309 2601 9321 2604
rect 9355 2601 9367 2635
rect 9309 2595 9367 2601
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10137 2635 10195 2641
rect 10137 2632 10149 2635
rect 10100 2604 10149 2632
rect 10100 2592 10106 2604
rect 10137 2601 10149 2604
rect 10183 2601 10195 2635
rect 10137 2595 10195 2601
rect 11054 2592 11060 2644
rect 11112 2592 11118 2644
rect 11146 2592 11152 2644
rect 11204 2592 11210 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14185 2635 14243 2641
rect 14185 2632 14197 2635
rect 14056 2604 14197 2632
rect 14056 2592 14062 2604
rect 14185 2601 14197 2604
rect 14231 2601 14243 2635
rect 14185 2595 14243 2601
rect 14458 2592 14464 2644
rect 14516 2592 14522 2644
rect 16485 2635 16543 2641
rect 16485 2601 16497 2635
rect 16531 2632 16543 2635
rect 16758 2632 16764 2644
rect 16531 2604 16764 2632
rect 16531 2601 16543 2604
rect 16485 2595 16543 2601
rect 16758 2592 16764 2604
rect 16816 2592 16822 2644
rect 16850 2592 16856 2644
rect 16908 2592 16914 2644
rect 26421 2635 26479 2641
rect 22388 2604 26234 2632
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 4908 2564 4936 2592
rect 1627 2536 4936 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 6638 2524 6644 2576
rect 6696 2524 6702 2576
rect 6656 2496 6684 2524
rect 4448 2468 6684 2496
rect 11072 2496 11100 2592
rect 14090 2524 14096 2576
rect 14148 2524 14154 2576
rect 16574 2564 16580 2576
rect 16546 2524 16580 2564
rect 16632 2524 16638 2576
rect 16666 2524 16672 2576
rect 16724 2524 16730 2576
rect 11517 2499 11575 2505
rect 11517 2496 11529 2499
rect 11072 2468 11529 2496
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2038 2388 2044 2440
rect 2096 2388 2102 2440
rect 3050 2388 3056 2440
rect 3108 2388 3114 2440
rect 4062 2388 4068 2440
rect 4120 2388 4126 2440
rect 4448 2360 4476 2468
rect 11517 2465 11529 2468
rect 11563 2465 11575 2499
rect 11517 2459 11575 2465
rect 11790 2456 11796 2508
rect 11848 2456 11854 2508
rect 13538 2456 13544 2508
rect 13596 2456 13602 2508
rect 14108 2496 14136 2524
rect 14737 2499 14795 2505
rect 14737 2496 14749 2499
rect 14108 2468 14749 2496
rect 14737 2465 14749 2468
rect 14783 2465 14795 2499
rect 14737 2459 14795 2465
rect 15013 2499 15071 2505
rect 15013 2465 15025 2499
rect 15059 2496 15071 2499
rect 15470 2496 15476 2508
rect 15059 2468 15476 2496
rect 15059 2465 15071 2468
rect 15013 2459 15071 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 15562 2456 15568 2508
rect 15620 2496 15626 2508
rect 16546 2496 16574 2524
rect 15620 2468 16574 2496
rect 16868 2496 16896 2592
rect 17589 2499 17647 2505
rect 17589 2496 17601 2499
rect 16868 2468 17601 2496
rect 15620 2456 15626 2468
rect 4798 2388 4804 2440
rect 4856 2388 4862 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5994 2388 6000 2440
rect 6052 2428 6058 2440
rect 6365 2431 6423 2437
rect 6365 2428 6377 2431
rect 6052 2400 6377 2428
rect 6052 2388 6058 2400
rect 6365 2397 6377 2400
rect 6411 2397 6423 2431
rect 6365 2391 6423 2397
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7285 2431 7343 2437
rect 7285 2428 7297 2431
rect 7064 2400 7297 2428
rect 7064 2388 7070 2400
rect 7285 2397 7297 2400
rect 7331 2397 7343 2431
rect 7285 2391 7343 2397
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 10042 2388 10048 2440
rect 10100 2428 10106 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 10100 2400 10333 2428
rect 10100 2388 10106 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11112 2400 11345 2428
rect 11112 2388 11118 2400
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 13262 2428 13268 2440
rect 12926 2400 13268 2428
rect 11333 2391 11391 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 14090 2388 14096 2440
rect 14148 2428 14154 2440
rect 14369 2431 14427 2437
rect 14369 2428 14381 2431
rect 14148 2400 14381 2428
rect 14148 2388 14154 2400
rect 14369 2397 14381 2400
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 16132 2414 16160 2468
rect 17589 2465 17601 2468
rect 17635 2465 17647 2499
rect 17589 2459 17647 2465
rect 19061 2499 19119 2505
rect 19061 2465 19073 2499
rect 19107 2465 19119 2499
rect 19061 2459 19119 2465
rect 14645 2391 14703 2397
rect 2240 2332 4476 2360
rect 2240 2301 2268 2332
rect 2225 2295 2283 2301
rect 2225 2261 2237 2295
rect 2271 2261 2283 2295
rect 2225 2255 2283 2261
rect 4249 2295 4307 2301
rect 4249 2261 4261 2295
rect 4295 2292 4307 2295
rect 4816 2292 4844 2388
rect 14660 2360 14688 2391
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 16853 2431 16911 2437
rect 16853 2428 16865 2431
rect 16724 2400 16865 2428
rect 16724 2388 16730 2400
rect 16853 2397 16865 2400
rect 16899 2397 16911 2431
rect 16853 2391 16911 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 14918 2360 14924 2372
rect 14660 2332 14924 2360
rect 14918 2320 14924 2332
rect 14976 2320 14982 2372
rect 17328 2360 17356 2391
rect 18690 2388 18696 2440
rect 18748 2388 18754 2440
rect 19076 2428 19104 2459
rect 19334 2456 19340 2508
rect 19392 2496 19398 2508
rect 19705 2499 19763 2505
rect 19705 2496 19717 2499
rect 19392 2468 19717 2496
rect 19392 2456 19398 2468
rect 19705 2465 19717 2468
rect 19751 2465 19763 2499
rect 19705 2459 19763 2465
rect 20254 2456 20260 2508
rect 20312 2496 20318 2508
rect 22281 2499 22339 2505
rect 22281 2496 22293 2499
rect 20312 2468 22293 2496
rect 20312 2456 20318 2468
rect 22281 2465 22293 2468
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 19076 2400 19257 2428
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 21818 2388 21824 2440
rect 21876 2388 21882 2440
rect 17862 2360 17868 2372
rect 17328 2332 17868 2360
rect 17862 2320 17868 2332
rect 17920 2320 17926 2372
rect 4295 2264 4844 2292
rect 4295 2261 4307 2264
rect 4249 2255 4307 2261
rect 14366 2252 14372 2304
rect 14424 2292 14430 2304
rect 22388 2292 22416 2604
rect 26206 2564 26234 2604
rect 26421 2601 26433 2635
rect 26467 2632 26479 2635
rect 26694 2632 26700 2644
rect 26467 2604 26700 2632
rect 26467 2601 26479 2604
rect 26421 2595 26479 2601
rect 26694 2592 26700 2604
rect 26752 2592 26758 2644
rect 29273 2635 29331 2641
rect 27632 2604 29224 2632
rect 27632 2564 27660 2604
rect 26206 2536 27660 2564
rect 29196 2564 29224 2604
rect 29273 2601 29285 2635
rect 29319 2632 29331 2635
rect 31018 2632 31024 2644
rect 29319 2604 31024 2632
rect 29319 2601 29331 2604
rect 29273 2595 29331 2601
rect 31018 2592 31024 2604
rect 31076 2592 31082 2644
rect 34701 2567 34759 2573
rect 34701 2564 34713 2567
rect 29196 2536 34713 2564
rect 34701 2533 34713 2536
rect 34747 2533 34759 2567
rect 34701 2527 34759 2533
rect 23658 2456 23664 2508
rect 23716 2496 23722 2508
rect 24673 2499 24731 2505
rect 24673 2496 24685 2499
rect 23716 2468 24685 2496
rect 23716 2456 23722 2468
rect 24673 2465 24685 2468
rect 24719 2465 24731 2499
rect 24673 2459 24731 2465
rect 24946 2456 24952 2508
rect 25004 2456 25010 2508
rect 26970 2456 26976 2508
rect 27028 2496 27034 2508
rect 27522 2496 27528 2508
rect 27028 2468 27528 2496
rect 27028 2456 27034 2468
rect 27522 2456 27528 2468
rect 27580 2456 27586 2508
rect 27801 2499 27859 2505
rect 27801 2465 27813 2499
rect 27847 2496 27859 2499
rect 27890 2496 27896 2508
rect 27847 2468 27896 2496
rect 27847 2465 27859 2468
rect 27801 2459 27859 2465
rect 27890 2456 27896 2468
rect 27948 2456 27954 2508
rect 30466 2456 30472 2508
rect 30524 2496 30530 2508
rect 32585 2499 32643 2505
rect 32585 2496 32597 2499
rect 30524 2468 32597 2496
rect 30524 2456 30530 2468
rect 32585 2465 32597 2468
rect 32631 2465 32643 2499
rect 32585 2459 32643 2465
rect 34238 2456 34244 2508
rect 34296 2456 34302 2508
rect 29086 2388 29092 2440
rect 29144 2428 29150 2440
rect 29549 2431 29607 2437
rect 29549 2428 29561 2431
rect 29144 2400 29561 2428
rect 29144 2388 29150 2400
rect 29549 2397 29561 2400
rect 29595 2397 29607 2431
rect 29549 2391 29607 2397
rect 32122 2388 32128 2440
rect 32180 2388 32186 2440
rect 34514 2388 34520 2440
rect 34572 2388 34578 2440
rect 34885 2431 34943 2437
rect 34885 2397 34897 2431
rect 34931 2428 34943 2431
rect 35342 2428 35348 2440
rect 34931 2400 35348 2428
rect 34931 2397 34943 2400
rect 34885 2391 34943 2397
rect 35342 2388 35348 2400
rect 35400 2388 35406 2440
rect 25332 2332 25438 2360
rect 25332 2304 25360 2332
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 27764 2332 28290 2360
rect 27764 2320 27770 2332
rect 30374 2320 30380 2372
rect 30432 2360 30438 2372
rect 30469 2363 30527 2369
rect 30469 2360 30481 2363
rect 30432 2332 30481 2360
rect 30432 2320 30438 2332
rect 30469 2329 30481 2332
rect 30515 2329 30527 2363
rect 30469 2323 30527 2329
rect 14424 2264 22416 2292
rect 14424 2252 14430 2264
rect 25314 2252 25320 2304
rect 25372 2252 25378 2304
rect 1104 2202 35236 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 35236 2202
rect 1104 2128 35236 2150
<< via1 >>
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 18052 19320 18104 19372
rect 18236 19116 18288 19168
rect 18512 19159 18564 19168
rect 18512 19125 18521 19159
rect 18521 19125 18555 19159
rect 18555 19125 18564 19159
rect 18512 19116 18564 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 16580 18776 16632 18828
rect 18052 18819 18104 18828
rect 18052 18785 18061 18819
rect 18061 18785 18095 18819
rect 18095 18785 18104 18819
rect 18052 18776 18104 18785
rect 18512 18776 18564 18828
rect 20076 18844 20128 18896
rect 20996 18844 21048 18896
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 12716 18751 12768 18760
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 16488 18751 16540 18760
rect 16488 18717 16497 18751
rect 16497 18717 16531 18751
rect 16531 18717 16540 18751
rect 16488 18708 16540 18717
rect 18236 18751 18288 18760
rect 18236 18717 18245 18751
rect 18245 18717 18279 18751
rect 18279 18717 18288 18751
rect 18236 18708 18288 18717
rect 19984 18751 20036 18760
rect 19984 18717 19993 18751
rect 19993 18717 20027 18751
rect 20027 18717 20036 18751
rect 19984 18708 20036 18717
rect 20628 18751 20680 18760
rect 20628 18717 20637 18751
rect 20637 18717 20671 18751
rect 20671 18717 20680 18751
rect 20628 18708 20680 18717
rect 20996 18683 21048 18692
rect 20996 18649 21005 18683
rect 21005 18649 21039 18683
rect 21039 18649 21048 18683
rect 20996 18640 21048 18649
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 20352 18615 20404 18624
rect 20352 18581 20361 18615
rect 20361 18581 20395 18615
rect 20395 18581 20404 18615
rect 20352 18572 20404 18581
rect 20812 18615 20864 18624
rect 20812 18581 20821 18615
rect 20821 18581 20855 18615
rect 20855 18581 20864 18615
rect 20812 18572 20864 18581
rect 20904 18572 20956 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 12716 18368 12768 18420
rect 19984 18368 20036 18420
rect 20076 18368 20128 18420
rect 20628 18368 20680 18420
rect 11336 18232 11388 18284
rect 16580 18300 16632 18352
rect 17960 18300 18012 18352
rect 18420 18343 18472 18352
rect 18420 18309 18429 18343
rect 18429 18309 18463 18343
rect 18463 18309 18472 18343
rect 18420 18300 18472 18309
rect 14280 18232 14332 18284
rect 14832 18232 14884 18284
rect 15292 18232 15344 18284
rect 15752 18275 15804 18284
rect 15752 18241 15761 18275
rect 15761 18241 15795 18275
rect 15795 18241 15804 18275
rect 15752 18232 15804 18241
rect 11520 18164 11572 18216
rect 12624 18164 12676 18216
rect 18512 18232 18564 18284
rect 20444 18300 20496 18352
rect 20812 18300 20864 18352
rect 18328 18164 18380 18216
rect 20352 18232 20404 18284
rect 21640 18207 21692 18216
rect 21640 18173 21649 18207
rect 21649 18173 21683 18207
rect 21683 18173 21692 18207
rect 21640 18164 21692 18173
rect 13084 18071 13136 18080
rect 13084 18037 13093 18071
rect 13093 18037 13127 18071
rect 13127 18037 13136 18071
rect 13084 18028 13136 18037
rect 15200 18028 15252 18080
rect 15936 18071 15988 18080
rect 15936 18037 15945 18071
rect 15945 18037 15979 18071
rect 15979 18037 15988 18071
rect 15936 18028 15988 18037
rect 18696 18028 18748 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 14832 17867 14884 17876
rect 14832 17833 14841 17867
rect 14841 17833 14875 17867
rect 14875 17833 14884 17867
rect 14832 17824 14884 17833
rect 15936 17867 15988 17876
rect 15936 17833 15945 17867
rect 15945 17833 15979 17867
rect 15979 17833 15988 17867
rect 15936 17824 15988 17833
rect 16488 17824 16540 17876
rect 16580 17824 16632 17876
rect 15752 17756 15804 17808
rect 13084 17731 13136 17740
rect 13084 17697 13093 17731
rect 13093 17697 13127 17731
rect 13127 17697 13136 17731
rect 13084 17688 13136 17697
rect 10416 17620 10468 17672
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 11520 17663 11572 17672
rect 11520 17629 11529 17663
rect 11529 17629 11563 17663
rect 11563 17629 11572 17663
rect 11520 17620 11572 17629
rect 12072 17663 12124 17672
rect 12072 17629 12081 17663
rect 12081 17629 12115 17663
rect 12115 17629 12124 17663
rect 12072 17620 12124 17629
rect 11060 17552 11112 17604
rect 12164 17595 12216 17604
rect 12164 17561 12173 17595
rect 12173 17561 12207 17595
rect 12207 17561 12216 17595
rect 12164 17552 12216 17561
rect 10692 17484 10744 17536
rect 11520 17484 11572 17536
rect 12992 17620 13044 17672
rect 15200 17620 15252 17672
rect 15292 17620 15344 17672
rect 16396 17688 16448 17740
rect 16856 17688 16908 17740
rect 16304 17620 16356 17672
rect 16580 17663 16632 17672
rect 16580 17629 16589 17663
rect 16589 17629 16623 17663
rect 16623 17629 16632 17663
rect 16580 17620 16632 17629
rect 17960 17688 18012 17740
rect 18512 17688 18564 17740
rect 17040 17663 17092 17672
rect 17040 17629 17049 17663
rect 17049 17629 17083 17663
rect 17083 17629 17092 17663
rect 17040 17620 17092 17629
rect 17132 17620 17184 17672
rect 18328 17620 18380 17672
rect 18420 17663 18472 17672
rect 18420 17629 18429 17663
rect 18429 17629 18463 17663
rect 18463 17629 18472 17663
rect 18420 17620 18472 17629
rect 18696 17620 18748 17672
rect 18880 17731 18932 17740
rect 18880 17697 18889 17731
rect 18889 17697 18923 17731
rect 18923 17697 18932 17731
rect 18880 17688 18932 17697
rect 18972 17620 19024 17672
rect 12532 17484 12584 17536
rect 13176 17484 13228 17536
rect 13360 17527 13412 17536
rect 13360 17493 13369 17527
rect 13369 17493 13403 17527
rect 13403 17493 13412 17527
rect 13360 17484 13412 17493
rect 16028 17484 16080 17536
rect 16672 17484 16724 17536
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 18420 17484 18472 17536
rect 18972 17484 19024 17536
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 11336 17280 11388 17332
rect 12072 17280 12124 17332
rect 12164 17212 12216 17264
rect 12992 17280 13044 17332
rect 13084 17280 13136 17332
rect 15292 17280 15344 17332
rect 9956 17144 10008 17196
rect 9680 17119 9732 17128
rect 9680 17085 9689 17119
rect 9689 17085 9723 17119
rect 9723 17085 9732 17119
rect 9680 17076 9732 17085
rect 10048 17076 10100 17128
rect 12532 17187 12584 17196
rect 12532 17153 12541 17187
rect 12541 17153 12575 17187
rect 12575 17153 12584 17187
rect 12532 17144 12584 17153
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 15200 17212 15252 17264
rect 15384 17255 15436 17264
rect 15384 17221 15393 17255
rect 15393 17221 15427 17255
rect 15427 17221 15436 17255
rect 15384 17212 15436 17221
rect 15936 17280 15988 17332
rect 16304 17280 16356 17332
rect 16856 17280 16908 17332
rect 17040 17280 17092 17332
rect 16028 17144 16080 17196
rect 16672 17212 16724 17264
rect 18236 17280 18288 17332
rect 18880 17323 18932 17332
rect 18880 17289 18889 17323
rect 18889 17289 18923 17323
rect 18923 17289 18932 17323
rect 18880 17280 18932 17289
rect 19064 17280 19116 17332
rect 16488 17144 16540 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17960 17212 18012 17264
rect 17132 17076 17184 17128
rect 19984 17144 20036 17196
rect 20904 17187 20956 17196
rect 20904 17153 20913 17187
rect 20913 17153 20947 17187
rect 20947 17153 20956 17187
rect 20904 17144 20956 17153
rect 21180 17144 21232 17196
rect 18420 17008 18472 17060
rect 22100 17051 22152 17060
rect 22100 17017 22109 17051
rect 22109 17017 22143 17051
rect 22143 17017 22152 17051
rect 22100 17008 22152 17017
rect 15752 16940 15804 16992
rect 16580 16940 16632 16992
rect 16948 16940 17000 16992
rect 18512 16940 18564 16992
rect 20904 16983 20956 16992
rect 20904 16949 20913 16983
rect 20913 16949 20947 16983
rect 20947 16949 20956 16983
rect 20904 16940 20956 16949
rect 21180 16940 21232 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 10416 16736 10468 16788
rect 15752 16736 15804 16788
rect 9220 16643 9272 16652
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 14740 16668 14792 16720
rect 9772 16464 9824 16516
rect 9956 16575 10008 16584
rect 9956 16541 9965 16575
rect 9965 16541 9999 16575
rect 9999 16541 10008 16575
rect 9956 16532 10008 16541
rect 13728 16464 13780 16516
rect 14740 16532 14792 16584
rect 17684 16668 17736 16720
rect 22100 16668 22152 16720
rect 15384 16600 15436 16652
rect 16304 16600 16356 16652
rect 19248 16600 19300 16652
rect 16948 16575 17000 16584
rect 16948 16541 16957 16575
rect 16957 16541 16991 16575
rect 16991 16541 17000 16575
rect 16948 16532 17000 16541
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 22100 16575 22152 16584
rect 22100 16541 22109 16575
rect 22109 16541 22143 16575
rect 22143 16541 22152 16575
rect 22100 16532 22152 16541
rect 21364 16464 21416 16516
rect 22008 16507 22060 16516
rect 22008 16473 22017 16507
rect 22017 16473 22051 16507
rect 22051 16473 22060 16507
rect 22008 16464 22060 16473
rect 9864 16396 9916 16448
rect 10048 16396 10100 16448
rect 14464 16396 14516 16448
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 14832 16396 14884 16448
rect 15476 16396 15528 16448
rect 26056 16396 26108 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11060 16124 11112 16176
rect 13728 16167 13780 16176
rect 13728 16133 13737 16167
rect 13737 16133 13771 16167
rect 13771 16133 13780 16167
rect 13728 16124 13780 16133
rect 14280 16235 14332 16244
rect 14280 16201 14289 16235
rect 14289 16201 14323 16235
rect 14323 16201 14332 16235
rect 14280 16192 14332 16201
rect 14832 16192 14884 16244
rect 10324 16056 10376 16108
rect 10692 16056 10744 16108
rect 9772 15988 9824 16040
rect 13360 16056 13412 16108
rect 12900 16031 12952 16040
rect 12900 15997 12909 16031
rect 12909 15997 12943 16031
rect 12943 15997 12952 16031
rect 12900 15988 12952 15997
rect 13820 16031 13872 16040
rect 13820 15997 13829 16031
rect 13829 15997 13863 16031
rect 13863 15997 13872 16031
rect 13820 15988 13872 15997
rect 15476 16099 15528 16108
rect 15476 16065 15485 16099
rect 15485 16065 15519 16099
rect 15519 16065 15528 16099
rect 15476 16056 15528 16065
rect 15936 16099 15988 16108
rect 15936 16065 15945 16099
rect 15945 16065 15979 16099
rect 15979 16065 15988 16099
rect 15936 16056 15988 16065
rect 16028 16056 16080 16108
rect 17960 16099 18012 16108
rect 17960 16065 17969 16099
rect 17969 16065 18003 16099
rect 18003 16065 18012 16099
rect 17960 16056 18012 16065
rect 14648 15988 14700 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 15016 15988 15068 16040
rect 17408 16031 17460 16040
rect 17408 15997 17417 16031
rect 17417 15997 17451 16031
rect 17451 15997 17460 16031
rect 17408 15988 17460 15997
rect 18328 15988 18380 16040
rect 20996 16192 21048 16244
rect 19248 16056 19300 16108
rect 19800 16099 19852 16108
rect 19800 16065 19809 16099
rect 19809 16065 19843 16099
rect 19843 16065 19852 16099
rect 19800 16056 19852 16065
rect 11336 15852 11388 15904
rect 11428 15852 11480 15904
rect 16856 15920 16908 15972
rect 20076 16031 20128 16040
rect 20076 15997 20085 16031
rect 20085 15997 20119 16031
rect 20119 15997 20128 16031
rect 20076 15988 20128 15997
rect 20444 16056 20496 16108
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 20996 16099 21048 16108
rect 20996 16065 21005 16099
rect 21005 16065 21039 16099
rect 21039 16065 21048 16099
rect 20996 16056 21048 16065
rect 22100 16192 22152 16244
rect 22008 16124 22060 16176
rect 14372 15852 14424 15904
rect 14464 15852 14516 15904
rect 14924 15852 14976 15904
rect 19432 15895 19484 15904
rect 19432 15861 19441 15895
rect 19441 15861 19475 15895
rect 19475 15861 19484 15895
rect 19432 15852 19484 15861
rect 20720 15920 20772 15972
rect 21364 16056 21416 16108
rect 22100 16031 22152 16040
rect 22100 15997 22109 16031
rect 22109 15997 22143 16031
rect 22143 15997 22152 16031
rect 22100 15988 22152 15997
rect 26056 16167 26108 16176
rect 26056 16133 26065 16167
rect 26065 16133 26099 16167
rect 26099 16133 26108 16167
rect 26056 16124 26108 16133
rect 23296 16099 23348 16108
rect 23296 16065 23305 16099
rect 23305 16065 23339 16099
rect 23339 16065 23348 16099
rect 23296 16056 23348 16065
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 24860 16056 24912 16108
rect 26976 16124 27028 16176
rect 25688 16031 25740 16040
rect 25688 15997 25697 16031
rect 25697 15997 25731 16031
rect 25731 15997 25740 16031
rect 25688 15988 25740 15997
rect 24308 15920 24360 15972
rect 28080 16031 28132 16040
rect 28080 15997 28089 16031
rect 28089 15997 28123 16031
rect 28123 15997 28132 16031
rect 28080 15988 28132 15997
rect 26516 15895 26568 15904
rect 26516 15861 26525 15895
rect 26525 15861 26559 15895
rect 26559 15861 26568 15895
rect 26516 15852 26568 15861
rect 28172 15895 28224 15904
rect 28172 15861 28181 15895
rect 28181 15861 28215 15895
rect 28215 15861 28224 15895
rect 28172 15852 28224 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 9680 15691 9732 15700
rect 9680 15657 9689 15691
rect 9689 15657 9723 15691
rect 9723 15657 9732 15691
rect 9680 15648 9732 15657
rect 10232 15648 10284 15700
rect 10692 15623 10744 15632
rect 10692 15589 10701 15623
rect 10701 15589 10735 15623
rect 10735 15589 10744 15623
rect 10692 15580 10744 15589
rect 9956 15444 10008 15496
rect 11428 15691 11480 15700
rect 11428 15657 11437 15691
rect 11437 15657 11471 15691
rect 11471 15657 11480 15691
rect 11428 15648 11480 15657
rect 12900 15648 12952 15700
rect 13820 15648 13872 15700
rect 15016 15648 15068 15700
rect 15292 15691 15344 15700
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 17960 15648 18012 15700
rect 19800 15648 19852 15700
rect 20996 15648 21048 15700
rect 22100 15648 22152 15700
rect 23296 15648 23348 15700
rect 25688 15648 25740 15700
rect 26056 15648 26108 15700
rect 26516 15648 26568 15700
rect 11336 15512 11388 15564
rect 12164 15555 12216 15564
rect 12164 15521 12173 15555
rect 12173 15521 12207 15555
rect 12207 15521 12216 15555
rect 12164 15512 12216 15521
rect 13360 15623 13412 15632
rect 13360 15589 13369 15623
rect 13369 15589 13403 15623
rect 13403 15589 13412 15623
rect 13360 15580 13412 15589
rect 14740 15580 14792 15632
rect 11980 15487 12032 15496
rect 11980 15453 11989 15487
rect 11989 15453 12023 15487
rect 12023 15453 12032 15487
rect 11980 15444 12032 15453
rect 14464 15444 14516 15496
rect 14832 15444 14884 15496
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 9772 15376 9824 15428
rect 10416 15376 10468 15428
rect 11060 15419 11112 15428
rect 11060 15385 11069 15419
rect 11069 15385 11103 15419
rect 11103 15385 11112 15419
rect 11060 15376 11112 15385
rect 11336 15376 11388 15428
rect 14924 15419 14976 15428
rect 14924 15385 14933 15419
rect 14933 15385 14967 15419
rect 14967 15385 14976 15419
rect 14924 15376 14976 15385
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16028 15487 16080 15496
rect 16028 15453 16037 15487
rect 16037 15453 16071 15487
rect 16071 15453 16080 15487
rect 16028 15444 16080 15453
rect 16672 15444 16724 15496
rect 16764 15487 16816 15496
rect 16764 15453 16773 15487
rect 16773 15453 16807 15487
rect 16807 15453 16816 15487
rect 16764 15444 16816 15453
rect 24860 15512 24912 15564
rect 17592 15444 17644 15496
rect 20904 15444 20956 15496
rect 21180 15487 21232 15496
rect 21180 15453 21189 15487
rect 21189 15453 21223 15487
rect 21223 15453 21232 15487
rect 21180 15444 21232 15453
rect 21824 15444 21876 15496
rect 24676 15444 24728 15496
rect 28172 15648 28224 15700
rect 26976 15512 27028 15564
rect 15476 15376 15528 15428
rect 10692 15308 10744 15360
rect 12900 15308 12952 15360
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 27436 15444 27488 15496
rect 28172 15376 28224 15428
rect 27804 15351 27856 15360
rect 27804 15317 27813 15351
rect 27813 15317 27847 15351
rect 27847 15317 27856 15351
rect 27804 15308 27856 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 9496 15104 9548 15156
rect 9956 15104 10008 15156
rect 10232 15147 10284 15156
rect 10232 15113 10241 15147
rect 10241 15113 10275 15147
rect 10275 15113 10284 15147
rect 10232 15104 10284 15113
rect 9772 15036 9824 15088
rect 10416 15104 10468 15156
rect 11060 15104 11112 15156
rect 11980 15104 12032 15156
rect 17132 15147 17184 15156
rect 17132 15113 17141 15147
rect 17141 15113 17175 15147
rect 17175 15113 17184 15147
rect 17132 15104 17184 15113
rect 17408 15104 17460 15156
rect 21180 15104 21232 15156
rect 9220 14968 9272 15020
rect 9588 14968 9640 15020
rect 9680 14968 9732 15020
rect 10140 14968 10192 15020
rect 10692 14968 10744 15020
rect 11704 14968 11756 15020
rect 12072 14968 12124 15020
rect 15200 15036 15252 15088
rect 15844 15036 15896 15088
rect 20904 15036 20956 15088
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 16948 15011 17000 15020
rect 16948 14977 16957 15011
rect 16957 14977 16991 15011
rect 16991 14977 17000 15011
rect 16948 14968 17000 14977
rect 17500 15011 17552 15020
rect 12624 14900 12676 14952
rect 17500 14977 17509 15011
rect 17509 14977 17543 15011
rect 17543 14977 17552 15011
rect 17500 14968 17552 14977
rect 17592 15011 17644 15020
rect 17592 14977 17601 15011
rect 17601 14977 17635 15011
rect 17635 14977 17644 15011
rect 17592 14968 17644 14977
rect 17868 14968 17920 15020
rect 18052 14968 18104 15020
rect 20076 14968 20128 15020
rect 20720 14968 20772 15020
rect 21824 14968 21876 15020
rect 19432 14900 19484 14952
rect 9956 14832 10008 14884
rect 24860 14900 24912 14952
rect 19984 14875 20036 14884
rect 19984 14841 19993 14875
rect 19993 14841 20027 14875
rect 20027 14841 20036 14875
rect 19984 14832 20036 14841
rect 20812 14832 20864 14884
rect 23940 14832 23992 14884
rect 15292 14764 15344 14816
rect 16028 14764 16080 14816
rect 17960 14764 18012 14816
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 9772 14560 9824 14612
rect 10140 14560 10192 14612
rect 12164 14603 12216 14612
rect 12164 14569 12173 14603
rect 12173 14569 12207 14603
rect 12207 14569 12216 14603
rect 12164 14560 12216 14569
rect 14924 14560 14976 14612
rect 15660 14560 15712 14612
rect 9220 14492 9272 14544
rect 9588 14424 9640 14476
rect 9128 14399 9180 14408
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 9496 14399 9548 14408
rect 9496 14365 9505 14399
rect 9505 14365 9539 14399
rect 9539 14365 9548 14399
rect 9496 14356 9548 14365
rect 10324 14492 10376 14544
rect 11612 14492 11664 14544
rect 12072 14492 12124 14544
rect 9956 14424 10008 14476
rect 10508 14424 10560 14476
rect 12532 14492 12584 14544
rect 11612 14356 11664 14408
rect 11704 14399 11756 14408
rect 11704 14365 11713 14399
rect 11713 14365 11747 14399
rect 11747 14365 11756 14399
rect 11704 14356 11756 14365
rect 9220 14288 9272 14340
rect 9680 14220 9732 14272
rect 11060 14263 11112 14272
rect 11060 14229 11069 14263
rect 11069 14229 11103 14263
rect 11103 14229 11112 14263
rect 11060 14220 11112 14229
rect 11152 14220 11204 14272
rect 12440 14356 12492 14408
rect 12624 14424 12676 14476
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 16120 14492 16172 14544
rect 16764 14560 16816 14612
rect 17500 14603 17552 14612
rect 17500 14569 17509 14603
rect 17509 14569 17543 14603
rect 17543 14569 17552 14603
rect 17500 14560 17552 14569
rect 17868 14603 17920 14612
rect 17868 14569 17877 14603
rect 17877 14569 17911 14603
rect 17911 14569 17920 14603
rect 17868 14560 17920 14569
rect 18052 14560 18104 14612
rect 22100 14603 22152 14612
rect 14004 14356 14056 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 18144 14356 18196 14408
rect 20812 14356 20864 14408
rect 15752 14288 15804 14340
rect 11796 14220 11848 14272
rect 13636 14220 13688 14272
rect 13912 14220 13964 14272
rect 14556 14220 14608 14272
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 17960 14331 18012 14340
rect 17960 14297 17969 14331
rect 17969 14297 18003 14331
rect 18003 14297 18012 14331
rect 22100 14569 22109 14603
rect 22109 14569 22143 14603
rect 22143 14569 22152 14603
rect 22100 14560 22152 14569
rect 23664 14603 23716 14612
rect 23664 14569 23673 14603
rect 23673 14569 23707 14603
rect 23707 14569 23716 14603
rect 23664 14560 23716 14569
rect 23940 14560 23992 14612
rect 22192 14492 22244 14544
rect 21456 14424 21508 14476
rect 21548 14424 21600 14476
rect 17960 14288 18012 14297
rect 21916 14331 21968 14340
rect 23388 14424 23440 14476
rect 23020 14356 23072 14408
rect 23572 14356 23624 14408
rect 24400 14399 24452 14408
rect 24400 14365 24409 14399
rect 24409 14365 24443 14399
rect 24443 14365 24452 14399
rect 24400 14356 24452 14365
rect 24492 14399 24544 14408
rect 24492 14365 24501 14399
rect 24501 14365 24535 14399
rect 24535 14365 24544 14399
rect 24492 14356 24544 14365
rect 25044 14424 25096 14476
rect 24860 14356 24912 14408
rect 21916 14297 21951 14331
rect 21951 14297 21968 14331
rect 21916 14288 21968 14297
rect 21180 14220 21232 14272
rect 21272 14220 21324 14272
rect 22376 14288 22428 14340
rect 25320 14331 25372 14340
rect 25320 14297 25329 14331
rect 25329 14297 25363 14331
rect 25363 14297 25372 14331
rect 26056 14399 26108 14408
rect 26056 14365 26065 14399
rect 26065 14365 26099 14399
rect 26099 14365 26108 14399
rect 26056 14356 26108 14365
rect 25320 14288 25372 14297
rect 22284 14263 22336 14272
rect 22284 14229 22293 14263
rect 22293 14229 22327 14263
rect 22327 14229 22336 14263
rect 22284 14220 22336 14229
rect 23020 14220 23072 14272
rect 24124 14220 24176 14272
rect 25412 14263 25464 14272
rect 25412 14229 25421 14263
rect 25421 14229 25455 14263
rect 25455 14229 25464 14263
rect 25412 14220 25464 14229
rect 25872 14263 25924 14272
rect 25872 14229 25881 14263
rect 25881 14229 25915 14263
rect 25915 14229 25924 14263
rect 25872 14220 25924 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 9496 14016 9548 14068
rect 9680 14016 9732 14068
rect 11060 14016 11112 14068
rect 11796 14016 11848 14068
rect 12440 14016 12492 14068
rect 13268 14059 13320 14068
rect 13268 14025 13277 14059
rect 13277 14025 13311 14059
rect 13311 14025 13320 14059
rect 13268 14016 13320 14025
rect 14464 14059 14516 14068
rect 14464 14025 14473 14059
rect 14473 14025 14507 14059
rect 14507 14025 14516 14059
rect 14464 14016 14516 14025
rect 8852 13744 8904 13796
rect 9956 13812 10008 13864
rect 10324 13812 10376 13864
rect 10508 13855 10560 13864
rect 10508 13821 10517 13855
rect 10517 13821 10551 13855
rect 10551 13821 10560 13855
rect 10508 13812 10560 13821
rect 10784 13880 10836 13932
rect 13912 13948 13964 14000
rect 12440 13812 12492 13864
rect 10876 13744 10928 13796
rect 11796 13744 11848 13796
rect 12900 13855 12952 13864
rect 12900 13821 12909 13855
rect 12909 13821 12943 13855
rect 12943 13821 12952 13855
rect 13636 13855 13688 13864
rect 12900 13812 12952 13821
rect 13636 13821 13645 13855
rect 13645 13821 13679 13855
rect 13679 13821 13688 13855
rect 13636 13812 13688 13821
rect 14740 13948 14792 14000
rect 14464 13880 14516 13932
rect 14648 13880 14700 13932
rect 14924 13923 14976 13932
rect 14924 13889 14933 13923
rect 14933 13889 14967 13923
rect 14967 13889 14976 13923
rect 14924 13880 14976 13889
rect 15200 13991 15252 14000
rect 15200 13957 15209 13991
rect 15209 13957 15243 13991
rect 15243 13957 15252 13991
rect 15200 13948 15252 13957
rect 14372 13812 14424 13864
rect 16948 14016 17000 14068
rect 17684 13948 17736 14000
rect 15292 13855 15344 13864
rect 15292 13821 15301 13855
rect 15301 13821 15335 13855
rect 15335 13821 15344 13855
rect 15292 13812 15344 13821
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 20076 14016 20128 14068
rect 20812 14059 20864 14068
rect 20812 14025 20821 14059
rect 20821 14025 20855 14059
rect 20855 14025 20864 14059
rect 20812 14016 20864 14025
rect 21916 14059 21968 14068
rect 21916 14025 21925 14059
rect 21925 14025 21959 14059
rect 21959 14025 21968 14059
rect 21916 14016 21968 14025
rect 22468 14016 22520 14068
rect 23112 14016 23164 14068
rect 19340 13923 19392 13932
rect 19340 13889 19349 13923
rect 19349 13889 19383 13923
rect 19383 13889 19392 13923
rect 19340 13880 19392 13889
rect 19432 13880 19484 13932
rect 20720 13923 20772 13932
rect 20720 13889 20729 13923
rect 20729 13889 20763 13923
rect 20763 13889 20772 13923
rect 20720 13880 20772 13889
rect 19892 13812 19944 13864
rect 15936 13744 15988 13796
rect 17960 13744 18012 13796
rect 18604 13787 18656 13796
rect 18604 13753 18613 13787
rect 18613 13753 18647 13787
rect 18647 13753 18656 13787
rect 18604 13744 18656 13753
rect 18972 13744 19024 13796
rect 21272 13880 21324 13932
rect 21916 13880 21968 13932
rect 11060 13676 11112 13728
rect 14832 13676 14884 13728
rect 22100 13812 22152 13864
rect 22376 13991 22428 14000
rect 22376 13957 22385 13991
rect 22385 13957 22419 13991
rect 22419 13957 22428 13991
rect 22376 13948 22428 13957
rect 22560 13855 22612 13864
rect 22560 13821 22569 13855
rect 22569 13821 22603 13855
rect 22603 13821 22612 13855
rect 22560 13812 22612 13821
rect 23112 13880 23164 13932
rect 23664 14016 23716 14068
rect 24400 14016 24452 14068
rect 23480 13812 23532 13864
rect 24032 13880 24084 13932
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 25320 14016 25372 14068
rect 25412 14016 25464 14068
rect 25872 14016 25924 14068
rect 25228 13923 25280 13932
rect 25228 13889 25237 13923
rect 25237 13889 25271 13923
rect 25271 13889 25280 13923
rect 25228 13880 25280 13889
rect 25780 13855 25832 13864
rect 25780 13821 25789 13855
rect 25789 13821 25823 13855
rect 25823 13821 25832 13855
rect 25780 13812 25832 13821
rect 26976 13812 27028 13864
rect 21180 13719 21232 13728
rect 21180 13685 21189 13719
rect 21189 13685 21223 13719
rect 21223 13685 21232 13719
rect 21180 13676 21232 13685
rect 23296 13676 23348 13728
rect 26424 13744 26476 13796
rect 24492 13719 24544 13728
rect 24492 13685 24501 13719
rect 24501 13685 24535 13719
rect 24535 13685 24544 13719
rect 24492 13676 24544 13685
rect 24676 13676 24728 13728
rect 25412 13719 25464 13728
rect 25412 13685 25421 13719
rect 25421 13685 25455 13719
rect 25455 13685 25464 13719
rect 25412 13676 25464 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10784 13472 10836 13524
rect 11980 13472 12032 13524
rect 14832 13472 14884 13524
rect 14464 13404 14516 13456
rect 15016 13515 15068 13524
rect 15016 13481 15025 13515
rect 15025 13481 15059 13515
rect 15059 13481 15068 13515
rect 15016 13472 15068 13481
rect 23112 13472 23164 13524
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 24492 13472 24544 13524
rect 10508 13336 10560 13388
rect 9956 13268 10008 13320
rect 11060 13268 11112 13320
rect 9772 13200 9824 13252
rect 8944 13132 8996 13184
rect 10232 13132 10284 13184
rect 10968 13200 11020 13252
rect 13820 13200 13872 13252
rect 14832 13336 14884 13388
rect 14924 13336 14976 13388
rect 16304 13379 16356 13388
rect 16304 13345 16313 13379
rect 16313 13345 16347 13379
rect 16347 13345 16356 13379
rect 16304 13336 16356 13345
rect 14648 13268 14700 13320
rect 14740 13268 14792 13320
rect 15844 13268 15896 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 17316 13268 17368 13320
rect 17592 13311 17644 13320
rect 17592 13277 17601 13311
rect 17601 13277 17635 13311
rect 17635 13277 17644 13311
rect 17592 13268 17644 13277
rect 21916 13404 21968 13456
rect 18604 13379 18656 13388
rect 18604 13345 18613 13379
rect 18613 13345 18647 13379
rect 18647 13345 18656 13379
rect 18604 13336 18656 13345
rect 19984 13379 20036 13388
rect 19984 13345 19993 13379
rect 19993 13345 20027 13379
rect 20027 13345 20036 13379
rect 19984 13336 20036 13345
rect 19892 13311 19944 13320
rect 19892 13277 19901 13311
rect 19901 13277 19935 13311
rect 19935 13277 19944 13311
rect 19892 13268 19944 13277
rect 20076 13268 20128 13320
rect 21180 13268 21232 13320
rect 23388 13404 23440 13456
rect 24400 13336 24452 13388
rect 25780 13472 25832 13524
rect 26056 13472 26108 13524
rect 26976 13515 27028 13524
rect 26976 13481 26985 13515
rect 26985 13481 27019 13515
rect 27019 13481 27028 13515
rect 26976 13472 27028 13481
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 23296 13311 23348 13320
rect 23296 13277 23305 13311
rect 23305 13277 23339 13311
rect 23339 13277 23348 13311
rect 23296 13268 23348 13277
rect 24032 13268 24084 13320
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 25044 13311 25096 13320
rect 25044 13277 25053 13311
rect 25053 13277 25087 13311
rect 25087 13277 25096 13311
rect 25044 13268 25096 13277
rect 25596 13311 25648 13320
rect 25596 13277 25605 13311
rect 25605 13277 25639 13311
rect 25639 13277 25648 13311
rect 25596 13268 25648 13277
rect 15384 13243 15436 13252
rect 15384 13209 15393 13243
rect 15393 13209 15427 13243
rect 15427 13209 15436 13243
rect 15384 13200 15436 13209
rect 16764 13243 16816 13252
rect 16764 13209 16773 13243
rect 16773 13209 16807 13243
rect 16807 13209 16816 13243
rect 16764 13200 16816 13209
rect 10416 13132 10468 13184
rect 11152 13132 11204 13184
rect 11428 13132 11480 13184
rect 12256 13132 12308 13184
rect 13912 13132 13964 13184
rect 14740 13175 14792 13184
rect 14740 13141 14749 13175
rect 14749 13141 14783 13175
rect 14783 13141 14792 13175
rect 14740 13132 14792 13141
rect 14832 13132 14884 13184
rect 17684 13175 17736 13184
rect 17684 13141 17693 13175
rect 17693 13141 17727 13175
rect 17727 13141 17736 13175
rect 17684 13132 17736 13141
rect 18144 13200 18196 13252
rect 18328 13200 18380 13252
rect 18420 13243 18472 13252
rect 18420 13209 18429 13243
rect 18429 13209 18463 13243
rect 18463 13209 18472 13243
rect 18420 13200 18472 13209
rect 21272 13200 21324 13252
rect 22100 13200 22152 13252
rect 22468 13200 22520 13252
rect 24676 13200 24728 13252
rect 25228 13200 25280 13252
rect 26148 13268 26200 13320
rect 26332 13379 26384 13388
rect 26332 13345 26341 13379
rect 26341 13345 26375 13379
rect 26375 13345 26384 13379
rect 26332 13336 26384 13345
rect 18972 13132 19024 13184
rect 21180 13132 21232 13184
rect 27436 13311 27488 13320
rect 27436 13277 27445 13311
rect 27445 13277 27479 13311
rect 27479 13277 27488 13311
rect 27436 13268 27488 13277
rect 22928 13132 22980 13184
rect 23204 13132 23256 13184
rect 24124 13132 24176 13184
rect 24768 13175 24820 13184
rect 24768 13141 24777 13175
rect 24777 13141 24811 13175
rect 24811 13141 24820 13175
rect 24768 13132 24820 13141
rect 26516 13132 26568 13184
rect 26608 13175 26660 13184
rect 26608 13141 26617 13175
rect 26617 13141 26651 13175
rect 26651 13141 26660 13175
rect 26608 13132 26660 13141
rect 27804 13175 27856 13184
rect 27804 13141 27813 13175
rect 27813 13141 27847 13175
rect 27847 13141 27856 13175
rect 27804 13132 27856 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 9772 12928 9824 12980
rect 11152 12971 11204 12980
rect 11152 12937 11161 12971
rect 11161 12937 11195 12971
rect 11195 12937 11204 12971
rect 11152 12928 11204 12937
rect 9220 12903 9272 12912
rect 9220 12869 9245 12903
rect 9245 12869 9272 12903
rect 9220 12860 9272 12869
rect 8852 12792 8904 12844
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 9864 12903 9916 12912
rect 9864 12869 9873 12903
rect 9873 12869 9907 12903
rect 9907 12869 9916 12903
rect 9864 12860 9916 12869
rect 10692 12860 10744 12912
rect 10784 12792 10836 12844
rect 9956 12767 10008 12776
rect 9956 12733 9965 12767
rect 9965 12733 9999 12767
rect 9999 12733 10008 12767
rect 9956 12724 10008 12733
rect 10416 12767 10468 12776
rect 10416 12733 10425 12767
rect 10425 12733 10459 12767
rect 10459 12733 10468 12767
rect 10416 12724 10468 12733
rect 11152 12835 11204 12844
rect 11152 12801 11161 12835
rect 11161 12801 11195 12835
rect 11195 12801 11204 12835
rect 11152 12792 11204 12801
rect 11428 12792 11480 12844
rect 10048 12588 10100 12640
rect 11244 12656 11296 12708
rect 11520 12656 11572 12708
rect 11796 12792 11848 12844
rect 11888 12699 11940 12708
rect 11888 12665 11897 12699
rect 11897 12665 11931 12699
rect 11931 12665 11940 12699
rect 11888 12656 11940 12665
rect 11980 12656 12032 12708
rect 12256 12835 12308 12844
rect 12256 12801 12265 12835
rect 12265 12801 12299 12835
rect 12299 12801 12308 12835
rect 12256 12792 12308 12801
rect 14372 12792 14424 12844
rect 15200 12928 15252 12980
rect 15384 12928 15436 12980
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 16672 12971 16724 12980
rect 16672 12937 16681 12971
rect 16681 12937 16715 12971
rect 16715 12937 16724 12971
rect 16672 12928 16724 12937
rect 19984 12928 20036 12980
rect 26608 12928 26660 12980
rect 26792 12971 26844 12980
rect 26792 12937 26801 12971
rect 26801 12937 26835 12971
rect 26835 12937 26844 12971
rect 26792 12928 26844 12937
rect 27436 12928 27488 12980
rect 17592 12860 17644 12912
rect 19340 12860 19392 12912
rect 22284 12860 22336 12912
rect 15844 12835 15896 12844
rect 15844 12801 15853 12835
rect 15853 12801 15887 12835
rect 15887 12801 15896 12835
rect 15844 12792 15896 12801
rect 15936 12792 15988 12844
rect 15200 12767 15252 12776
rect 15200 12733 15209 12767
rect 15209 12733 15243 12767
rect 15243 12733 15252 12767
rect 15200 12724 15252 12733
rect 14740 12656 14792 12708
rect 15016 12699 15068 12708
rect 15016 12665 15025 12699
rect 15025 12665 15059 12699
rect 15059 12665 15068 12699
rect 15016 12656 15068 12665
rect 15476 12656 15528 12708
rect 16856 12724 16908 12776
rect 17224 12835 17276 12844
rect 17224 12801 17233 12835
rect 17233 12801 17267 12835
rect 17267 12801 17276 12835
rect 17224 12792 17276 12801
rect 17316 12792 17368 12844
rect 18972 12835 19024 12844
rect 18972 12801 18981 12835
rect 18981 12801 19015 12835
rect 19015 12801 19024 12835
rect 18972 12792 19024 12801
rect 26516 12835 26568 12844
rect 17960 12724 18012 12776
rect 21916 12724 21968 12776
rect 26516 12801 26525 12835
rect 26525 12801 26559 12835
rect 26559 12801 26568 12835
rect 26516 12792 26568 12801
rect 28080 12792 28132 12844
rect 28356 12792 28408 12844
rect 27804 12767 27856 12776
rect 27804 12733 27813 12767
rect 27813 12733 27847 12767
rect 27847 12733 27856 12767
rect 27804 12724 27856 12733
rect 16672 12656 16724 12708
rect 19432 12656 19484 12708
rect 22192 12699 22244 12708
rect 22192 12665 22201 12699
rect 22201 12665 22235 12699
rect 22235 12665 22244 12699
rect 22192 12656 22244 12665
rect 16580 12588 16632 12640
rect 19340 12588 19392 12640
rect 22652 12588 22704 12640
rect 26976 12588 27028 12640
rect 28540 12588 28592 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 9312 12427 9364 12436
rect 9312 12393 9321 12427
rect 9321 12393 9355 12427
rect 9355 12393 9364 12427
rect 9312 12384 9364 12393
rect 10784 12384 10836 12436
rect 11244 12427 11296 12436
rect 11244 12393 11253 12427
rect 11253 12393 11287 12427
rect 11287 12393 11296 12427
rect 11244 12384 11296 12393
rect 11888 12384 11940 12436
rect 12256 12384 12308 12436
rect 15108 12384 15160 12436
rect 9864 12316 9916 12368
rect 11060 12316 11112 12368
rect 11612 12316 11664 12368
rect 11796 12316 11848 12368
rect 9588 12291 9640 12300
rect 9588 12257 9597 12291
rect 9597 12257 9631 12291
rect 9631 12257 9640 12291
rect 9588 12248 9640 12257
rect 9312 12180 9364 12232
rect 9772 12180 9824 12232
rect 10416 12180 10468 12232
rect 11060 12223 11112 12232
rect 11060 12189 11069 12223
rect 11069 12189 11103 12223
rect 11103 12189 11112 12223
rect 11060 12180 11112 12189
rect 11244 12180 11296 12232
rect 11428 12180 11480 12232
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 9404 12044 9456 12096
rect 9864 12044 9916 12096
rect 10232 12044 10284 12096
rect 11980 12180 12032 12232
rect 11244 12044 11296 12096
rect 14464 12248 14516 12300
rect 12348 12180 12400 12232
rect 13360 12180 13412 12232
rect 13820 12180 13872 12232
rect 14188 12112 14240 12164
rect 14372 12155 14424 12164
rect 14372 12121 14381 12155
rect 14381 12121 14415 12155
rect 14415 12121 14424 12155
rect 14372 12112 14424 12121
rect 15476 12316 15528 12368
rect 15844 12316 15896 12368
rect 16028 12291 16080 12300
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 15016 12180 15068 12232
rect 16028 12257 16037 12291
rect 16037 12257 16071 12291
rect 16071 12257 16080 12291
rect 16028 12248 16080 12257
rect 16212 12223 16264 12232
rect 16212 12189 16221 12223
rect 16221 12189 16255 12223
rect 16255 12189 16264 12223
rect 16212 12180 16264 12189
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 16764 12384 16816 12436
rect 20076 12384 20128 12436
rect 22284 12427 22336 12436
rect 22284 12393 22293 12427
rect 22293 12393 22327 12427
rect 22327 12393 22336 12427
rect 22284 12384 22336 12393
rect 25780 12427 25832 12436
rect 25780 12393 25789 12427
rect 25789 12393 25823 12427
rect 25823 12393 25832 12427
rect 25780 12384 25832 12393
rect 26332 12384 26384 12436
rect 16580 12316 16632 12368
rect 16396 12180 16448 12232
rect 16672 12223 16724 12232
rect 16672 12189 16681 12223
rect 16681 12189 16715 12223
rect 16715 12189 16724 12223
rect 16672 12180 16724 12189
rect 16856 12180 16908 12232
rect 16948 12223 17000 12232
rect 16948 12189 16957 12223
rect 16957 12189 16991 12223
rect 16991 12189 17000 12223
rect 16948 12180 17000 12189
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 15844 12112 15896 12164
rect 16580 12112 16632 12164
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 18788 12223 18840 12232
rect 18788 12189 18797 12223
rect 18797 12189 18831 12223
rect 18831 12189 18840 12223
rect 18788 12180 18840 12189
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 18696 12112 18748 12164
rect 17592 12087 17644 12096
rect 17592 12053 17601 12087
rect 17601 12053 17635 12087
rect 17635 12053 17644 12087
rect 19432 12180 19484 12232
rect 17592 12044 17644 12053
rect 22192 12180 22244 12232
rect 22652 12223 22704 12232
rect 22652 12189 22661 12223
rect 22661 12189 22695 12223
rect 22695 12189 22704 12223
rect 22652 12180 22704 12189
rect 23204 12248 23256 12300
rect 23112 12180 23164 12232
rect 22560 12112 22612 12164
rect 24308 12180 24360 12232
rect 24768 12223 24820 12232
rect 24768 12189 24777 12223
rect 24777 12189 24811 12223
rect 24811 12189 24820 12223
rect 24768 12180 24820 12189
rect 25504 12180 25556 12232
rect 26148 12223 26200 12232
rect 26148 12189 26157 12223
rect 26157 12189 26191 12223
rect 26191 12189 26200 12223
rect 26148 12180 26200 12189
rect 26332 12223 26384 12232
rect 26332 12189 26341 12223
rect 26341 12189 26375 12223
rect 26375 12189 26384 12223
rect 26332 12180 26384 12189
rect 27804 12180 27856 12232
rect 28264 12316 28316 12368
rect 28080 12180 28132 12232
rect 28356 12180 28408 12232
rect 19984 12044 20036 12096
rect 23572 12044 23624 12096
rect 24308 12044 24360 12096
rect 24584 12044 24636 12096
rect 24860 12087 24912 12096
rect 24860 12053 24869 12087
rect 24869 12053 24903 12087
rect 24903 12053 24912 12087
rect 24860 12044 24912 12053
rect 25596 12044 25648 12096
rect 27712 12087 27764 12096
rect 27712 12053 27721 12087
rect 27721 12053 27755 12087
rect 27755 12053 27764 12087
rect 27712 12044 27764 12053
rect 27896 12044 27948 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 9220 11840 9272 11892
rect 9588 11840 9640 11892
rect 11152 11840 11204 11892
rect 9404 11636 9456 11688
rect 9772 11747 9824 11756
rect 9772 11713 9781 11747
rect 9781 11713 9815 11747
rect 9815 11713 9824 11747
rect 9772 11704 9824 11713
rect 9956 11747 10008 11756
rect 9956 11713 9965 11747
rect 9965 11713 9999 11747
rect 9999 11713 10008 11747
rect 9956 11704 10008 11713
rect 10784 11704 10836 11756
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 11060 11704 11112 11756
rect 11244 11704 11296 11756
rect 14188 11840 14240 11892
rect 17408 11840 17460 11892
rect 17592 11840 17644 11892
rect 18696 11840 18748 11892
rect 18788 11840 18840 11892
rect 19984 11840 20036 11892
rect 11612 11679 11664 11688
rect 11612 11645 11621 11679
rect 11621 11645 11655 11679
rect 11655 11645 11664 11679
rect 11612 11636 11664 11645
rect 12164 11704 12216 11756
rect 13360 11636 13412 11688
rect 13820 11679 13872 11688
rect 13820 11645 13829 11679
rect 13829 11645 13863 11679
rect 13863 11645 13872 11679
rect 13820 11636 13872 11645
rect 9312 11500 9364 11552
rect 10232 11500 10284 11552
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 11704 11500 11756 11552
rect 12624 11500 12676 11552
rect 13636 11500 13688 11552
rect 14464 11704 14516 11756
rect 16028 11772 16080 11824
rect 16304 11704 16356 11756
rect 23112 11840 23164 11892
rect 23204 11840 23256 11892
rect 23572 11840 23624 11892
rect 24860 11840 24912 11892
rect 26332 11840 26384 11892
rect 15108 11636 15160 11688
rect 18420 11636 18472 11688
rect 21640 11704 21692 11756
rect 22560 11747 22612 11756
rect 22560 11713 22569 11747
rect 22569 11713 22603 11747
rect 22603 11713 22612 11747
rect 22560 11704 22612 11713
rect 18880 11636 18932 11688
rect 21732 11636 21784 11688
rect 24584 11704 24636 11756
rect 25136 11704 25188 11756
rect 25504 11704 25556 11756
rect 25596 11704 25648 11756
rect 28080 11840 28132 11892
rect 28172 11840 28224 11892
rect 28264 11840 28316 11892
rect 27896 11747 27948 11756
rect 27896 11713 27905 11747
rect 27905 11713 27939 11747
rect 27939 11713 27948 11747
rect 27896 11704 27948 11713
rect 25320 11679 25372 11688
rect 25320 11645 25329 11679
rect 25329 11645 25363 11679
rect 25363 11645 25372 11679
rect 25320 11636 25372 11645
rect 26056 11679 26108 11688
rect 26056 11645 26065 11679
rect 26065 11645 26099 11679
rect 26099 11645 26108 11679
rect 26056 11636 26108 11645
rect 28540 11679 28592 11688
rect 28540 11645 28549 11679
rect 28549 11645 28583 11679
rect 28583 11645 28592 11679
rect 28540 11636 28592 11645
rect 28080 11568 28132 11620
rect 14188 11500 14240 11552
rect 14832 11500 14884 11552
rect 15200 11500 15252 11552
rect 16856 11543 16908 11552
rect 16856 11509 16865 11543
rect 16865 11509 16899 11543
rect 16899 11509 16908 11543
rect 16856 11500 16908 11509
rect 19524 11500 19576 11552
rect 19616 11500 19668 11552
rect 20076 11500 20128 11552
rect 20812 11543 20864 11552
rect 20812 11509 20821 11543
rect 20821 11509 20855 11543
rect 20855 11509 20864 11543
rect 20812 11500 20864 11509
rect 22468 11500 22520 11552
rect 23756 11500 23808 11552
rect 27804 11500 27856 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 11060 11296 11112 11348
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 12164 11296 12216 11348
rect 11520 11228 11572 11280
rect 15016 11296 15068 11348
rect 16396 11339 16448 11348
rect 16396 11305 16405 11339
rect 16405 11305 16439 11339
rect 16439 11305 16448 11339
rect 16396 11296 16448 11305
rect 19432 11296 19484 11348
rect 19616 11339 19668 11348
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 24860 11296 24912 11348
rect 25136 11296 25188 11348
rect 9312 11135 9364 11144
rect 9312 11101 9321 11135
rect 9321 11101 9355 11135
rect 9355 11101 9364 11135
rect 9312 11092 9364 11101
rect 9772 11135 9824 11144
rect 9772 11101 9781 11135
rect 9781 11101 9815 11135
rect 9815 11101 9824 11135
rect 9772 11092 9824 11101
rect 10232 11092 10284 11144
rect 11612 11160 11664 11212
rect 12072 11160 12124 11212
rect 12716 11203 12768 11212
rect 12716 11169 12725 11203
rect 12725 11169 12759 11203
rect 12759 11169 12768 11203
rect 12716 11160 12768 11169
rect 14648 11160 14700 11212
rect 15476 11160 15528 11212
rect 15568 11203 15620 11212
rect 15568 11169 15577 11203
rect 15577 11169 15611 11203
rect 15611 11169 15620 11203
rect 15568 11160 15620 11169
rect 10324 11024 10376 11076
rect 11060 11067 11112 11076
rect 11060 11033 11069 11067
rect 11069 11033 11103 11067
rect 11103 11033 11112 11067
rect 11060 11024 11112 11033
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 13360 11092 13412 11144
rect 14832 11135 14884 11144
rect 14832 11101 14841 11135
rect 14841 11101 14875 11135
rect 14875 11101 14884 11135
rect 14832 11092 14884 11101
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 15200 11092 15252 11101
rect 9404 10956 9456 11008
rect 14832 10956 14884 11008
rect 16120 11160 16172 11212
rect 19524 11228 19576 11280
rect 20444 11228 20496 11280
rect 25320 11339 25372 11348
rect 25320 11305 25329 11339
rect 25329 11305 25363 11339
rect 25363 11305 25372 11339
rect 25320 11296 25372 11305
rect 26148 11296 26200 11348
rect 27436 11339 27488 11348
rect 27436 11305 27445 11339
rect 27445 11305 27479 11339
rect 27479 11305 27488 11339
rect 27436 11296 27488 11305
rect 27712 11296 27764 11348
rect 16304 11092 16356 11144
rect 18512 11092 18564 11144
rect 19524 11135 19576 11144
rect 19524 11101 19533 11135
rect 19533 11101 19567 11135
rect 19567 11101 19576 11135
rect 19524 11092 19576 11101
rect 25504 11092 25556 11144
rect 25596 11135 25648 11144
rect 25596 11101 25605 11135
rect 25605 11101 25639 11135
rect 25639 11101 25648 11135
rect 25596 11092 25648 11101
rect 16672 11067 16724 11076
rect 16672 11033 16681 11067
rect 16681 11033 16715 11067
rect 16715 11033 16724 11067
rect 16672 11024 16724 11033
rect 25320 11024 25372 11076
rect 27988 11067 28040 11076
rect 27988 11033 27997 11067
rect 27997 11033 28031 11067
rect 28031 11033 28040 11067
rect 27988 11024 28040 11033
rect 28172 11067 28224 11076
rect 28172 11033 28181 11067
rect 28181 11033 28215 11067
rect 28215 11033 28224 11067
rect 28172 11024 28224 11033
rect 15752 10956 15804 11008
rect 16028 10956 16080 11008
rect 16212 10999 16264 11008
rect 16212 10965 16221 10999
rect 16221 10965 16255 10999
rect 16255 10965 16264 10999
rect 16212 10956 16264 10965
rect 25504 10956 25556 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 13728 10752 13780 10804
rect 16212 10752 16264 10804
rect 21640 10795 21692 10804
rect 21640 10761 21649 10795
rect 21649 10761 21683 10795
rect 21683 10761 21692 10795
rect 21640 10752 21692 10761
rect 21824 10795 21876 10804
rect 21824 10761 21833 10795
rect 21833 10761 21867 10795
rect 21867 10761 21876 10795
rect 21824 10752 21876 10761
rect 23296 10752 23348 10804
rect 25320 10752 25372 10804
rect 11244 10684 11296 10736
rect 14372 10684 14424 10736
rect 10416 10659 10468 10668
rect 10416 10625 10425 10659
rect 10425 10625 10459 10659
rect 10459 10625 10468 10659
rect 10416 10616 10468 10625
rect 10784 10616 10836 10668
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 14004 10616 14056 10668
rect 13452 10480 13504 10532
rect 13912 10480 13964 10532
rect 16028 10727 16080 10736
rect 16028 10693 16037 10727
rect 16037 10693 16071 10727
rect 16071 10693 16080 10727
rect 16028 10684 16080 10693
rect 14832 10659 14884 10668
rect 14832 10625 14841 10659
rect 14841 10625 14875 10659
rect 14875 10625 14884 10659
rect 14832 10616 14884 10625
rect 9404 10412 9456 10464
rect 11336 10412 11388 10464
rect 12164 10412 12216 10464
rect 15384 10548 15436 10600
rect 15660 10480 15712 10532
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 21456 10659 21508 10668
rect 21456 10625 21465 10659
rect 21465 10625 21499 10659
rect 21499 10625 21508 10659
rect 21456 10616 21508 10625
rect 22100 10659 22152 10668
rect 22100 10625 22109 10659
rect 22109 10625 22143 10659
rect 22143 10625 22152 10659
rect 22100 10616 22152 10625
rect 17684 10480 17736 10532
rect 21916 10548 21968 10600
rect 22468 10659 22520 10668
rect 22468 10625 22477 10659
rect 22477 10625 22511 10659
rect 22511 10625 22520 10659
rect 22468 10616 22520 10625
rect 22928 10616 22980 10668
rect 26424 10616 26476 10668
rect 26792 10616 26844 10668
rect 23848 10548 23900 10600
rect 24676 10548 24728 10600
rect 23940 10480 23992 10532
rect 24032 10480 24084 10532
rect 16120 10412 16172 10464
rect 16396 10455 16448 10464
rect 16396 10421 16405 10455
rect 16405 10421 16439 10455
rect 16439 10421 16448 10455
rect 16396 10412 16448 10421
rect 17776 10412 17828 10464
rect 19892 10412 19944 10464
rect 21272 10412 21324 10464
rect 23572 10412 23624 10464
rect 26516 10455 26568 10464
rect 26516 10421 26525 10455
rect 26525 10421 26559 10455
rect 26559 10421 26568 10455
rect 26516 10412 26568 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 14556 10208 14608 10260
rect 15384 10208 15436 10260
rect 16028 10208 16080 10260
rect 17316 10208 17368 10260
rect 18328 10251 18380 10260
rect 18328 10217 18337 10251
rect 18337 10217 18371 10251
rect 18371 10217 18380 10251
rect 18328 10208 18380 10217
rect 21272 10208 21324 10260
rect 7748 10047 7800 10056
rect 7748 10013 7757 10047
rect 7757 10013 7791 10047
rect 7791 10013 7800 10047
rect 7748 10004 7800 10013
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 11060 10004 11112 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11888 10004 11940 10056
rect 12440 10004 12492 10056
rect 13544 10072 13596 10124
rect 13728 10140 13780 10192
rect 14280 10072 14332 10124
rect 9404 9868 9456 9920
rect 13452 9936 13504 9988
rect 14188 10004 14240 10056
rect 15660 10072 15712 10124
rect 11796 9868 11848 9920
rect 14372 9979 14424 9988
rect 14372 9945 14381 9979
rect 14381 9945 14415 9979
rect 14415 9945 14424 9979
rect 14924 10004 14976 10056
rect 16028 10004 16080 10056
rect 16120 10047 16172 10056
rect 16120 10013 16129 10047
rect 16129 10013 16163 10047
rect 16163 10013 16172 10047
rect 16120 10004 16172 10013
rect 16212 10004 16264 10056
rect 16304 10047 16356 10056
rect 16304 10013 16313 10047
rect 16313 10013 16347 10047
rect 16347 10013 16356 10047
rect 16304 10004 16356 10013
rect 19340 10140 19392 10192
rect 21456 10140 21508 10192
rect 17776 10004 17828 10056
rect 18236 10072 18288 10124
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 14372 9936 14424 9945
rect 18052 9936 18104 9988
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 20536 10047 20588 10056
rect 20536 10013 20545 10047
rect 20545 10013 20579 10047
rect 20579 10013 20588 10047
rect 20536 10004 20588 10013
rect 22928 10208 22980 10260
rect 23848 10251 23900 10260
rect 23848 10217 23857 10251
rect 23857 10217 23891 10251
rect 23891 10217 23900 10251
rect 23848 10208 23900 10217
rect 24124 10251 24176 10260
rect 24124 10217 24133 10251
rect 24133 10217 24167 10251
rect 24167 10217 24176 10251
rect 24124 10208 24176 10217
rect 25504 10208 25556 10260
rect 22100 10140 22152 10192
rect 23296 10140 23348 10192
rect 23572 10115 23624 10124
rect 23572 10081 23581 10115
rect 23581 10081 23615 10115
rect 23615 10081 23624 10115
rect 23572 10072 23624 10081
rect 17592 9868 17644 9920
rect 20260 9936 20312 9988
rect 21916 10047 21968 10056
rect 21916 10013 21944 10047
rect 21944 10013 21968 10047
rect 21916 10004 21968 10013
rect 22100 10047 22152 10056
rect 22100 10013 22106 10047
rect 22106 10013 22140 10047
rect 22140 10013 22152 10047
rect 26792 10115 26844 10124
rect 26792 10081 26801 10115
rect 26801 10081 26835 10115
rect 26835 10081 26844 10115
rect 26792 10072 26844 10081
rect 22100 10004 22152 10013
rect 23940 10004 23992 10056
rect 24492 10047 24544 10056
rect 24492 10013 24501 10047
rect 24501 10013 24535 10047
rect 24535 10013 24544 10047
rect 24492 10004 24544 10013
rect 24584 10047 24636 10056
rect 24584 10013 24593 10047
rect 24593 10013 24627 10047
rect 24627 10013 24636 10047
rect 24584 10004 24636 10013
rect 24860 10004 24912 10056
rect 24952 10047 25004 10056
rect 24952 10013 24961 10047
rect 24961 10013 24995 10047
rect 24995 10013 25004 10047
rect 24952 10004 25004 10013
rect 23296 9936 23348 9988
rect 26424 10004 26476 10056
rect 26516 9936 26568 9988
rect 18880 9911 18932 9920
rect 18880 9877 18889 9911
rect 18889 9877 18923 9911
rect 18923 9877 18932 9911
rect 18880 9868 18932 9877
rect 19892 9868 19944 9920
rect 21364 9868 21416 9920
rect 22100 9868 22152 9920
rect 22284 9911 22336 9920
rect 22284 9877 22293 9911
rect 22293 9877 22327 9911
rect 22327 9877 22336 9911
rect 22284 9868 22336 9877
rect 22744 9911 22796 9920
rect 22744 9877 22753 9911
rect 22753 9877 22787 9911
rect 22787 9877 22796 9911
rect 22744 9868 22796 9877
rect 25504 9868 25556 9920
rect 27344 9911 27396 9920
rect 27344 9877 27353 9911
rect 27353 9877 27387 9911
rect 27387 9877 27396 9911
rect 27344 9868 27396 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 10876 9664 10928 9716
rect 15844 9664 15896 9716
rect 8760 9571 8812 9580
rect 8760 9537 8769 9571
rect 8769 9537 8803 9571
rect 8803 9537 8812 9571
rect 8760 9528 8812 9537
rect 9220 9571 9272 9580
rect 9220 9537 9229 9571
rect 9229 9537 9263 9571
rect 9263 9537 9272 9571
rect 9220 9528 9272 9537
rect 11704 9596 11756 9648
rect 10968 9528 11020 9580
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 15568 9596 15620 9648
rect 17592 9596 17644 9648
rect 15384 9528 15436 9580
rect 18328 9664 18380 9716
rect 20536 9707 20588 9716
rect 20536 9673 20545 9707
rect 20545 9673 20579 9707
rect 20579 9673 20588 9707
rect 20536 9664 20588 9673
rect 21916 9664 21968 9716
rect 22284 9664 22336 9716
rect 22744 9664 22796 9716
rect 21180 9639 21232 9648
rect 21180 9605 21189 9639
rect 21189 9605 21223 9639
rect 21223 9605 21232 9639
rect 21180 9596 21232 9605
rect 15844 9460 15896 9512
rect 16672 9460 16724 9512
rect 17868 9460 17920 9512
rect 18512 9528 18564 9580
rect 19340 9528 19392 9580
rect 20536 9528 20588 9580
rect 23020 9639 23072 9648
rect 23020 9605 23029 9639
rect 23029 9605 23063 9639
rect 23063 9605 23072 9639
rect 23020 9596 23072 9605
rect 12440 9392 12492 9444
rect 15752 9324 15804 9376
rect 17960 9324 18012 9376
rect 19984 9460 20036 9512
rect 20996 9460 21048 9512
rect 24584 9664 24636 9716
rect 24492 9596 24544 9648
rect 23480 9503 23532 9512
rect 23480 9469 23489 9503
rect 23489 9469 23523 9503
rect 23523 9469 23532 9503
rect 23480 9460 23532 9469
rect 23848 9571 23900 9580
rect 23848 9537 23857 9571
rect 23857 9537 23891 9571
rect 23891 9537 23900 9571
rect 23848 9528 23900 9537
rect 23940 9528 23992 9580
rect 24216 9528 24268 9580
rect 24676 9528 24728 9580
rect 26516 9596 26568 9648
rect 25504 9460 25556 9512
rect 24124 9392 24176 9444
rect 25412 9392 25464 9444
rect 26976 9528 27028 9580
rect 27344 9460 27396 9512
rect 27528 9503 27580 9512
rect 27528 9469 27537 9503
rect 27537 9469 27571 9503
rect 27571 9469 27580 9503
rect 27528 9460 27580 9469
rect 19432 9324 19484 9376
rect 22468 9324 22520 9376
rect 23388 9324 23440 9376
rect 23848 9324 23900 9376
rect 24860 9324 24912 9376
rect 25228 9367 25280 9376
rect 25228 9333 25237 9367
rect 25237 9333 25271 9367
rect 25271 9333 25280 9367
rect 25228 9324 25280 9333
rect 25780 9367 25832 9376
rect 25780 9333 25789 9367
rect 25789 9333 25823 9367
rect 25823 9333 25832 9367
rect 25780 9324 25832 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 15752 9120 15804 9172
rect 15844 9163 15896 9172
rect 15844 9129 15853 9163
rect 15853 9129 15887 9163
rect 15887 9129 15896 9163
rect 15844 9120 15896 9129
rect 14280 9052 14332 9104
rect 14740 9052 14792 9104
rect 10232 8959 10284 8968
rect 10232 8925 10241 8959
rect 10241 8925 10275 8959
rect 10275 8925 10284 8959
rect 10232 8916 10284 8925
rect 10324 8916 10376 8968
rect 14832 8984 14884 9036
rect 15016 9027 15068 9036
rect 15016 8993 15025 9027
rect 15025 8993 15059 9027
rect 15059 8993 15068 9027
rect 15016 8984 15068 8993
rect 14188 8848 14240 8900
rect 14556 8959 14608 8968
rect 14556 8925 14565 8959
rect 14565 8925 14599 8959
rect 14599 8925 14608 8959
rect 14556 8916 14608 8925
rect 15200 8848 15252 8900
rect 14556 8780 14608 8832
rect 14648 8823 14700 8832
rect 14648 8789 14657 8823
rect 14657 8789 14691 8823
rect 14691 8789 14700 8823
rect 14648 8780 14700 8789
rect 14740 8780 14792 8832
rect 15660 8916 15712 8968
rect 16304 8916 16356 8968
rect 21364 9120 21416 9172
rect 23480 9120 23532 9172
rect 24124 9120 24176 9172
rect 24952 9163 25004 9172
rect 24952 9129 24961 9163
rect 24961 9129 24995 9163
rect 24995 9129 25004 9163
rect 24952 9120 25004 9129
rect 25780 9120 25832 9172
rect 27620 9120 27672 9172
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 21180 9052 21232 9104
rect 23664 9052 23716 9104
rect 24676 8984 24728 9036
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 21180 8916 21232 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 21916 8916 21968 8968
rect 24216 8916 24268 8968
rect 24492 8916 24544 8968
rect 17592 8891 17644 8900
rect 17592 8857 17601 8891
rect 17601 8857 17635 8891
rect 17635 8857 17644 8891
rect 17592 8848 17644 8857
rect 25228 8959 25280 8968
rect 25228 8925 25237 8959
rect 25237 8925 25271 8959
rect 25271 8925 25280 8959
rect 25228 8916 25280 8925
rect 27712 9052 27764 9104
rect 27988 9052 28040 9104
rect 27896 8959 27948 8968
rect 27896 8925 27905 8959
rect 27905 8925 27939 8959
rect 27939 8925 27948 8959
rect 27896 8916 27948 8925
rect 16764 8780 16816 8832
rect 16856 8780 16908 8832
rect 21180 8780 21232 8832
rect 27804 8848 27856 8900
rect 22192 8823 22244 8832
rect 22192 8789 22201 8823
rect 22201 8789 22235 8823
rect 22235 8789 22244 8823
rect 22192 8780 22244 8789
rect 23940 8780 23992 8832
rect 24584 8780 24636 8832
rect 25872 8780 25924 8832
rect 27988 8780 28040 8832
rect 28908 8823 28960 8832
rect 28908 8789 28917 8823
rect 28917 8789 28951 8823
rect 28951 8789 28960 8823
rect 28908 8780 28960 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 10232 8576 10284 8628
rect 7748 8508 7800 8560
rect 7288 8483 7340 8492
rect 7288 8449 7297 8483
rect 7297 8449 7331 8483
rect 7331 8449 7340 8483
rect 7288 8440 7340 8449
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 9220 8508 9272 8560
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 11980 8576 12032 8628
rect 10140 8415 10192 8424
rect 10140 8381 10149 8415
rect 10149 8381 10183 8415
rect 10183 8381 10192 8415
rect 10140 8372 10192 8381
rect 10876 8415 10928 8424
rect 10876 8381 10885 8415
rect 10885 8381 10919 8415
rect 10919 8381 10928 8415
rect 10876 8372 10928 8381
rect 11060 8440 11112 8492
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 12072 8508 12124 8560
rect 14648 8576 14700 8628
rect 14740 8619 14792 8628
rect 14740 8585 14749 8619
rect 14749 8585 14783 8619
rect 14783 8585 14792 8619
rect 14740 8576 14792 8585
rect 15384 8619 15436 8628
rect 15384 8585 15393 8619
rect 15393 8585 15427 8619
rect 15427 8585 15436 8619
rect 15384 8576 15436 8585
rect 15568 8576 15620 8628
rect 18880 8576 18932 8628
rect 19984 8576 20036 8628
rect 23664 8619 23716 8628
rect 23664 8585 23673 8619
rect 23673 8585 23707 8619
rect 23707 8585 23716 8619
rect 23664 8576 23716 8585
rect 9128 8304 9180 8356
rect 8852 8236 8904 8288
rect 9588 8304 9640 8356
rect 10232 8304 10284 8356
rect 12532 8440 12584 8492
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 14188 8440 14240 8492
rect 17500 8551 17552 8560
rect 17500 8517 17509 8551
rect 17509 8517 17543 8551
rect 17543 8517 17552 8551
rect 17500 8508 17552 8517
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 16856 8440 16908 8492
rect 18696 8483 18748 8492
rect 18696 8449 18705 8483
rect 18705 8449 18739 8483
rect 18739 8449 18748 8483
rect 18696 8440 18748 8449
rect 18880 8483 18932 8492
rect 18880 8449 18889 8483
rect 18889 8449 18923 8483
rect 18923 8449 18932 8483
rect 18880 8440 18932 8449
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 23572 8440 23624 8492
rect 23940 8440 23992 8492
rect 26516 8551 26568 8560
rect 26516 8517 26525 8551
rect 26525 8517 26559 8551
rect 26559 8517 26568 8551
rect 26516 8508 26568 8517
rect 26976 8551 27028 8560
rect 24860 8440 24912 8492
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25780 8440 25832 8492
rect 26976 8517 26985 8551
rect 26985 8517 27019 8551
rect 27019 8517 27028 8551
rect 26976 8508 27028 8517
rect 27068 8508 27120 8560
rect 27620 8576 27672 8628
rect 27896 8576 27948 8628
rect 27344 8440 27396 8492
rect 11980 8304 12032 8356
rect 12348 8304 12400 8356
rect 15108 8415 15160 8424
rect 15108 8381 15117 8415
rect 15117 8381 15151 8415
rect 15151 8381 15160 8415
rect 15108 8372 15160 8381
rect 15660 8372 15712 8424
rect 19984 8372 20036 8424
rect 20168 8415 20220 8424
rect 20168 8381 20177 8415
rect 20177 8381 20211 8415
rect 20211 8381 20220 8415
rect 20168 8372 20220 8381
rect 24952 8372 25004 8424
rect 27712 8483 27764 8492
rect 27712 8449 27721 8483
rect 27721 8449 27755 8483
rect 27755 8449 27764 8483
rect 27712 8440 27764 8449
rect 27804 8483 27856 8492
rect 27804 8449 27814 8483
rect 27814 8449 27848 8483
rect 27848 8449 27856 8483
rect 27804 8440 27856 8449
rect 15292 8304 15344 8356
rect 12624 8236 12676 8288
rect 25320 8304 25372 8356
rect 23020 8236 23072 8288
rect 24584 8236 24636 8288
rect 25228 8279 25280 8288
rect 25228 8245 25237 8279
rect 25237 8245 25271 8279
rect 25271 8245 25280 8279
rect 25228 8236 25280 8245
rect 27252 8236 27304 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 11520 8032 11572 8084
rect 12256 8075 12308 8084
rect 12256 8041 12265 8075
rect 12265 8041 12299 8075
rect 12299 8041 12308 8075
rect 12256 8032 12308 8041
rect 12532 8032 12584 8084
rect 19984 8032 20036 8084
rect 7288 7896 7340 7948
rect 9220 7939 9272 7948
rect 9220 7905 9229 7939
rect 9229 7905 9263 7939
rect 9263 7905 9272 7939
rect 9220 7896 9272 7905
rect 11060 7964 11112 8016
rect 7564 7828 7616 7880
rect 11152 7896 11204 7948
rect 8852 7760 8904 7812
rect 9772 7692 9824 7744
rect 10508 7828 10560 7880
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 10692 7803 10744 7812
rect 10692 7769 10701 7803
rect 10701 7769 10735 7803
rect 10735 7769 10744 7803
rect 10692 7760 10744 7769
rect 12072 7803 12124 7812
rect 12072 7769 12081 7803
rect 12081 7769 12115 7803
rect 12115 7769 12124 7803
rect 12072 7760 12124 7769
rect 12348 7828 12400 7880
rect 13084 7896 13136 7948
rect 20168 7964 20220 8016
rect 14372 7896 14424 7948
rect 15108 7896 15160 7948
rect 18880 7939 18932 7948
rect 18880 7905 18889 7939
rect 18889 7905 18923 7939
rect 18923 7905 18932 7939
rect 18880 7896 18932 7905
rect 18972 7896 19024 7948
rect 14740 7828 14792 7880
rect 15200 7871 15252 7880
rect 15200 7837 15209 7871
rect 15209 7837 15243 7871
rect 15243 7837 15252 7871
rect 15200 7828 15252 7837
rect 17592 7828 17644 7880
rect 17960 7828 18012 7880
rect 18696 7828 18748 7880
rect 19892 7828 19944 7880
rect 20444 7896 20496 7948
rect 20168 7871 20220 7880
rect 20168 7837 20177 7871
rect 20177 7837 20211 7871
rect 20211 7837 20220 7871
rect 20168 7828 20220 7837
rect 20352 7828 20404 7880
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 20904 7871 20956 7880
rect 20904 7837 20913 7871
rect 20913 7837 20947 7871
rect 20947 7837 20956 7871
rect 20904 7828 20956 7837
rect 21456 7896 21508 7948
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 23296 8075 23348 8084
rect 23296 8041 23305 8075
rect 23305 8041 23339 8075
rect 23339 8041 23348 8075
rect 23296 8032 23348 8041
rect 25136 8032 25188 8084
rect 25688 8032 25740 8084
rect 23664 7896 23716 7948
rect 24860 8007 24912 8016
rect 24860 7973 24869 8007
rect 24869 7973 24903 8007
rect 24903 7973 24912 8007
rect 24860 7964 24912 7973
rect 25964 8032 26016 8084
rect 25964 7896 26016 7948
rect 23940 7871 23992 7880
rect 23940 7837 23949 7871
rect 23949 7837 23983 7871
rect 23983 7837 23992 7871
rect 23940 7828 23992 7837
rect 24584 7828 24636 7880
rect 24952 7871 25004 7880
rect 24952 7837 24961 7871
rect 24961 7837 24995 7871
rect 24995 7837 25004 7871
rect 24952 7828 25004 7837
rect 11336 7692 11388 7744
rect 14740 7692 14792 7744
rect 15384 7735 15436 7744
rect 15384 7701 15393 7735
rect 15393 7701 15427 7735
rect 15427 7701 15436 7735
rect 15384 7692 15436 7701
rect 18328 7692 18380 7744
rect 20260 7692 20312 7744
rect 20536 7692 20588 7744
rect 21088 7735 21140 7744
rect 21088 7701 21097 7735
rect 21097 7701 21131 7735
rect 21131 7701 21140 7735
rect 21088 7692 21140 7701
rect 21272 7735 21324 7744
rect 21272 7701 21281 7735
rect 21281 7701 21315 7735
rect 21315 7701 21324 7735
rect 21272 7692 21324 7701
rect 21824 7735 21876 7744
rect 21824 7701 21833 7735
rect 21833 7701 21867 7735
rect 21867 7701 21876 7735
rect 21824 7692 21876 7701
rect 23848 7692 23900 7744
rect 25780 7828 25832 7880
rect 26516 8075 26568 8084
rect 26516 8041 26525 8075
rect 26525 8041 26559 8075
rect 26559 8041 26568 8075
rect 26516 8032 26568 8041
rect 25320 7803 25372 7812
rect 25320 7769 25329 7803
rect 25329 7769 25363 7803
rect 25363 7769 25372 7803
rect 25320 7760 25372 7769
rect 25688 7803 25740 7812
rect 25688 7769 25697 7803
rect 25697 7769 25731 7803
rect 25731 7769 25740 7803
rect 25688 7760 25740 7769
rect 25872 7735 25924 7744
rect 25872 7701 25897 7735
rect 25897 7701 25924 7735
rect 25872 7692 25924 7701
rect 26516 7692 26568 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 16028 7488 16080 7540
rect 16396 7488 16448 7540
rect 18972 7488 19024 7540
rect 20260 7531 20312 7540
rect 20260 7497 20269 7531
rect 20269 7497 20303 7531
rect 20303 7497 20312 7531
rect 20260 7488 20312 7497
rect 8484 7352 8536 7404
rect 8852 7395 8904 7404
rect 8852 7361 8861 7395
rect 8861 7361 8895 7395
rect 8895 7361 8904 7395
rect 8852 7352 8904 7361
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 10600 7420 10652 7472
rect 12072 7420 12124 7472
rect 10508 7352 10560 7404
rect 10968 7352 11020 7404
rect 12808 7352 12860 7404
rect 12992 7352 13044 7404
rect 13452 7352 13504 7404
rect 10416 7327 10468 7336
rect 10416 7293 10425 7327
rect 10425 7293 10459 7327
rect 10459 7293 10468 7327
rect 10416 7284 10468 7293
rect 10600 7284 10652 7336
rect 12440 7284 12492 7336
rect 9312 7259 9364 7268
rect 9312 7225 9321 7259
rect 9321 7225 9355 7259
rect 9355 7225 9364 7259
rect 9312 7216 9364 7225
rect 11152 7216 11204 7268
rect 12348 7216 12400 7268
rect 12716 7191 12768 7200
rect 12716 7157 12725 7191
rect 12725 7157 12759 7191
rect 12759 7157 12768 7191
rect 12716 7148 12768 7157
rect 14372 7420 14424 7472
rect 14740 7352 14792 7404
rect 15108 7395 15160 7404
rect 15108 7361 15117 7395
rect 15117 7361 15151 7395
rect 15151 7361 15160 7395
rect 15108 7352 15160 7361
rect 14924 7327 14976 7336
rect 14924 7293 14933 7327
rect 14933 7293 14967 7327
rect 14967 7293 14976 7327
rect 14924 7284 14976 7293
rect 15384 7420 15436 7472
rect 17592 7420 17644 7472
rect 18328 7420 18380 7472
rect 16120 7352 16172 7404
rect 17500 7352 17552 7404
rect 18420 7395 18472 7404
rect 18420 7361 18429 7395
rect 18429 7361 18463 7395
rect 18463 7361 18472 7395
rect 18420 7352 18472 7361
rect 20536 7488 20588 7540
rect 20812 7488 20864 7540
rect 20628 7463 20680 7472
rect 20628 7429 20637 7463
rect 20637 7429 20671 7463
rect 20671 7429 20680 7463
rect 20628 7420 20680 7429
rect 20904 7420 20956 7472
rect 14832 7148 14884 7200
rect 15292 7191 15344 7200
rect 15292 7157 15301 7191
rect 15301 7157 15335 7191
rect 15335 7157 15344 7191
rect 15292 7148 15344 7157
rect 16304 7216 16356 7268
rect 17960 7284 18012 7336
rect 19984 7284 20036 7336
rect 20536 7216 20588 7268
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 21364 7488 21416 7540
rect 21824 7488 21876 7540
rect 23020 7531 23072 7540
rect 23020 7497 23029 7531
rect 23029 7497 23063 7531
rect 23063 7497 23072 7531
rect 23020 7488 23072 7497
rect 23940 7488 23992 7540
rect 23848 7395 23900 7404
rect 23848 7361 23857 7395
rect 23857 7361 23891 7395
rect 23891 7361 23900 7395
rect 23848 7352 23900 7361
rect 21364 7284 21416 7336
rect 22192 7216 22244 7268
rect 23664 7216 23716 7268
rect 25228 7352 25280 7404
rect 25964 7488 26016 7540
rect 26516 7327 26568 7336
rect 26516 7293 26525 7327
rect 26525 7293 26559 7327
rect 26559 7293 26568 7327
rect 26516 7284 26568 7293
rect 27068 7327 27120 7336
rect 27068 7293 27077 7327
rect 27077 7293 27111 7327
rect 27111 7293 27120 7327
rect 27068 7284 27120 7293
rect 27988 7395 28040 7404
rect 27988 7361 27997 7395
rect 27997 7361 28031 7395
rect 28031 7361 28040 7395
rect 27988 7352 28040 7361
rect 28172 7284 28224 7336
rect 22376 7191 22428 7200
rect 22376 7157 22385 7191
rect 22385 7157 22419 7191
rect 22419 7157 22428 7191
rect 22376 7148 22428 7157
rect 28264 7191 28316 7200
rect 28264 7157 28273 7191
rect 28273 7157 28307 7191
rect 28307 7157 28316 7191
rect 28264 7148 28316 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 8300 6987 8352 6996
rect 8300 6953 8309 6987
rect 8309 6953 8343 6987
rect 8343 6953 8352 6987
rect 8300 6944 8352 6953
rect 8944 6944 8996 6996
rect 10232 6944 10284 6996
rect 7288 6808 7340 6860
rect 9128 6808 9180 6860
rect 12440 6876 12492 6928
rect 12716 6876 12768 6928
rect 13084 6876 13136 6928
rect 7196 6740 7248 6792
rect 7564 6740 7616 6792
rect 8208 6740 8260 6792
rect 8576 6740 8628 6792
rect 8668 6740 8720 6792
rect 9588 6808 9640 6860
rect 10600 6740 10652 6792
rect 10692 6783 10744 6792
rect 10692 6749 10701 6783
rect 10701 6749 10735 6783
rect 10735 6749 10744 6783
rect 10692 6740 10744 6749
rect 12624 6783 12676 6792
rect 12624 6749 12633 6783
rect 12633 6749 12667 6783
rect 12667 6749 12676 6783
rect 12624 6740 12676 6749
rect 13084 6740 13136 6792
rect 15936 6944 15988 6996
rect 17776 6987 17828 6996
rect 17776 6953 17785 6987
rect 17785 6953 17819 6987
rect 17819 6953 17828 6987
rect 17776 6944 17828 6953
rect 21180 6987 21232 6996
rect 21180 6953 21189 6987
rect 21189 6953 21223 6987
rect 21223 6953 21232 6987
rect 21180 6944 21232 6953
rect 23664 6944 23716 6996
rect 23940 6876 23992 6928
rect 16028 6808 16080 6860
rect 9036 6672 9088 6724
rect 10324 6672 10376 6724
rect 11612 6672 11664 6724
rect 14188 6783 14240 6792
rect 14188 6749 14197 6783
rect 14197 6749 14231 6783
rect 14231 6749 14240 6783
rect 14188 6740 14240 6749
rect 18420 6808 18472 6860
rect 19340 6808 19392 6860
rect 16304 6740 16356 6792
rect 17592 6740 17644 6792
rect 10508 6604 10560 6656
rect 10692 6604 10744 6656
rect 12164 6604 12216 6656
rect 13912 6604 13964 6656
rect 16488 6672 16540 6724
rect 17684 6715 17736 6724
rect 17684 6681 17693 6715
rect 17693 6681 17727 6715
rect 17727 6681 17736 6715
rect 17684 6672 17736 6681
rect 18328 6740 18380 6792
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 21088 6808 21140 6860
rect 28172 6851 28224 6860
rect 28172 6817 28181 6851
rect 28181 6817 28215 6851
rect 28215 6817 28224 6851
rect 28172 6808 28224 6817
rect 28448 6851 28500 6860
rect 28448 6817 28457 6851
rect 28457 6817 28491 6851
rect 28491 6817 28500 6851
rect 28448 6808 28500 6817
rect 20168 6783 20220 6792
rect 20168 6749 20177 6783
rect 20177 6749 20211 6783
rect 20211 6749 20220 6783
rect 20168 6740 20220 6749
rect 20352 6783 20404 6792
rect 20352 6749 20361 6783
rect 20361 6749 20395 6783
rect 20395 6749 20404 6783
rect 20352 6740 20404 6749
rect 20812 6740 20864 6792
rect 21364 6783 21416 6792
rect 21364 6749 21373 6783
rect 21373 6749 21407 6783
rect 21407 6749 21416 6783
rect 21364 6740 21416 6749
rect 27988 6740 28040 6792
rect 14464 6604 14516 6656
rect 16120 6604 16172 6656
rect 16580 6647 16632 6656
rect 16580 6613 16589 6647
rect 16589 6613 16623 6647
rect 16623 6613 16632 6647
rect 16580 6604 16632 6613
rect 17776 6604 17828 6656
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 9772 6400 9824 6452
rect 9956 6332 10008 6384
rect 10692 6332 10744 6384
rect 11336 6375 11388 6384
rect 11336 6341 11345 6375
rect 11345 6341 11379 6375
rect 11379 6341 11388 6375
rect 11336 6332 11388 6341
rect 12808 6332 12860 6384
rect 13912 6400 13964 6452
rect 14832 6443 14884 6452
rect 14832 6409 14841 6443
rect 14841 6409 14875 6443
rect 14875 6409 14884 6443
rect 14832 6400 14884 6409
rect 15108 6400 15160 6452
rect 15292 6400 15344 6452
rect 15568 6400 15620 6452
rect 16028 6400 16080 6452
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8484 6264 8536 6316
rect 9680 6307 9732 6316
rect 9680 6273 9689 6307
rect 9689 6273 9723 6307
rect 9723 6273 9732 6307
rect 9680 6264 9732 6273
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 12072 6307 12124 6316
rect 12072 6273 12081 6307
rect 12081 6273 12115 6307
rect 12115 6273 12124 6307
rect 12072 6264 12124 6273
rect 11612 6239 11664 6248
rect 11612 6205 11621 6239
rect 11621 6205 11655 6239
rect 11655 6205 11664 6239
rect 11612 6196 11664 6205
rect 11704 6196 11756 6248
rect 12256 6196 12308 6248
rect 12532 6171 12584 6180
rect 12532 6137 12541 6171
rect 12541 6137 12575 6171
rect 12575 6137 12584 6171
rect 12532 6128 12584 6137
rect 11060 6060 11112 6112
rect 13728 6307 13780 6316
rect 13728 6273 13737 6307
rect 13737 6273 13771 6307
rect 13771 6273 13780 6307
rect 13728 6264 13780 6273
rect 14004 6375 14056 6384
rect 14004 6341 14013 6375
rect 14013 6341 14047 6375
rect 14047 6341 14056 6375
rect 14004 6332 14056 6341
rect 14740 6375 14792 6384
rect 14740 6341 14749 6375
rect 14749 6341 14783 6375
rect 14783 6341 14792 6375
rect 14740 6332 14792 6341
rect 16212 6332 16264 6384
rect 12992 6239 13044 6248
rect 12992 6205 13001 6239
rect 13001 6205 13035 6239
rect 13035 6205 13044 6239
rect 12992 6196 13044 6205
rect 16488 6264 16540 6316
rect 18328 6400 18380 6452
rect 19340 6400 19392 6452
rect 20352 6400 20404 6452
rect 17408 6332 17460 6384
rect 17776 6264 17828 6316
rect 14556 6171 14608 6180
rect 14556 6137 14565 6171
rect 14565 6137 14599 6171
rect 14599 6137 14608 6171
rect 14556 6128 14608 6137
rect 14832 6128 14884 6180
rect 15936 6128 15988 6180
rect 17684 6196 17736 6248
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 16580 6128 16632 6180
rect 16212 6060 16264 6112
rect 16396 6060 16448 6112
rect 17960 6128 18012 6180
rect 18144 6103 18196 6112
rect 18144 6069 18153 6103
rect 18153 6069 18187 6103
rect 18187 6069 18196 6103
rect 18144 6060 18196 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 8484 5856 8536 5908
rect 8760 5856 8812 5908
rect 9680 5856 9732 5908
rect 10416 5856 10468 5908
rect 10600 5856 10652 5908
rect 11060 5856 11112 5908
rect 11612 5856 11664 5908
rect 14188 5856 14240 5908
rect 14924 5856 14976 5908
rect 15384 5856 15436 5908
rect 17408 5899 17460 5908
rect 17408 5865 17417 5899
rect 17417 5865 17451 5899
rect 17451 5865 17460 5899
rect 17408 5856 17460 5865
rect 17960 5856 18012 5908
rect 18144 5856 18196 5908
rect 12808 5831 12860 5840
rect 5172 5695 5224 5704
rect 5172 5661 5181 5695
rect 5181 5661 5215 5695
rect 5215 5661 5224 5695
rect 5172 5652 5224 5661
rect 6552 5652 6604 5704
rect 8208 5652 8260 5704
rect 9772 5720 9824 5772
rect 12808 5797 12817 5831
rect 12817 5797 12851 5831
rect 12851 5797 12860 5831
rect 12808 5788 12860 5797
rect 10232 5652 10284 5704
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 10508 5695 10560 5704
rect 10508 5661 10517 5695
rect 10517 5661 10551 5695
rect 10551 5661 10560 5695
rect 10508 5652 10560 5661
rect 4804 5584 4856 5636
rect 8944 5627 8996 5636
rect 8944 5593 8953 5627
rect 8953 5593 8987 5627
rect 8987 5593 8996 5627
rect 8944 5584 8996 5593
rect 9404 5584 9456 5636
rect 10692 5652 10744 5704
rect 10968 5652 11020 5704
rect 12624 5720 12676 5772
rect 10784 5516 10836 5568
rect 12900 5695 12952 5704
rect 12900 5661 12909 5695
rect 12909 5661 12943 5695
rect 12943 5661 12952 5695
rect 12900 5652 12952 5661
rect 13452 5652 13504 5704
rect 14740 5695 14792 5704
rect 14740 5661 14749 5695
rect 14749 5661 14783 5695
rect 14783 5661 14792 5695
rect 14740 5652 14792 5661
rect 14832 5652 14884 5704
rect 15200 5695 15252 5704
rect 15200 5661 15209 5695
rect 15209 5661 15243 5695
rect 15243 5661 15252 5695
rect 15200 5652 15252 5661
rect 15568 5652 15620 5704
rect 18328 5695 18380 5704
rect 18328 5661 18337 5695
rect 18337 5661 18371 5695
rect 18371 5661 18380 5695
rect 18328 5652 18380 5661
rect 20444 5720 20496 5772
rect 21272 5856 21324 5908
rect 23480 5856 23532 5908
rect 23756 5899 23808 5908
rect 23756 5865 23765 5899
rect 23765 5865 23799 5899
rect 23799 5865 23808 5899
rect 23756 5856 23808 5865
rect 27436 5856 27488 5908
rect 27160 5831 27212 5840
rect 27160 5797 27169 5831
rect 27169 5797 27203 5831
rect 27203 5797 27212 5831
rect 27160 5788 27212 5797
rect 21364 5720 21416 5772
rect 22468 5763 22520 5772
rect 22468 5729 22477 5763
rect 22477 5729 22511 5763
rect 22511 5729 22520 5763
rect 22468 5720 22520 5729
rect 23020 5763 23072 5772
rect 23020 5729 23029 5763
rect 23029 5729 23063 5763
rect 23063 5729 23072 5763
rect 23020 5720 23072 5729
rect 19984 5652 20036 5704
rect 23572 5763 23624 5772
rect 23572 5729 23581 5763
rect 23581 5729 23615 5763
rect 23615 5729 23624 5763
rect 23572 5720 23624 5729
rect 20076 5584 20128 5636
rect 22928 5584 22980 5636
rect 24584 5652 24636 5704
rect 26424 5652 26476 5704
rect 12808 5516 12860 5568
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 19984 5559 20036 5568
rect 19984 5525 19993 5559
rect 19993 5525 20027 5559
rect 20027 5525 20036 5559
rect 19984 5516 20036 5525
rect 24124 5516 24176 5568
rect 25136 5559 25188 5568
rect 25136 5525 25145 5559
rect 25145 5525 25179 5559
rect 25179 5525 25188 5559
rect 25136 5516 25188 5525
rect 27528 5652 27580 5704
rect 28080 5652 28132 5704
rect 28264 5695 28316 5704
rect 28264 5661 28273 5695
rect 28273 5661 28307 5695
rect 28307 5661 28316 5695
rect 28264 5652 28316 5661
rect 28908 5652 28960 5704
rect 27252 5516 27304 5568
rect 27712 5516 27764 5568
rect 28172 5516 28224 5568
rect 28540 5516 28592 5568
rect 29552 5516 29604 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 12072 5312 12124 5364
rect 15200 5312 15252 5364
rect 15476 5312 15528 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 26056 5312 26108 5364
rect 26884 5312 26936 5364
rect 27436 5312 27488 5364
rect 8760 5244 8812 5296
rect 8300 5176 8352 5228
rect 11152 5176 11204 5228
rect 11704 5176 11756 5228
rect 12808 5287 12860 5296
rect 12808 5253 12817 5287
rect 12817 5253 12851 5287
rect 12851 5253 12860 5287
rect 12808 5244 12860 5253
rect 12348 5219 12400 5228
rect 6368 5108 6420 5160
rect 6736 5151 6788 5160
rect 6736 5117 6745 5151
rect 6745 5117 6779 5151
rect 6779 5117 6788 5151
rect 6736 5108 6788 5117
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 13544 5176 13596 5228
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 10968 5040 11020 5092
rect 16580 5244 16632 5296
rect 15936 5176 15988 5228
rect 16212 5176 16264 5228
rect 16304 5219 16356 5228
rect 16304 5185 16313 5219
rect 16313 5185 16347 5219
rect 16347 5185 16356 5219
rect 16304 5176 16356 5185
rect 19984 5219 20036 5228
rect 19984 5185 19993 5219
rect 19993 5185 20027 5219
rect 20027 5185 20036 5219
rect 19984 5176 20036 5185
rect 20076 5176 20128 5228
rect 22376 5176 22428 5228
rect 23020 5176 23072 5228
rect 23572 5219 23624 5228
rect 23572 5185 23581 5219
rect 23581 5185 23615 5219
rect 23615 5185 23624 5219
rect 23572 5176 23624 5185
rect 24124 5176 24176 5228
rect 25136 5176 25188 5228
rect 23756 5108 23808 5160
rect 24400 5151 24452 5160
rect 24400 5117 24409 5151
rect 24409 5117 24443 5151
rect 24443 5117 24452 5151
rect 24400 5108 24452 5117
rect 26424 5219 26476 5228
rect 26424 5185 26433 5219
rect 26433 5185 26467 5219
rect 26467 5185 26476 5219
rect 26424 5176 26476 5185
rect 27160 5176 27212 5228
rect 14740 4972 14792 5024
rect 16028 5015 16080 5024
rect 16028 4981 16037 5015
rect 16037 4981 16071 5015
rect 16071 4981 16080 5015
rect 16028 4972 16080 4981
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 19984 5015 20036 5024
rect 19984 4981 19993 5015
rect 19993 4981 20027 5015
rect 20027 4981 20036 5015
rect 19984 4972 20036 4981
rect 20812 4972 20864 5024
rect 24952 5040 25004 5092
rect 26240 5040 26292 5092
rect 21364 5015 21416 5024
rect 21364 4981 21373 5015
rect 21373 4981 21407 5015
rect 21407 4981 21416 5015
rect 21364 4972 21416 4981
rect 22008 4972 22060 5024
rect 24308 4972 24360 5024
rect 27252 5108 27304 5160
rect 27804 5176 27856 5228
rect 28172 5287 28224 5296
rect 28172 5253 28181 5287
rect 28181 5253 28215 5287
rect 28215 5253 28224 5287
rect 28172 5244 28224 5253
rect 27528 5108 27580 5160
rect 28448 5219 28500 5228
rect 28448 5185 28457 5219
rect 28457 5185 28491 5219
rect 28491 5185 28500 5219
rect 28448 5176 28500 5185
rect 28540 5108 28592 5160
rect 28908 5176 28960 5228
rect 29552 5244 29604 5296
rect 30840 5244 30892 5296
rect 30104 5151 30156 5160
rect 30104 5117 30113 5151
rect 30113 5117 30147 5151
rect 30147 5117 30156 5151
rect 30104 5108 30156 5117
rect 29092 5040 29144 5092
rect 29000 5015 29052 5024
rect 29000 4981 29009 5015
rect 29009 4981 29043 5015
rect 29043 4981 29052 5015
rect 29000 4972 29052 4981
rect 31852 5015 31904 5024
rect 31852 4981 31861 5015
rect 31861 4981 31895 5015
rect 31895 4981 31904 5015
rect 31852 4972 31904 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 11152 4811 11204 4820
rect 11152 4777 11161 4811
rect 11161 4777 11195 4811
rect 11195 4777 11204 4811
rect 11152 4768 11204 4777
rect 16304 4768 16356 4820
rect 16580 4768 16632 4820
rect 17132 4768 17184 4820
rect 18236 4768 18288 4820
rect 19984 4768 20036 4820
rect 27160 4811 27212 4820
rect 27160 4777 27169 4811
rect 27169 4777 27203 4811
rect 27203 4777 27212 4811
rect 27160 4768 27212 4777
rect 7196 4675 7248 4684
rect 7196 4641 7205 4675
rect 7205 4641 7239 4675
rect 7239 4641 7248 4675
rect 7196 4632 7248 4641
rect 9312 4632 9364 4684
rect 10416 4632 10468 4684
rect 12256 4632 12308 4684
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 6552 4564 6604 4616
rect 5448 4539 5500 4548
rect 5448 4505 5457 4539
rect 5457 4505 5491 4539
rect 5491 4505 5500 4539
rect 5448 4496 5500 4505
rect 8300 4496 8352 4548
rect 9220 4539 9272 4548
rect 9220 4505 9229 4539
rect 9229 4505 9263 4539
rect 9263 4505 9272 4539
rect 9220 4496 9272 4505
rect 6368 4428 6420 4480
rect 13728 4564 13780 4616
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 19432 4700 19484 4752
rect 14464 4496 14516 4548
rect 15936 4496 15988 4548
rect 22100 4700 22152 4752
rect 21364 4632 21416 4684
rect 22008 4632 22060 4684
rect 20812 4607 20864 4616
rect 20812 4573 20821 4607
rect 20821 4573 20855 4607
rect 20855 4573 20864 4607
rect 20812 4564 20864 4573
rect 22376 4632 22428 4684
rect 27252 4675 27304 4684
rect 27252 4641 27261 4675
rect 27261 4641 27295 4675
rect 27295 4641 27304 4675
rect 27252 4632 27304 4641
rect 25596 4607 25648 4616
rect 25596 4573 25605 4607
rect 25605 4573 25639 4607
rect 25639 4573 25648 4607
rect 25596 4564 25648 4573
rect 27436 4564 27488 4616
rect 27712 4564 27764 4616
rect 13268 4428 13320 4480
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 18144 4471 18196 4480
rect 18144 4437 18153 4471
rect 18153 4437 18187 4471
rect 18187 4437 18196 4471
rect 18144 4428 18196 4437
rect 22468 4471 22520 4480
rect 22468 4437 22477 4471
rect 22477 4437 22511 4471
rect 22511 4437 22520 4471
rect 22468 4428 22520 4437
rect 24860 4539 24912 4548
rect 24860 4505 24869 4539
rect 24869 4505 24903 4539
rect 24903 4505 24912 4539
rect 24860 4496 24912 4505
rect 27804 4428 27856 4480
rect 27988 4471 28040 4480
rect 27988 4437 27997 4471
rect 27997 4437 28031 4471
rect 28031 4437 28040 4471
rect 27988 4428 28040 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 15936 4224 15988 4276
rect 8208 4156 8260 4208
rect 12072 4156 12124 4208
rect 13268 4156 13320 4208
rect 8300 4088 8352 4140
rect 10508 4088 10560 4140
rect 6368 4063 6420 4072
rect 6368 4029 6377 4063
rect 6377 4029 6411 4063
rect 6411 4029 6420 4063
rect 6368 4020 6420 4029
rect 6644 4063 6696 4072
rect 6644 4029 6653 4063
rect 6653 4029 6687 4063
rect 6687 4029 6696 4063
rect 6644 4020 6696 4029
rect 8760 4063 8812 4072
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 10232 4063 10284 4072
rect 10232 4029 10241 4063
rect 10241 4029 10275 4063
rect 10275 4029 10284 4063
rect 10232 4020 10284 4029
rect 14096 4020 14148 4072
rect 15476 4088 15528 4140
rect 29184 4224 29236 4276
rect 30104 4224 30156 4276
rect 16764 4131 16816 4140
rect 16764 4097 16773 4131
rect 16773 4097 16807 4131
rect 16807 4097 16816 4131
rect 16764 4088 16816 4097
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 23572 4131 23624 4140
rect 23572 4097 23581 4131
rect 23581 4097 23615 4131
rect 23615 4097 23624 4131
rect 23572 4088 23624 4097
rect 23940 4131 23992 4140
rect 23940 4097 23949 4131
rect 23949 4097 23983 4131
rect 23983 4097 23992 4131
rect 23940 4088 23992 4097
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 26700 4088 26752 4140
rect 17224 4063 17276 4072
rect 17224 4029 17233 4063
rect 17233 4029 17267 4063
rect 17267 4029 17276 4063
rect 17224 4020 17276 4029
rect 18420 4020 18472 4072
rect 22192 4020 22244 4072
rect 23296 4020 23348 4072
rect 25228 4020 25280 4072
rect 26424 4020 26476 4072
rect 29092 4063 29144 4072
rect 29092 4029 29101 4063
rect 29101 4029 29135 4063
rect 29135 4029 29144 4063
rect 29092 4020 29144 4029
rect 16028 3952 16080 4004
rect 6828 3884 6880 3936
rect 8484 3884 8536 3936
rect 9312 3884 9364 3936
rect 14372 3927 14424 3936
rect 14372 3893 14381 3927
rect 14381 3893 14415 3927
rect 14415 3893 14424 3927
rect 14372 3884 14424 3893
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 27712 3884 27764 3936
rect 30380 4156 30432 4208
rect 30840 4156 30892 4208
rect 30564 3927 30616 3936
rect 30564 3893 30573 3927
rect 30573 3893 30607 3927
rect 30607 3893 30616 3927
rect 30564 3884 30616 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4160 3544 4212 3596
rect 5080 3680 5132 3732
rect 6000 3476 6052 3528
rect 6552 3476 6604 3528
rect 8668 3680 8720 3732
rect 9036 3544 9088 3596
rect 4896 3451 4948 3460
rect 4896 3417 4905 3451
rect 4905 3417 4939 3451
rect 4939 3417 4948 3451
rect 4896 3408 4948 3417
rect 8300 3476 8352 3528
rect 10508 3544 10560 3596
rect 13268 3680 13320 3732
rect 15660 3680 15712 3732
rect 18236 3680 18288 3732
rect 9312 3476 9364 3528
rect 12900 3544 12952 3596
rect 7012 3451 7064 3460
rect 7012 3417 7021 3451
rect 7021 3417 7055 3451
rect 7055 3417 7064 3451
rect 7012 3408 7064 3417
rect 6828 3340 6880 3392
rect 12348 3476 12400 3528
rect 14096 3476 14148 3528
rect 10048 3451 10100 3460
rect 10048 3417 10057 3451
rect 10057 3417 10091 3451
rect 10091 3417 10100 3451
rect 10048 3408 10100 3417
rect 12900 3408 12952 3460
rect 14004 3408 14056 3460
rect 11060 3340 11112 3392
rect 12256 3340 12308 3392
rect 16580 3408 16632 3460
rect 16488 3340 16540 3392
rect 18696 3544 18748 3596
rect 23664 3680 23716 3732
rect 23940 3723 23992 3732
rect 23940 3689 23949 3723
rect 23949 3689 23983 3723
rect 23983 3689 23992 3723
rect 23940 3680 23992 3689
rect 24308 3680 24360 3732
rect 24400 3680 24452 3732
rect 22468 3587 22520 3596
rect 22468 3553 22477 3587
rect 22477 3553 22511 3587
rect 22511 3553 22520 3587
rect 22468 3544 22520 3553
rect 17868 3408 17920 3460
rect 19892 3519 19944 3528
rect 19892 3485 19901 3519
rect 19901 3485 19935 3519
rect 19935 3485 19944 3519
rect 19892 3476 19944 3485
rect 21824 3476 21876 3528
rect 21916 3519 21968 3528
rect 21916 3485 21925 3519
rect 21925 3485 21959 3519
rect 21959 3485 21968 3519
rect 21916 3476 21968 3485
rect 26516 3680 26568 3732
rect 28816 3680 28868 3732
rect 29184 3680 29236 3732
rect 26240 3612 26292 3664
rect 28724 3612 28776 3664
rect 24400 3519 24452 3528
rect 24400 3485 24409 3519
rect 24409 3485 24443 3519
rect 24443 3485 24452 3519
rect 24400 3476 24452 3485
rect 29092 3544 29144 3596
rect 29276 3612 29328 3664
rect 32312 3544 32364 3596
rect 26240 3519 26292 3528
rect 26240 3485 26249 3519
rect 26249 3485 26283 3519
rect 26283 3485 26292 3519
rect 26240 3476 26292 3485
rect 21088 3451 21140 3460
rect 21088 3417 21097 3451
rect 21097 3417 21131 3451
rect 21131 3417 21140 3451
rect 21088 3408 21140 3417
rect 22928 3408 22980 3460
rect 25320 3408 25372 3460
rect 26976 3408 27028 3460
rect 28816 3340 28868 3392
rect 29184 3476 29236 3528
rect 31024 3519 31076 3528
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 31852 3476 31904 3528
rect 33600 3340 33652 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 6828 3136 6880 3188
rect 6000 3068 6052 3120
rect 8484 3136 8536 3188
rect 8760 3136 8812 3188
rect 13268 3136 13320 3188
rect 8944 3111 8996 3120
rect 8944 3077 8953 3111
rect 8953 3077 8987 3111
rect 8987 3077 8996 3111
rect 8944 3068 8996 3077
rect 10508 3068 10560 3120
rect 11152 3068 11204 3120
rect 12900 3068 12952 3120
rect 13544 3111 13596 3120
rect 13544 3077 13553 3111
rect 13553 3077 13587 3111
rect 13587 3077 13596 3111
rect 13544 3068 13596 3077
rect 15568 3136 15620 3188
rect 16580 3136 16632 3188
rect 16672 3068 16724 3120
rect 8300 3000 8352 3052
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 12256 3000 12308 3052
rect 13084 3000 13136 3052
rect 17868 3136 17920 3188
rect 18144 3068 18196 3120
rect 21916 3136 21968 3188
rect 22100 3111 22152 3120
rect 22100 3077 22109 3111
rect 22109 3077 22143 3111
rect 22143 3077 22152 3111
rect 22100 3068 22152 3077
rect 22928 3136 22980 3188
rect 23480 3068 23532 3120
rect 25320 3136 25372 3188
rect 25596 3136 25648 3188
rect 27528 3136 27580 3188
rect 26976 3068 27028 3120
rect 27712 3068 27764 3120
rect 4160 2975 4212 2984
rect 4160 2941 4169 2975
rect 4169 2941 4203 2975
rect 4203 2941 4212 2975
rect 4160 2932 4212 2941
rect 4436 2975 4488 2984
rect 4436 2941 4445 2975
rect 4445 2941 4479 2975
rect 4479 2941 4488 2975
rect 4436 2932 4488 2941
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 10324 2932 10376 2984
rect 11060 2975 11112 2984
rect 11060 2941 11069 2975
rect 11069 2941 11103 2975
rect 11103 2941 11112 2975
rect 11060 2932 11112 2941
rect 14096 2932 14148 2984
rect 23572 3000 23624 3052
rect 23664 3043 23716 3052
rect 23664 3009 23673 3043
rect 23673 3009 23707 3043
rect 23707 3009 23716 3043
rect 23664 3000 23716 3009
rect 26240 3000 26292 3052
rect 29184 3136 29236 3188
rect 30564 3136 30616 3188
rect 29000 3068 29052 3120
rect 30380 3068 30432 3120
rect 28816 3043 28868 3052
rect 19800 2975 19852 2984
rect 19800 2941 19809 2975
rect 19809 2941 19843 2975
rect 19843 2941 19852 2975
rect 19800 2932 19852 2941
rect 19432 2864 19484 2916
rect 20168 2932 20220 2984
rect 21824 2975 21876 2984
rect 21824 2941 21833 2975
rect 21833 2941 21867 2975
rect 21867 2941 21876 2975
rect 21824 2932 21876 2941
rect 28816 3009 28825 3043
rect 28825 3009 28859 3043
rect 28859 3009 28868 3043
rect 28816 3000 28868 3009
rect 33600 3179 33652 3188
rect 33600 3145 33609 3179
rect 33609 3145 33643 3179
rect 33643 3145 33652 3179
rect 33600 3136 33652 3145
rect 26884 2932 26936 2984
rect 26976 2975 27028 2984
rect 26976 2941 26985 2975
rect 26985 2941 27019 2975
rect 27019 2941 27028 2975
rect 26976 2932 27028 2941
rect 27804 2932 27856 2984
rect 33324 3000 33376 3052
rect 31300 2932 31352 2984
rect 8576 2796 8628 2848
rect 11796 2839 11848 2848
rect 11796 2805 11805 2839
rect 11805 2805 11839 2839
rect 11839 2805 11848 2839
rect 11796 2796 11848 2805
rect 21824 2796 21876 2848
rect 27436 2796 27488 2848
rect 30380 2796 30432 2848
rect 32128 2796 32180 2848
rect 34244 2796 34296 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4620 2592 4672 2644
rect 4896 2592 4948 2644
rect 5448 2592 5500 2644
rect 6736 2592 6788 2644
rect 7012 2592 7064 2644
rect 7196 2592 7248 2644
rect 9220 2592 9272 2644
rect 10048 2592 10100 2644
rect 11060 2592 11112 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 14004 2592 14056 2644
rect 14464 2635 14516 2644
rect 14464 2601 14473 2635
rect 14473 2601 14507 2635
rect 14507 2601 14516 2635
rect 14464 2592 14516 2601
rect 16764 2592 16816 2644
rect 16856 2592 16908 2644
rect 6644 2524 6696 2576
rect 14096 2524 14148 2576
rect 16580 2524 16632 2576
rect 16672 2567 16724 2576
rect 16672 2533 16681 2567
rect 16681 2533 16715 2567
rect 16715 2533 16724 2567
rect 16672 2524 16724 2533
rect 940 2388 992 2440
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 11796 2499 11848 2508
rect 11796 2465 11805 2499
rect 11805 2465 11839 2499
rect 11839 2465 11848 2499
rect 11796 2456 11848 2465
rect 13544 2499 13596 2508
rect 13544 2465 13553 2499
rect 13553 2465 13587 2499
rect 13587 2465 13596 2499
rect 13544 2456 13596 2465
rect 15476 2456 15528 2508
rect 15568 2456 15620 2508
rect 4804 2388 4856 2440
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 6000 2388 6052 2440
rect 7012 2388 7064 2440
rect 8300 2431 8352 2440
rect 8300 2397 8309 2431
rect 8309 2397 8343 2431
rect 8343 2397 8352 2431
rect 8300 2388 8352 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 10048 2388 10100 2440
rect 11060 2388 11112 2440
rect 13268 2388 13320 2440
rect 14096 2388 14148 2440
rect 16672 2388 16724 2440
rect 14924 2320 14976 2372
rect 18696 2388 18748 2440
rect 19340 2456 19392 2508
rect 20260 2456 20312 2508
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 17868 2320 17920 2372
rect 14372 2252 14424 2304
rect 26700 2592 26752 2644
rect 31024 2592 31076 2644
rect 23664 2456 23716 2508
rect 24952 2499 25004 2508
rect 24952 2465 24961 2499
rect 24961 2465 24995 2499
rect 24995 2465 25004 2499
rect 24952 2456 25004 2465
rect 26976 2456 27028 2508
rect 27528 2499 27580 2508
rect 27528 2465 27537 2499
rect 27537 2465 27571 2499
rect 27571 2465 27580 2499
rect 27528 2456 27580 2465
rect 27896 2456 27948 2508
rect 30472 2456 30524 2508
rect 34244 2499 34296 2508
rect 34244 2465 34253 2499
rect 34253 2465 34287 2499
rect 34287 2465 34296 2499
rect 34244 2456 34296 2465
rect 29092 2388 29144 2440
rect 32128 2431 32180 2440
rect 32128 2397 32137 2431
rect 32137 2397 32171 2431
rect 32171 2397 32180 2431
rect 32128 2388 32180 2397
rect 34520 2431 34572 2440
rect 34520 2397 34529 2431
rect 34529 2397 34563 2431
rect 34563 2397 34572 2431
rect 34520 2388 34572 2397
rect 35348 2388 35400 2440
rect 27712 2320 27764 2372
rect 30380 2320 30432 2372
rect 25320 2252 25372 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 18052 19372 18104 19378
rect 18052 19314 18104 19320
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 18064 18834 18092 19314
rect 18236 19168 18288 19174
rect 18236 19110 18288 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 16488 18760 16540 18766
rect 16488 18702 16540 18708
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 11348 17678 11376 18226
rect 12636 18222 12664 18702
rect 12728 18426 12756 18702
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 11532 17678 11560 18158
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11520 17672 11572 17678
rect 11520 17614 11572 17620
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 9956 17196 10008 17202
rect 9876 17156 9956 17184
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 9232 15026 9260 16594
rect 9692 15706 9720 17070
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9784 16046 9812 16458
rect 9876 16454 9904 17156
rect 9956 17138 10008 17144
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 9784 15586 9812 15982
rect 9692 15558 9812 15586
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 9232 14550 9260 14962
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 8864 12850 8892 13738
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12850 8984 13126
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 9140 11354 9168 14350
rect 9232 14346 9260 14486
rect 9508 14414 9536 15098
rect 9692 15026 9720 15558
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9784 15094 9812 15370
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9588 15020 9640 15026
rect 9588 14962 9640 14968
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9600 14482 9628 14962
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9496 14408 9548 14414
rect 9496 14350 9548 14356
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 9232 13954 9260 14282
rect 9508 14074 9536 14350
rect 9692 14278 9720 14962
rect 9784 14618 9812 15030
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 14074 9720 14214
rect 9496 14068 9548 14074
rect 9496 14010 9548 14016
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9232 13926 9352 13954
rect 9220 12912 9272 12918
rect 9220 12854 9272 12860
rect 9232 11898 9260 12854
rect 9324 12442 9352 13926
rect 9772 13252 9824 13258
rect 9772 13194 9824 13200
rect 9784 12986 9812 13194
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9876 12918 9904 16390
rect 9968 15502 9996 16526
rect 10060 16454 10088 17070
rect 10428 16794 10456 17614
rect 11060 17604 11112 17610
rect 11060 17546 11112 17552
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9956 15496 10008 15502
rect 9956 15438 10008 15444
rect 9968 15162 9996 15438
rect 9956 15156 10008 15162
rect 9956 15098 10008 15104
rect 9956 14884 10008 14890
rect 9956 14826 10008 14832
rect 9968 14482 9996 14826
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 9956 13864 10008 13870
rect 9956 13806 10008 13812
rect 9968 13326 9996 13806
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9968 12594 9996 12718
rect 10060 12646 10088 16390
rect 10704 16114 10732 17478
rect 11072 16182 11100 17546
rect 11348 17338 11376 17614
rect 11532 17542 11560 17614
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 12084 17338 12112 17614
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12176 17270 12204 17546
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 12544 17202 12572 17478
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10244 15162 10272 15642
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10152 14618 10180 14962
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 10336 14550 10364 16050
rect 10704 15638 10732 16050
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11428 15904 11480 15910
rect 11428 15846 11480 15852
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 11348 15570 11376 15846
rect 11440 15706 11468 15846
rect 11428 15700 11480 15706
rect 11428 15642 11480 15648
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 12164 15564 12216 15570
rect 12164 15506 12216 15512
rect 11980 15496 12032 15502
rect 11980 15438 12032 15444
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11336 15428 11388 15434
rect 11336 15370 11388 15376
rect 10428 15162 10456 15370
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10704 15026 10732 15302
rect 11072 15162 11100 15370
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10324 14544 10376 14550
rect 10324 14486 10376 14492
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10520 13870 10548 14418
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 10508 13864 10560 13870
rect 10508 13806 10560 13812
rect 10232 13184 10284 13190
rect 10232 13126 10284 13132
rect 9876 12566 9996 12594
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 9312 12436 9364 12442
rect 9876 12434 9904 12566
rect 9876 12406 9996 12434
rect 9312 12378 9364 12384
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9220 11892 9272 11898
rect 9220 11834 9272 11840
rect 9324 11558 9352 12174
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9416 11694 9444 12038
rect 9600 11898 9628 12242
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9784 11762 9812 12174
rect 9876 12102 9904 12310
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9968 11762 9996 12406
rect 10244 12102 10272 13126
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9956 11756 10008 11762
rect 9956 11698 10008 11704
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 9324 11150 9352 11494
rect 9312 11144 9364 11150
rect 9312 11086 9364 11092
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 7748 10056 7800 10062
rect 7748 9998 7800 10004
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 7760 8566 7788 9998
rect 8760 9580 8812 9586
rect 8760 9522 8812 9528
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 8772 8498 8800 9522
rect 9232 8566 9260 9522
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 7300 7954 7328 8434
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 7300 6866 7328 7890
rect 7576 7886 7604 8434
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7288 6860 7340 6866
rect 7288 6802 7340 6808
rect 7576 6798 7604 7822
rect 8220 6798 8248 8434
rect 8484 7404 8536 7410
rect 8484 7346 8536 7352
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4160 3596 4212 3602
rect 4160 3538 4212 3544
rect 4172 2990 4200 3538
rect 4160 2984 4212 2990
rect 4160 2926 4212 2932
rect 4436 2984 4488 2990
rect 4488 2932 4660 2938
rect 4436 2926 4660 2932
rect 4448 2910 4660 2926
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4632 2650 4660 2910
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4816 2446 4844 5578
rect 5184 4622 5212 5646
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5184 3754 5212 4558
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5092 3738 5212 3754
rect 5080 3732 5212 3738
rect 5132 3726 5212 3732
rect 5080 3674 5132 3680
rect 4896 3460 4948 3466
rect 4896 3402 4948 3408
rect 4908 2650 4936 3402
rect 5460 2650 5488 4490
rect 6380 4486 6408 5102
rect 6564 4622 6592 5646
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 4078 6408 4422
rect 6368 4072 6420 4078
rect 6368 4014 6420 4020
rect 6564 3534 6592 4558
rect 6644 4072 6696 4078
rect 6644 4014 6696 4020
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6012 3126 6040 3470
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 6656 2582 6684 4014
rect 6748 2650 6776 5102
rect 7208 4690 7236 6734
rect 8220 5710 8248 6734
rect 8312 6322 8340 6938
rect 8496 6322 8524 7346
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8300 6316 8352 6322
rect 8300 6258 8352 6264
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8496 5914 8524 6258
rect 8484 5908 8536 5914
rect 8484 5850 8536 5856
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 8220 4214 8248 5646
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8312 4554 8340 5170
rect 8300 4548 8352 4554
rect 8300 4490 8352 4496
rect 8208 4208 8260 4214
rect 8208 4150 8260 4156
rect 8312 4146 8340 4490
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6840 3398 6868 3878
rect 8312 3534 8340 4082
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 7012 3460 7064 3466
rect 7012 3402 7064 3408
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6840 3194 6868 3334
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 7024 2650 7052 3402
rect 8312 3058 8340 3470
rect 8496 3194 8524 3878
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7208 2650 7236 2926
rect 8588 2854 8616 6734
rect 8680 3738 8708 6734
rect 8772 5914 8800 8434
rect 9128 8356 9180 8362
rect 9128 8298 9180 8304
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 8864 7818 8892 8230
rect 8852 7812 8904 7818
rect 8852 7754 8904 7760
rect 8864 7410 8892 7754
rect 8852 7404 8904 7410
rect 8852 7346 8904 7352
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8956 7002 8984 7346
rect 8944 6996 8996 7002
rect 8944 6938 8996 6944
rect 9140 6866 9168 8298
rect 9232 7954 9260 8502
rect 9220 7948 9272 7954
rect 9220 7890 9272 7896
rect 9324 7274 9352 11086
rect 9416 11014 9444 11630
rect 9784 11150 9812 11698
rect 9772 11144 9824 11150
rect 9772 11086 9824 11092
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10470 9444 10950
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9926 9444 9998
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 9036 6724 9088 6730
rect 9036 6666 9088 6672
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8772 5302 8800 5850
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8772 3194 8800 4014
rect 8760 3188 8812 3194
rect 8760 3130 8812 3136
rect 8956 3126 8984 5578
rect 9048 3602 9076 6666
rect 9416 5642 9444 9862
rect 9588 8356 9640 8362
rect 9588 8298 9640 8304
rect 9600 6866 9628 8298
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9784 6458 9812 7686
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9692 5914 9720 6258
rect 9680 5908 9732 5914
rect 9680 5850 9732 5856
rect 9784 5778 9812 6394
rect 9968 6390 9996 11698
rect 10232 11552 10284 11558
rect 10230 11520 10232 11529
rect 10336 11540 10364 13806
rect 10520 13394 10548 13806
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10428 12782 10456 13126
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10428 12238 10456 12718
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10520 11778 10548 13330
rect 10704 12918 10732 14962
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11072 14074 11100 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 13530 10824 13874
rect 11072 13818 11100 14010
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10980 13790 11100 13818
rect 10784 13524 10836 13530
rect 10784 13466 10836 13472
rect 10692 12912 10744 12918
rect 10692 12854 10744 12860
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10796 12442 10824 12786
rect 10784 12436 10836 12442
rect 10784 12378 10836 12384
rect 10284 11520 10364 11540
rect 10286 11512 10364 11520
rect 10428 11750 10548 11778
rect 10784 11756 10836 11762
rect 10230 11455 10286 11464
rect 10428 11370 10456 11750
rect 10784 11698 10836 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10152 11342 10456 11370
rect 10152 8430 10180 11342
rect 10232 11144 10284 11150
rect 10232 11086 10284 11092
rect 10244 8974 10272 11086
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10336 8974 10364 11018
rect 10520 10690 10548 11630
rect 10428 10674 10548 10690
rect 10796 10674 10824 11698
rect 10416 10668 10548 10674
rect 10468 10662 10548 10668
rect 10784 10668 10836 10674
rect 10416 10610 10468 10616
rect 10784 10610 10836 10616
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10244 8634 10272 8910
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10244 7002 10272 8298
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10336 6730 10364 8910
rect 10428 7342 10456 10610
rect 10508 7880 10560 7886
rect 10508 7822 10560 7828
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10520 7410 10548 7822
rect 10612 7478 10640 7822
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10324 6724 10376 6730
rect 10324 6666 10376 6672
rect 10520 6662 10548 7346
rect 10600 7336 10652 7342
rect 10600 7278 10652 7284
rect 10612 6798 10640 7278
rect 10704 6798 10732 7754
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 9956 6384 10008 6390
rect 9956 6326 10008 6332
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 9772 5772 9824 5778
rect 9772 5714 9824 5720
rect 10244 5710 10272 6258
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10428 5710 10456 5850
rect 10520 5710 10548 6598
rect 10612 5914 10640 6734
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6390 10732 6598
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10508 5704 10560 5710
rect 10692 5704 10744 5710
rect 10560 5652 10692 5658
rect 10508 5646 10744 5652
rect 9404 5636 9456 5642
rect 9404 5578 9456 5584
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 9232 2650 9260 4490
rect 9324 3942 9352 4626
rect 10244 4078 10272 5646
rect 10232 4072 10284 4078
rect 10232 4014 10284 4020
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9324 3534 9352 3878
rect 9312 3528 9364 3534
rect 9312 3470 9364 3476
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10060 2650 10088 3402
rect 10336 2990 10364 5646
rect 10428 4690 10456 5646
rect 10520 5630 10732 5646
rect 10796 5574 10824 10610
rect 10888 10266 10916 13738
rect 10980 13258 11008 13790
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 13326 11100 13670
rect 11060 13320 11112 13326
rect 11060 13262 11112 13268
rect 10968 13252 11020 13258
rect 10968 13194 11020 13200
rect 11072 12374 11100 13262
rect 11164 13190 11192 14214
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11348 13002 11376 15370
rect 11992 15162 12020 15438
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11624 14414 11652 14486
rect 11716 14414 11744 14962
rect 12084 14550 12112 14962
rect 12176 14618 12204 15506
rect 12164 14612 12216 14618
rect 12164 14554 12216 14560
rect 12544 14550 12572 17138
rect 12636 14958 12664 18158
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17746 13124 18022
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13004 17338 13032 17614
rect 13096 17338 13124 17682
rect 13176 17536 13228 17542
rect 13176 17478 13228 17484
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 13188 17202 13216 17478
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13372 16114 13400 17478
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13740 16182 13768 16458
rect 14292 16250 14320 18226
rect 14844 17882 14872 18226
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 15212 17678 15240 18022
rect 15304 17678 15332 18226
rect 15764 17814 15792 18226
rect 15936 18080 15988 18086
rect 15936 18022 15988 18028
rect 15948 17882 15976 18022
rect 16500 17882 16528 18702
rect 16592 18358 16620 18770
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 16592 17882 16620 18294
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15212 17270 15240 17614
rect 15304 17338 15332 17614
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15200 17264 15252 17270
rect 15200 17206 15252 17212
rect 14740 16720 14792 16726
rect 14740 16662 14792 16668
rect 14752 16590 14780 16662
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14280 16244 14332 16250
rect 14280 16186 14332 16192
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 12912 15706 12940 15982
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 13372 15638 13400 16050
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15706 13860 15982
rect 14476 15910 14504 16390
rect 14660 16046 14688 16390
rect 14752 16046 14780 16526
rect 14832 16448 14884 16454
rect 14832 16390 14884 16396
rect 14844 16250 14872 16390
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14372 15904 14424 15910
rect 14372 15846 14424 15852
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12072 14544 12124 14550
rect 12072 14486 12124 14492
rect 12532 14544 12584 14550
rect 12532 14486 12584 14492
rect 12636 14482 12664 14894
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12912 14414 12940 15302
rect 13280 15026 13308 15302
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 11612 14408 11664 14414
rect 11612 14350 11664 14356
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 12440 14408 12492 14414
rect 12440 14350 12492 14356
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 14004 14408 14056 14414
rect 14004 14350 14056 14356
rect 11624 14260 11652 14350
rect 11796 14272 11848 14278
rect 11624 14232 11744 14260
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11164 12986 11376 13002
rect 11152 12980 11376 12986
rect 11204 12974 11376 12980
rect 11152 12922 11204 12928
rect 11440 12850 11468 13126
rect 11152 12844 11204 12850
rect 11152 12786 11204 12792
rect 11428 12844 11480 12850
rect 11428 12786 11480 12792
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11072 11762 11100 12174
rect 11164 11898 11192 12786
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11256 12442 11284 12650
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11256 12238 11284 12378
rect 11532 12238 11560 12650
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11428 12232 11480 12238
rect 11428 12174 11480 12180
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 11256 11762 11284 12038
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11072 11354 11100 11698
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10888 9722 10916 10202
rect 11072 10062 11100 11018
rect 11256 10742 11284 11698
rect 11440 11540 11468 12174
rect 11624 11694 11652 12310
rect 11716 12220 11744 14232
rect 11796 14214 11848 14220
rect 11808 14074 11836 14214
rect 12452 14074 12480 14350
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 12440 14068 12492 14074
rect 12440 14010 12492 14016
rect 11808 13802 11836 14010
rect 12912 13870 12940 14350
rect 13280 14074 13308 14350
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13648 13870 13676 14214
rect 13924 14006 13952 14214
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 13636 13864 13688 13870
rect 13636 13806 13688 13812
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11808 12374 11836 12786
rect 11992 12714 12020 13466
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12268 12850 12296 13126
rect 12256 12844 12308 12850
rect 12256 12786 12308 12792
rect 11888 12708 11940 12714
rect 11888 12650 11940 12656
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11900 12442 11928 12650
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11796 12368 11848 12374
rect 11796 12310 11848 12316
rect 11992 12238 12020 12650
rect 12268 12442 12296 12786
rect 12256 12436 12308 12442
rect 12256 12378 12308 12384
rect 11980 12232 12032 12238
rect 11716 12192 11836 12220
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11520 11552 11572 11558
rect 11440 11512 11520 11540
rect 11520 11494 11572 11500
rect 11532 11286 11560 11494
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11624 11218 11652 11630
rect 11704 11552 11756 11558
rect 11704 11494 11756 11500
rect 11716 11354 11744 11494
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10968 9580 11020 9586
rect 10968 9522 11020 9528
rect 10980 9432 11008 9522
rect 10888 9404 11008 9432
rect 10888 8430 10916 9404
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11072 8022 11100 8434
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11152 7948 11204 7954
rect 11152 7890 11204 7896
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 5710 11008 7346
rect 11164 7274 11192 7890
rect 11348 7750 11376 10406
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11532 8090 11560 8434
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11348 6390 11376 7686
rect 11624 6730 11652 11154
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11716 9654 11744 9998
rect 11808 9926 11836 12192
rect 11980 12174 12032 12180
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12176 11354 12204 11698
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 11098 12112 11154
rect 12360 11150 12388 12174
rect 12348 11144 12400 11150
rect 12084 11092 12348 11098
rect 12084 11086 12400 11092
rect 12084 11070 12388 11086
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 11888 10056 11940 10062
rect 11888 9998 11940 10004
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11900 9586 11928 9998
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 8786 11928 9522
rect 11900 8758 12112 8786
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11992 8362 12020 8570
rect 12084 8566 12112 8758
rect 12072 8560 12124 8566
rect 12072 8502 12124 8508
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7478 12112 7754
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11612 6724 11664 6730
rect 11612 6666 11664 6672
rect 11336 6384 11388 6390
rect 11336 6326 11388 6332
rect 12084 6322 12112 7414
rect 12176 6662 12204 10406
rect 12452 10062 12480 13806
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 11694 13400 12174
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12714 11520 12770 11529
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12452 9450 12480 9998
rect 12440 9444 12492 9450
rect 12440 9386 12492 9392
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12072 6316 12124 6322
rect 12072 6258 12124 6264
rect 11612 6248 11664 6254
rect 11612 6190 11664 6196
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5914 11100 6054
rect 11624 5914 11652 6190
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10980 5098 11008 5646
rect 11716 5234 11744 6190
rect 12084 5370 12112 6258
rect 12268 6254 12296 8026
rect 12360 7886 12388 8298
rect 12544 8090 12572 8434
rect 12636 8294 12664 11494
rect 12714 11455 12770 11464
rect 12728 11218 12756 11455
rect 12716 11212 12768 11218
rect 12716 11154 12768 11160
rect 13372 11150 13400 11630
rect 13648 11558 13676 13806
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13832 12238 13860 13194
rect 13924 13190 13952 13942
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13820 11688 13872 11694
rect 13924 11676 13952 13126
rect 13872 11648 13952 11676
rect 13820 11630 13872 11636
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13832 10826 13860 11630
rect 14016 11540 14044 14350
rect 14384 13870 14412 15846
rect 14476 15502 14504 15846
rect 14752 15638 14780 15982
rect 14740 15632 14792 15638
rect 14740 15574 14792 15580
rect 14844 15502 14872 16186
rect 15016 16040 15068 16046
rect 15016 15982 15068 15988
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 14476 14074 14504 15438
rect 14936 15434 14964 15846
rect 15028 15706 15056 15982
rect 15304 15706 15332 17274
rect 15384 17264 15436 17270
rect 15384 17206 15436 17212
rect 15396 16658 15424 17206
rect 15764 16998 15792 17750
rect 15948 17338 15976 17818
rect 16396 17740 16448 17746
rect 16396 17682 16448 17688
rect 16304 17672 16356 17678
rect 16304 17614 16356 17620
rect 16028 17536 16080 17542
rect 16028 17478 16080 17484
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 16040 17202 16068 17478
rect 16316 17338 16344 17614
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16028 17196 16080 17202
rect 16028 17138 16080 17144
rect 15752 16992 15804 16998
rect 16408 16946 16436 17682
rect 16500 17202 16528 17818
rect 17972 17746 18000 18294
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16868 17626 16896 17682
rect 17040 17672 17092 17678
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16592 16998 16620 17614
rect 16868 17598 16988 17626
rect 17040 17614 17092 17620
rect 17132 17672 17184 17678
rect 17132 17614 17184 17620
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 17270 16712 17478
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16672 17264 16724 17270
rect 16672 17206 16724 17212
rect 15752 16934 15804 16940
rect 15764 16794 15792 16934
rect 16316 16918 16436 16946
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 16316 16658 16344 16918
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15488 16114 15516 16390
rect 15476 16108 15528 16114
rect 15476 16050 15528 16056
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 16028 16108 16080 16114
rect 16028 16050 16080 16056
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 14924 15428 14976 15434
rect 14924 15370 14976 15376
rect 14936 14618 14964 15370
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14464 13932 14516 13938
rect 14568 13920 14596 14214
rect 14752 14006 14780 14214
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14516 13892 14596 13920
rect 14648 13932 14700 13938
rect 14464 13874 14516 13880
rect 14648 13874 14700 13880
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 14476 13462 14504 13874
rect 14464 13456 14516 13462
rect 14464 13398 14516 13404
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14384 12170 14412 12786
rect 14476 12306 14504 13398
rect 14660 13326 14688 13874
rect 14752 13326 14780 13942
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14844 13530 14872 13670
rect 14832 13524 14884 13530
rect 14832 13466 14884 13472
rect 14936 13394 14964 13874
rect 15028 13530 15056 15642
rect 15948 15502 15976 16050
rect 16040 15502 16068 16050
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 16028 15496 16080 15502
rect 16028 15438 16080 15444
rect 15016 13524 15068 13530
rect 15016 13466 15068 13472
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14648 13320 14700 13326
rect 14648 13262 14700 13268
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14844 13190 14872 13330
rect 14740 13184 14792 13190
rect 14660 13144 14740 13172
rect 14464 12300 14516 12306
rect 14464 12242 14516 12248
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14200 11898 14228 12106
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14200 11558 14228 11834
rect 13740 10810 13860 10826
rect 13728 10804 13860 10810
rect 13780 10798 13860 10804
rect 13924 11512 14044 11540
rect 14188 11552 14240 11558
rect 13728 10746 13780 10752
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12636 7970 12664 8230
rect 12544 7942 12664 7970
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 10968 5092 11020 5098
rect 10968 5034 11020 5040
rect 11164 4826 11192 5170
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 12084 4214 12112 5306
rect 12360 5234 12388 7210
rect 12452 6934 12480 7278
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12256 4684 12308 4690
rect 12256 4626 12308 4632
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10520 3602 10548 4082
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10520 3126 10548 3538
rect 12268 3398 12296 4626
rect 12452 3618 12480 6870
rect 12544 6186 12572 7942
rect 13004 7410 13032 10610
rect 13924 10538 13952 11512
rect 14188 11494 14240 11500
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13912 10532 13964 10538
rect 13912 10474 13964 10480
rect 13464 9994 13492 10474
rect 13728 10192 13780 10198
rect 13556 10140 13728 10146
rect 13556 10134 13780 10140
rect 13556 10130 13768 10134
rect 13544 10124 13768 10130
rect 13596 10118 13768 10124
rect 13544 10066 13596 10072
rect 13452 9988 13504 9994
rect 13452 9930 13504 9936
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13096 7954 13124 8434
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12728 6934 12756 7142
rect 12716 6928 12768 6934
rect 12716 6870 12768 6876
rect 12624 6792 12676 6798
rect 12624 6734 12676 6740
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12636 5778 12664 6734
rect 12820 6390 12848 7346
rect 13084 6928 13136 6934
rect 13084 6870 13136 6876
rect 13096 6798 13124 6870
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12820 5846 12848 6326
rect 12992 6248 13044 6254
rect 12912 6208 12992 6236
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12912 5710 12940 6208
rect 13096 6236 13124 6734
rect 13044 6208 13124 6236
rect 12992 6190 13044 6196
rect 13464 5710 13492 7346
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 6458 13952 6598
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 14016 6390 14044 10610
rect 14200 10062 14228 11494
rect 14384 11121 14412 12106
rect 14476 11762 14504 12242
rect 14464 11756 14516 11762
rect 14464 11698 14516 11704
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14370 10976 14426 10985
rect 14370 10911 14426 10920
rect 14384 10742 14412 10911
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 8906 14228 9998
rect 14292 9110 14320 10066
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 14200 8498 14228 8842
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14384 7954 14412 9930
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14370 7848 14426 7857
rect 14370 7783 14426 7792
rect 14384 7478 14412 7783
rect 14372 7472 14424 7478
rect 14372 7414 14424 7420
rect 14188 6792 14240 6798
rect 14188 6734 14240 6740
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 12900 5704 12952 5710
rect 12900 5646 12952 5652
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12820 5302 12848 5510
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12360 3590 12480 3618
rect 12912 3602 12940 5646
rect 13268 4480 13320 4486
rect 13268 4422 13320 4428
rect 13280 4214 13308 4422
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13280 3738 13308 4150
rect 13268 3732 13320 3738
rect 13268 3674 13320 3680
rect 12900 3596 12952 3602
rect 12360 3534 12388 3590
rect 12900 3538 12952 3544
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 11060 3392 11112 3398
rect 11060 3334 11112 3340
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 11072 2990 11100 3334
rect 11152 3120 11204 3126
rect 11152 3062 11204 3068
rect 10324 2984 10376 2990
rect 10324 2926 10376 2932
rect 11060 2984 11112 2990
rect 11060 2926 11112 2932
rect 11072 2650 11100 2926
rect 11164 2650 11192 3062
rect 12268 3058 12296 3334
rect 12912 3126 12940 3402
rect 13280 3194 13308 3674
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 12256 3052 12308 3058
rect 12256 2994 12308 3000
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 9220 2644 9272 2650
rect 9220 2586 9272 2592
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 11808 2514 11836 2790
rect 11992 2774 12020 2994
rect 11992 2746 12112 2774
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 940 2440 992 2446
rect 2044 2440 2096 2446
rect 940 2382 992 2388
rect 1964 2400 2044 2428
rect 952 800 980 2382
rect 1964 800 1992 2400
rect 3056 2440 3108 2446
rect 2044 2382 2096 2388
rect 2976 2400 3056 2428
rect 2976 800 3004 2400
rect 4068 2440 4120 2446
rect 3056 2382 3108 2388
rect 3988 2400 4068 2428
rect 3988 800 4016 2400
rect 4068 2382 4120 2388
rect 4804 2440 4856 2446
rect 5080 2440 5132 2446
rect 4804 2382 4856 2388
rect 5000 2400 5080 2428
rect 5000 800 5028 2400
rect 5080 2382 5132 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 7012 2440 7064 2446
rect 8300 2440 8352 2446
rect 7012 2382 7064 2388
rect 8036 2400 8300 2428
rect 6012 800 6040 2382
rect 7024 800 7052 2382
rect 8036 800 8064 2400
rect 9128 2440 9180 2446
rect 8300 2382 8352 2388
rect 9048 2400 9128 2428
rect 9048 800 9076 2400
rect 9128 2382 9180 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 11060 2440 11112 2446
rect 11060 2382 11112 2388
rect 10060 800 10088 2382
rect 11072 800 11100 2382
rect 12084 800 12112 2746
rect 13096 800 13124 2994
rect 13280 2446 13308 3130
rect 13464 2774 13492 5646
rect 13740 5234 13768 6258
rect 14200 5914 14228 6734
rect 14476 6662 14504 11698
rect 14660 11218 14688 13144
rect 14740 13126 14792 13132
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14740 12708 14792 12714
rect 14740 12650 14792 12656
rect 14752 12238 14780 12650
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14832 11552 14884 11558
rect 14832 11494 14884 11500
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14844 11150 14872 11494
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 10674 14872 10950
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14568 8974 14596 10202
rect 14740 9104 14792 9110
rect 14740 9046 14792 9052
rect 14556 8968 14608 8974
rect 14556 8910 14608 8916
rect 14752 8838 14780 9046
rect 14844 9042 14872 10610
rect 14936 10062 14964 13330
rect 15014 12744 15070 12753
rect 15014 12679 15016 12688
rect 15068 12679 15070 12688
rect 15016 12650 15068 12656
rect 15120 12442 15148 15438
rect 15476 15428 15528 15434
rect 15476 15370 15528 15376
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15212 14006 15240 15030
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15304 14414 15332 14758
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15212 12986 15240 13942
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15200 12776 15252 12782
rect 15200 12718 15252 12724
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15016 12232 15068 12238
rect 15068 12180 15148 12186
rect 15016 12174 15148 12180
rect 15028 12158 15148 12174
rect 15120 11694 15148 12158
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 15028 9042 15056 11290
rect 15120 11132 15148 11630
rect 15212 11558 15240 12718
rect 15304 12434 15332 13806
rect 15384 13252 15436 13258
rect 15384 13194 15436 13200
rect 15396 12986 15424 13194
rect 15488 12986 15516 15370
rect 15844 15088 15896 15094
rect 15844 15030 15896 15036
rect 15660 14612 15712 14618
rect 15660 14554 15712 14560
rect 15672 13870 15700 14554
rect 15856 14414 15884 15030
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16040 14414 16068 14758
rect 16120 14544 16172 14550
rect 16120 14486 16172 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15752 14340 15804 14346
rect 15752 14282 15804 14288
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15384 12980 15436 12986
rect 15384 12922 15436 12928
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15476 12708 15528 12714
rect 15476 12650 15528 12656
rect 15304 12406 15424 12434
rect 15200 11552 15252 11558
rect 15200 11494 15252 11500
rect 15200 11144 15252 11150
rect 15120 11104 15200 11132
rect 15200 11086 15252 11092
rect 15212 9674 15240 11086
rect 15396 10606 15424 12406
rect 15488 12374 15516 12650
rect 15476 12368 15528 12374
rect 15476 12310 15528 12316
rect 15476 11212 15528 11218
rect 15476 11154 15528 11160
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10266 15424 10542
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15120 9646 15240 9674
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14568 6186 14596 8774
rect 14660 8634 14688 8774
rect 14752 8634 14780 8774
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14752 7886 14780 8570
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14752 7410 14780 7686
rect 14740 7404 14792 7410
rect 14740 7346 14792 7352
rect 14844 7290 14872 8978
rect 15028 8498 15056 8978
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15120 8430 15148 9646
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15108 8424 15160 8430
rect 15108 8366 15160 8372
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15120 7410 15148 7890
rect 15212 7886 15240 8842
rect 15396 8634 15424 9522
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8356 15344 8362
rect 15292 8298 15344 8304
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14752 7262 14872 7290
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14752 6390 14780 7262
rect 14832 7200 14884 7206
rect 14832 7142 14884 7148
rect 14844 6458 14872 7142
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14740 6384 14792 6390
rect 14740 6326 14792 6332
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14188 5908 14240 5914
rect 14188 5850 14240 5856
rect 14752 5710 14780 6326
rect 14832 6180 14884 6186
rect 14832 6122 14884 6128
rect 14844 5710 14872 6122
rect 14936 5914 14964 7278
rect 15120 6458 15148 7346
rect 15304 7290 15332 8298
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7478 15424 7686
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15304 7262 15424 7290
rect 15292 7200 15344 7206
rect 15292 7142 15344 7148
rect 15304 6458 15332 7142
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15396 5914 15424 7262
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 14740 5704 14792 5710
rect 14740 5646 14792 5652
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5370 15240 5646
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13556 3126 13584 5170
rect 13740 4622 13768 5170
rect 14740 5024 14792 5030
rect 14740 4966 14792 4972
rect 14752 4622 14780 4966
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 14108 3534 14136 4014
rect 14372 3936 14424 3942
rect 14372 3878 14424 3884
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14004 3460 14056 3466
rect 14004 3402 14056 3408
rect 13544 3120 13596 3126
rect 13544 3062 13596 3068
rect 13464 2746 13584 2774
rect 13556 2514 13584 2746
rect 14016 2650 14044 3402
rect 14108 2990 14136 3470
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14108 2582 14136 2926
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 14108 800 14136 2382
rect 14384 2310 14412 3878
rect 14476 2650 14504 4490
rect 15396 4162 15424 5850
rect 15488 5370 15516 11154
rect 15580 9654 15608 11154
rect 15672 11098 15700 13806
rect 15764 12152 15792 14282
rect 15856 13326 15884 14350
rect 15948 13802 15976 14350
rect 15936 13796 15988 13802
rect 15936 13738 15988 13744
rect 15844 13320 15896 13326
rect 15844 13262 15896 13268
rect 15948 12850 15976 13738
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15856 12374 15884 12786
rect 15948 12753 15976 12786
rect 15934 12744 15990 12753
rect 15934 12679 15990 12688
rect 15844 12368 15896 12374
rect 15844 12310 15896 12316
rect 15844 12164 15896 12170
rect 15764 12124 15844 12152
rect 15844 12106 15896 12112
rect 15672 11070 15792 11098
rect 15764 11014 15792 11070
rect 15752 11008 15804 11014
rect 15856 10985 15884 12106
rect 15752 10950 15804 10956
rect 15842 10976 15898 10985
rect 15660 10532 15712 10538
rect 15660 10474 15712 10480
rect 15672 10130 15700 10474
rect 15660 10124 15712 10130
rect 15660 10066 15712 10072
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15764 9382 15792 10950
rect 15842 10911 15898 10920
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15856 9518 15884 9658
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 9178 15792 9318
rect 15856 9178 15884 9454
rect 15752 9172 15804 9178
rect 15752 9114 15804 9120
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15580 6458 15608 8570
rect 15672 8430 15700 8910
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15948 7002 15976 12679
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16040 11830 16068 12242
rect 16028 11824 16080 11830
rect 16028 11766 16080 11772
rect 16132 11218 16160 14486
rect 16316 13394 16344 16594
rect 16684 15502 16712 17206
rect 16868 17202 16896 17274
rect 16960 17202 16988 17598
rect 17052 17338 17080 17614
rect 17040 17332 17092 17338
rect 17040 17274 17092 17280
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16868 15978 16896 17138
rect 17144 17134 17172 17614
rect 17972 17270 18000 17682
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 16948 16992 17000 16998
rect 16948 16934 17000 16940
rect 16960 16590 16988 16934
rect 16948 16584 17000 16590
rect 16948 16526 17000 16532
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16672 15496 16724 15502
rect 16672 15438 16724 15444
rect 16764 15496 16816 15502
rect 16764 15438 16816 15444
rect 16776 14618 16804 15438
rect 17144 15162 17172 17070
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17420 15162 17448 15982
rect 17592 15496 17644 15502
rect 17592 15438 17644 15444
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 17408 15156 17460 15162
rect 17408 15098 17460 15104
rect 17604 15026 17632 15438
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 16764 14612 16816 14618
rect 16764 14554 16816 14560
rect 16960 14074 16988 14962
rect 17512 14618 17540 14962
rect 17500 14612 17552 14618
rect 17500 14554 17552 14560
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 17696 14006 17724 16662
rect 17960 16108 18012 16114
rect 17960 16050 18012 16056
rect 17972 15706 18000 16050
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18064 15026 18092 18770
rect 18248 18766 18276 19110
rect 18524 18834 18552 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 20076 18896 20128 18902
rect 20076 18838 20128 18844
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18432 18358 18460 18566
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18426 20024 18702
rect 20088 18426 20116 18838
rect 20628 18760 20680 18766
rect 20628 18702 20680 18708
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 19984 18420 20036 18426
rect 19984 18362 20036 18368
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 18420 18352 18472 18358
rect 18420 18294 18472 18300
rect 20364 18290 20392 18566
rect 20640 18426 20668 18702
rect 21008 18698 21036 18838
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20812 18624 20864 18630
rect 20812 18566 20864 18572
rect 20904 18624 20956 18630
rect 20904 18566 20956 18572
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20824 18358 20852 18566
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 18328 18216 18380 18222
rect 18328 18158 18380 18164
rect 18340 17678 18368 18158
rect 18524 17746 18552 18226
rect 18696 18080 18748 18086
rect 18696 18022 18748 18028
rect 18512 17740 18564 17746
rect 18512 17682 18564 17688
rect 18328 17672 18380 17678
rect 18248 17632 18328 17660
rect 18248 17338 18276 17632
rect 18328 17614 18380 17620
rect 18420 17672 18472 17678
rect 18420 17614 18472 17620
rect 18432 17542 18460 17614
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18340 16046 18368 17478
rect 18432 17066 18460 17478
rect 18420 17060 18472 17066
rect 18420 17002 18472 17008
rect 18524 16998 18552 17682
rect 18708 17678 18736 18022
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18892 17338 18920 17682
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18984 17542 19012 17614
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19076 17338 19104 17478
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 18880 17332 18932 17338
rect 18880 17274 18932 17280
rect 19064 17332 19116 17338
rect 19064 17274 19116 17280
rect 19996 17202 20024 17478
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16114 19288 16594
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20456 16114 20484 18294
rect 20916 17218 20944 18566
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 20916 17202 21220 17218
rect 20904 17196 21232 17202
rect 20956 17190 21180 17196
rect 20904 17138 20956 17144
rect 21180 17138 21232 17144
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19800 16108 19852 16114
rect 19800 16050 19852 16056
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 19432 15904 19484 15910
rect 19432 15846 19484 15852
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 17880 14618 17908 14962
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17972 14346 18000 14758
rect 18064 14618 18092 14962
rect 19444 14958 19472 15846
rect 19812 15706 19840 16050
rect 20076 16040 20128 16046
rect 20076 15982 20128 15988
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 20088 15026 20116 15982
rect 20732 15978 20760 16050
rect 20720 15972 20772 15978
rect 20720 15914 20772 15920
rect 20916 15502 20944 16934
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21008 16250 21036 16526
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21008 15706 21036 16050
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21192 15502 21220 16934
rect 21364 16516 21416 16522
rect 21364 16458 21416 16464
rect 21376 16114 21404 16458
rect 21364 16108 21416 16114
rect 21364 16050 21416 16056
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 20916 15094 20944 15438
rect 21192 15162 21220 15438
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19984 14884 20036 14890
rect 19984 14826 20036 14832
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 17960 14340 18012 14346
rect 17960 14282 18012 14288
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 16304 13388 16356 13394
rect 16304 13330 16356 13336
rect 16396 13320 16448 13326
rect 16396 13262 16448 13268
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 16408 12442 16436 13262
rect 16684 12986 16712 13262
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16672 12980 16724 12986
rect 16672 12922 16724 12928
rect 16672 12708 16724 12714
rect 16672 12650 16724 12656
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16592 12374 16620 12582
rect 16580 12368 16632 12374
rect 16580 12310 16632 12316
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16224 11744 16252 12174
rect 16304 11756 16356 11762
rect 16224 11716 16304 11744
rect 16304 11698 16356 11704
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16316 11150 16344 11698
rect 16408 11354 16436 12174
rect 16592 12170 16620 12310
rect 16684 12238 16712 12650
rect 16776 12442 16804 13194
rect 17328 12850 17356 13262
rect 17604 12918 17632 13262
rect 17696 13190 17724 13942
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17592 12912 17644 12918
rect 17592 12854 17644 12860
rect 17224 12844 17276 12850
rect 17224 12786 17276 12792
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 16856 12776 16908 12782
rect 16856 12718 16908 12724
rect 16764 12436 16816 12442
rect 16764 12378 16816 12384
rect 16868 12238 16896 12718
rect 17236 12434 17264 12786
rect 17052 12406 17264 12434
rect 16672 12232 16724 12238
rect 16672 12174 16724 12180
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16948 12232 17000 12238
rect 17052 12220 17080 12406
rect 17000 12192 17080 12220
rect 17132 12232 17184 12238
rect 16948 12174 17000 12180
rect 17328 12220 17356 12786
rect 17972 12782 18000 13738
rect 18156 13258 18184 14350
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 18604 13796 18656 13802
rect 18604 13738 18656 13744
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18616 13394 18644 13738
rect 18604 13388 18656 13394
rect 18604 13330 18656 13336
rect 18144 13252 18196 13258
rect 18144 13194 18196 13200
rect 18328 13252 18380 13258
rect 18328 13194 18380 13200
rect 18420 13252 18472 13258
rect 18420 13194 18472 13200
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17184 12192 17356 12220
rect 17408 12232 17460 12238
rect 17132 12174 17184 12180
rect 17408 12174 17460 12180
rect 16580 12164 16632 12170
rect 16580 12106 16632 12112
rect 16868 11558 16896 12174
rect 17420 11898 17448 12174
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11898 17632 12038
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16396 11348 16448 11354
rect 16396 11290 16448 11296
rect 16304 11144 16356 11150
rect 16304 11086 16356 11092
rect 16672 11076 16724 11082
rect 16672 11018 16724 11024
rect 16028 11008 16080 11014
rect 16028 10950 16080 10956
rect 16212 11008 16264 11014
rect 16212 10950 16264 10956
rect 16040 10742 16068 10950
rect 16224 10810 16252 10950
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16028 10736 16080 10742
rect 16028 10678 16080 10684
rect 16040 10266 16068 10678
rect 16120 10464 16172 10470
rect 16120 10406 16172 10412
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16040 10062 16068 10202
rect 16132 10062 16160 10406
rect 16224 10062 16252 10746
rect 16396 10464 16448 10470
rect 16396 10406 16448 10412
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16212 10056 16264 10062
rect 16212 9998 16264 10004
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16316 8974 16344 9998
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 16040 6866 16068 7482
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16132 6662 16160 7346
rect 16316 7274 16344 8910
rect 16408 7546 16436 10406
rect 16684 9518 16712 11018
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17328 10266 17356 10542
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 9654 17632 9862
rect 17592 9648 17644 9654
rect 17592 9590 17644 9596
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 17696 8974 17724 10474
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17788 10062 17816 10406
rect 18340 10266 18368 13194
rect 18432 11694 18460 13194
rect 18984 13190 19012 13738
rect 18972 13184 19024 13190
rect 18972 13126 19024 13132
rect 19352 12918 19380 13874
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 18972 12844 19024 12850
rect 18972 12786 19024 12792
rect 18984 12434 19012 12786
rect 19444 12714 19472 13874
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19904 13326 19932 13806
rect 19996 13682 20024 14826
rect 20088 14074 20116 14962
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20732 13938 20760 14962
rect 20812 14884 20864 14890
rect 20812 14826 20864 14832
rect 20824 14414 20852 14826
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14482 21496 14758
rect 21456 14476 21508 14482
rect 21548 14476 21600 14482
rect 21508 14436 21548 14464
rect 21456 14418 21508 14424
rect 21548 14418 21600 14424
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14074 20852 14350
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 21192 13734 21220 14214
rect 21284 13938 21312 14214
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21180 13728 21232 13734
rect 19996 13654 20208 13682
rect 21180 13670 21232 13676
rect 19984 13388 20036 13394
rect 19984 13330 20036 13336
rect 19892 13320 19944 13326
rect 19892 13262 19944 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19996 12986 20024 13330
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19432 12708 19484 12714
rect 19432 12650 19484 12656
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 18708 12406 19012 12434
rect 18708 12170 18736 12406
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18696 12164 18748 12170
rect 18696 12106 18748 12112
rect 18708 11898 18736 12106
rect 18800 11898 18828 12174
rect 18696 11892 18748 11898
rect 18696 11834 18748 11840
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18892 11694 18920 12174
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18880 11688 18932 11694
rect 18880 11630 18932 11636
rect 18512 11144 18564 11150
rect 19352 11132 19380 12582
rect 20088 12442 20116 13262
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19444 11354 19472 12174
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19996 11898 20024 12038
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19616 11552 19668 11558
rect 19616 11494 19668 11500
rect 20076 11552 20128 11558
rect 20076 11494 20128 11500
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19536 11286 19564 11494
rect 19628 11354 19656 11494
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19524 11144 19576 11150
rect 19352 11104 19524 11132
rect 18512 11086 18564 11092
rect 19524 11086 19576 11092
rect 18328 10260 18380 10266
rect 18328 10202 18380 10208
rect 17880 10130 18276 10146
rect 17880 10124 18288 10130
rect 17880 10118 18236 10124
rect 17776 10056 17828 10062
rect 17776 9998 17828 10004
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 16764 8832 16816 8838
rect 16764 8774 16816 8780
rect 16856 8832 16908 8838
rect 16856 8774 16908 8780
rect 16776 8498 16804 8774
rect 16868 8498 16896 8774
rect 17500 8560 17552 8566
rect 17500 8502 17552 8508
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16304 7268 16356 7274
rect 16304 7210 16356 7216
rect 16316 6798 16344 7210
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6474 16160 6598
rect 16040 6458 16160 6474
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 16028 6452 16160 6458
rect 16080 6446 16160 6452
rect 16028 6394 16080 6400
rect 15580 5710 15608 6394
rect 16132 6236 16160 6446
rect 16212 6384 16264 6390
rect 16316 6372 16344 6734
rect 16264 6344 16344 6372
rect 16212 6326 16264 6332
rect 16132 6208 16344 6236
rect 15936 6180 15988 6186
rect 15936 6122 15988 6128
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15948 5234 15976 6122
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5234 16252 6054
rect 16316 5234 16344 6208
rect 16408 6118 16436 7482
rect 17512 7410 17540 8502
rect 17604 7886 17632 8842
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 7478 17632 7822
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17604 6798 17632 7414
rect 17788 7002 17816 9998
rect 17880 9518 17908 10118
rect 18236 10066 18288 10072
rect 18052 9988 18104 9994
rect 18052 9930 18104 9936
rect 17868 9512 17920 9518
rect 17868 9454 17920 9460
rect 17960 9376 18012 9382
rect 18064 9364 18092 9930
rect 18340 9722 18368 10202
rect 18524 10062 18552 11086
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19340 10192 19392 10198
rect 19340 10134 19392 10140
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18524 9586 18552 9998
rect 18880 9920 18932 9926
rect 18880 9862 18932 9868
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18012 9336 18092 9364
rect 17960 9318 18012 9324
rect 18892 8634 18920 9862
rect 19352 9586 19380 10134
rect 19904 10062 19932 10406
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19904 9926 19932 9998
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 19432 9376 19484 9382
rect 19432 9318 19484 9324
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18708 7886 18736 8434
rect 18892 7954 18920 8434
rect 18984 7954 19012 8434
rect 18880 7948 18932 7954
rect 18880 7890 18932 7896
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 17972 7342 18000 7822
rect 18328 7744 18380 7750
rect 18328 7686 18380 7692
rect 18340 7478 18368 7686
rect 18984 7546 19012 7890
rect 18972 7540 19024 7546
rect 18972 7482 19024 7488
rect 18328 7472 18380 7478
rect 18328 7414 18380 7420
rect 17960 7336 18012 7342
rect 17960 7278 18012 7284
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 18340 6798 18368 7414
rect 18420 7404 18472 7410
rect 18420 7346 18472 7352
rect 18432 6866 18460 7346
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 16488 6724 16540 6730
rect 16488 6666 16540 6672
rect 17684 6724 17736 6730
rect 17684 6666 17736 6672
rect 16500 6322 16528 6666
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16488 6316 16540 6322
rect 16488 6258 16540 6264
rect 16592 6186 16620 6598
rect 17408 6384 17460 6390
rect 17408 6326 17460 6332
rect 16580 6180 16632 6186
rect 16580 6122 16632 6128
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 17420 5914 17448 6326
rect 17696 6254 17724 6666
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17788 6322 17816 6598
rect 18340 6458 18368 6734
rect 19352 6458 19380 6802
rect 19444 6798 19472 9318
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19996 8634 20024 9454
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20088 8514 20116 11494
rect 20180 10010 20208 13654
rect 21192 13326 21220 13670
rect 21180 13320 21232 13326
rect 21180 13262 21232 13268
rect 21284 13258 21312 13874
rect 21272 13252 21324 13258
rect 21272 13194 21324 13200
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 20812 11552 20864 11558
rect 20812 11494 20864 11500
rect 20444 11280 20496 11286
rect 20444 11222 20496 11228
rect 20180 9994 20300 10010
rect 20180 9988 20312 9994
rect 20180 9982 20260 9988
rect 20260 9930 20312 9936
rect 19904 8486 20116 8514
rect 19904 7886 19932 8486
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 19996 8090 20024 8366
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19996 7342 20024 8026
rect 20180 8022 20208 8366
rect 20168 8016 20220 8022
rect 20168 7958 20220 7964
rect 20180 7886 20208 7958
rect 20456 7954 20484 11222
rect 20536 10056 20588 10062
rect 20536 9998 20588 10004
rect 20548 9722 20576 9998
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20548 8498 20576 9522
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20444 7948 20496 7954
rect 20444 7890 20496 7896
rect 20168 7880 20220 7886
rect 20168 7822 20220 7828
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19984 7336 20036 7342
rect 19984 7278 20036 7284
rect 20180 6798 20208 7822
rect 20260 7744 20312 7750
rect 20260 7686 20312 7692
rect 20272 7546 20300 7686
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20364 6798 20392 7822
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 20352 6792 20404 6798
rect 20352 6734 20404 6740
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17684 6248 17736 6254
rect 17684 6190 17736 6196
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17972 5914 18000 6122
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 18156 5914 18184 6054
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 18340 5710 18368 6394
rect 19444 6322 19472 6734
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19996 5710 20024 6598
rect 20364 6458 20392 6734
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20456 5778 20484 7890
rect 20548 7750 20576 8434
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7546 20576 7686
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20548 7274 20576 7482
rect 20640 7478 20668 7822
rect 20824 7546 20852 11494
rect 21192 9654 21220 13126
rect 21652 12434 21680 18158
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 22100 17060 22152 17066
rect 22100 17002 22152 17008
rect 22112 16726 22140 17002
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 22100 16720 22152 16726
rect 22152 16680 22232 16708
rect 22100 16662 22152 16668
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22008 16516 22060 16522
rect 22008 16458 22060 16464
rect 22020 16182 22048 16458
rect 22112 16250 22140 16526
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22008 16176 22060 16182
rect 22008 16118 22060 16124
rect 22100 16040 22152 16046
rect 22204 16028 22232 16680
rect 26056 16448 26108 16454
rect 26056 16390 26108 16396
rect 26068 16182 26096 16390
rect 26056 16176 26108 16182
rect 26056 16118 26108 16124
rect 26976 16176 27028 16182
rect 26976 16118 27028 16124
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 22152 16000 22232 16028
rect 22100 15982 22152 15988
rect 23308 15706 23336 16050
rect 24308 15972 24360 15978
rect 24308 15914 24360 15920
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 23296 15700 23348 15706
rect 23296 15642 23348 15648
rect 21824 15496 21876 15502
rect 21824 15438 21876 15444
rect 21836 15026 21864 15438
rect 21824 15020 21876 15026
rect 21824 14962 21876 14968
rect 21652 12406 21772 12434
rect 21640 11756 21692 11762
rect 21640 11698 21692 11704
rect 21652 10810 21680 11698
rect 21744 11694 21772 12406
rect 21732 11688 21784 11694
rect 21732 11630 21784 11636
rect 21836 10810 21864 14962
rect 22112 14618 22140 15642
rect 23940 14884 23992 14890
rect 23940 14826 23992 14832
rect 23952 14618 23980 14826
rect 22100 14612 22152 14618
rect 22100 14554 22152 14560
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23940 14612 23992 14618
rect 23940 14554 23992 14560
rect 22192 14544 22244 14550
rect 22192 14486 22244 14492
rect 21916 14340 21968 14346
rect 21916 14282 21968 14288
rect 21928 14074 21956 14282
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21928 13462 21956 13874
rect 22100 13864 22152 13870
rect 22100 13806 22152 13812
rect 21916 13456 21968 13462
rect 21916 13398 21968 13404
rect 21928 12782 21956 13398
rect 22112 13258 22140 13806
rect 22100 13252 22152 13258
rect 22100 13194 22152 13200
rect 21916 12776 21968 12782
rect 21916 12718 21968 12724
rect 22204 12714 22232 14486
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 12918 22324 14214
rect 22388 14006 22416 14282
rect 23032 14278 23060 14350
rect 23020 14272 23072 14278
rect 23020 14214 23072 14220
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22376 14000 22428 14006
rect 22376 13942 22428 13948
rect 22480 13258 22508 14010
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22284 12912 22336 12918
rect 22284 12854 22336 12860
rect 22192 12708 22244 12714
rect 22192 12650 22244 12656
rect 22204 12238 22232 12650
rect 22296 12442 22324 12854
rect 22284 12436 22336 12442
rect 22284 12378 22336 12384
rect 22192 12232 22244 12238
rect 22192 12174 22244 12180
rect 22572 12170 22600 13806
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22664 12238 22692 12582
rect 22652 12232 22704 12238
rect 22652 12174 22704 12180
rect 22560 12164 22612 12170
rect 22560 12106 22612 12112
rect 22572 11762 22600 12106
rect 22560 11756 22612 11762
rect 22560 11698 22612 11704
rect 22468 11552 22520 11558
rect 22468 11494 22520 11500
rect 21640 10804 21692 10810
rect 21640 10746 21692 10752
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 22480 10674 22508 11494
rect 22940 10674 22968 13126
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 22100 10668 22152 10674
rect 22100 10610 22152 10616
rect 22468 10668 22520 10674
rect 22468 10610 22520 10616
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21284 10266 21312 10406
rect 21272 10260 21324 10266
rect 21272 10202 21324 10208
rect 21376 9926 21404 10610
rect 21468 10198 21496 10610
rect 21916 10600 21968 10606
rect 21916 10542 21968 10548
rect 21456 10192 21508 10198
rect 21456 10134 21508 10140
rect 21928 10062 21956 10542
rect 22112 10198 22140 10610
rect 22940 10266 22968 10610
rect 22928 10260 22980 10266
rect 22928 10202 22980 10208
rect 22100 10192 22152 10198
rect 22100 10134 22152 10140
rect 22112 10062 22140 10134
rect 21916 10056 21968 10062
rect 21916 9998 21968 10004
rect 22100 10056 22152 10062
rect 22100 9998 22152 10004
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 20996 9512 21048 9518
rect 20996 9454 21048 9460
rect 21008 8974 21036 9454
rect 21192 9110 21220 9590
rect 21376 9178 21404 9862
rect 21928 9722 21956 9998
rect 22112 9926 22140 9998
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 22284 9920 22336 9926
rect 22284 9862 22336 9868
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22296 9722 22324 9862
rect 22756 9722 22784 9862
rect 21916 9716 21968 9722
rect 21916 9658 21968 9664
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22744 9716 22796 9722
rect 22744 9658 22796 9664
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21180 9104 21232 9110
rect 21180 9046 21232 9052
rect 21192 8974 21220 9046
rect 21928 8974 21956 9658
rect 23032 9654 23060 14214
rect 23112 14068 23164 14074
rect 23112 14010 23164 14016
rect 23124 13938 23152 14010
rect 23112 13932 23164 13938
rect 23112 13874 23164 13880
rect 23124 13530 23152 13874
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 23112 13524 23164 13530
rect 23112 13466 23164 13472
rect 23308 13326 23336 13670
rect 23400 13462 23428 14418
rect 23572 14408 23624 14414
rect 23492 14368 23572 14396
rect 23492 13870 23520 14368
rect 23572 14350 23624 14356
rect 23676 14074 23704 14554
rect 23664 14068 23716 14074
rect 23664 14010 23716 14016
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 23492 13530 23520 13806
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23388 13456 23440 13462
rect 23388 13398 23440 13404
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23216 13190 23244 13262
rect 23204 13184 23256 13190
rect 23204 13126 23256 13132
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23112 12232 23164 12238
rect 23112 12174 23164 12180
rect 23124 11898 23152 12174
rect 23216 11898 23244 12242
rect 23112 11892 23164 11898
rect 23112 11834 23164 11840
rect 23204 11892 23256 11898
rect 23204 11834 23256 11840
rect 23308 10810 23336 13262
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23308 10198 23336 10746
rect 23296 10192 23348 10198
rect 23296 10134 23348 10140
rect 23296 9988 23348 9994
rect 23296 9930 23348 9936
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 21180 8968 21232 8974
rect 21180 8910 21232 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21916 8968 21968 8974
rect 21916 8910 21968 8916
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21192 7886 21220 8774
rect 21468 7954 21496 8910
rect 22192 8832 22244 8838
rect 22192 8774 22244 8780
rect 21456 7948 21508 7954
rect 21456 7890 21508 7896
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20628 7472 20680 7478
rect 20628 7414 20680 7420
rect 20536 7268 20588 7274
rect 20536 7210 20588 7216
rect 20824 6798 20852 7482
rect 20916 7478 20944 7822
rect 21088 7744 21140 7750
rect 21088 7686 21140 7692
rect 20904 7472 20956 7478
rect 21100 7426 21128 7686
rect 20904 7414 20956 7420
rect 21008 7410 21128 7426
rect 20996 7404 21128 7410
rect 21048 7398 21128 7404
rect 20996 7346 21048 7352
rect 21100 6866 21128 7398
rect 21192 7002 21220 7822
rect 21272 7744 21324 7750
rect 21272 7686 21324 7692
rect 21180 6996 21232 7002
rect 21180 6938 21232 6944
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 21284 5914 21312 7686
rect 21376 7546 21404 7822
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21836 7546 21864 7686
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21376 6798 21404 7278
rect 22204 7274 22232 8774
rect 22192 7268 22244 7274
rect 22192 7210 22244 7216
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 21272 5908 21324 5914
rect 21272 5850 21324 5856
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 21364 5772 21416 5778
rect 21364 5714 21416 5720
rect 18328 5704 18380 5710
rect 18328 5646 18380 5652
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 20076 5636 20128 5642
rect 20076 5578 20128 5584
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16028 5024 16080 5030
rect 16028 4966 16080 4972
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15948 4282 15976 4490
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 15396 4146 15516 4162
rect 15396 4140 15528 4146
rect 15396 4134 15476 4140
rect 15476 4082 15528 4088
rect 14464 2644 14516 2650
rect 14464 2586 14516 2592
rect 15488 2514 15516 4082
rect 16040 4010 16068 4966
rect 16316 4826 16344 4966
rect 16592 4826 16620 5238
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17144 4826 17172 4966
rect 18248 4826 18276 5510
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19996 5234 20024 5510
rect 20088 5234 20116 5578
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 21376 5030 21404 5714
rect 22388 5234 22416 7142
rect 22480 5778 22508 9318
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7546 23060 8230
rect 23308 8090 23336 9930
rect 23400 9382 23428 13398
rect 23572 12096 23624 12102
rect 23572 12038 23624 12044
rect 23584 11898 23612 12038
rect 23572 11892 23624 11898
rect 23572 11834 23624 11840
rect 23756 11552 23808 11558
rect 23756 11494 23808 11500
rect 23572 10464 23624 10470
rect 23572 10406 23624 10412
rect 23584 10130 23612 10406
rect 23572 10124 23624 10130
rect 23572 10066 23624 10072
rect 23480 9512 23532 9518
rect 23480 9454 23532 9460
rect 23388 9376 23440 9382
rect 23388 9318 23440 9324
rect 23492 9178 23520 9454
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23584 8498 23612 10066
rect 23664 9104 23716 9110
rect 23664 9046 23716 9052
rect 23676 8634 23704 9046
rect 23664 8628 23716 8634
rect 23664 8570 23716 8576
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23676 7954 23704 8570
rect 23664 7948 23716 7954
rect 23664 7890 23716 7896
rect 23020 7540 23072 7546
rect 23020 7482 23072 7488
rect 23676 7274 23704 7890
rect 23664 7268 23716 7274
rect 23664 7210 23716 7216
rect 23676 7002 23704 7210
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23768 5914 23796 11494
rect 23848 10600 23900 10606
rect 23848 10542 23900 10548
rect 23860 10266 23888 10542
rect 23952 10538 23980 14554
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 13938 24164 14214
rect 24032 13932 24084 13938
rect 24032 13874 24084 13880
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24044 13682 24072 13874
rect 24136 13818 24164 13874
rect 24136 13790 24256 13818
rect 24044 13654 24164 13682
rect 24032 13320 24084 13326
rect 24032 13262 24084 13268
rect 24044 10538 24072 13262
rect 24136 13190 24164 13654
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 24032 10532 24084 10538
rect 24032 10474 24084 10480
rect 23848 10260 23900 10266
rect 23848 10202 23900 10208
rect 23952 10062 23980 10474
rect 24136 10266 24164 13126
rect 24124 10260 24176 10266
rect 24124 10202 24176 10208
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23940 9580 23992 9586
rect 23940 9522 23992 9528
rect 23860 9382 23888 9522
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23952 8838 23980 9522
rect 24136 9450 24164 10202
rect 24228 9586 24256 13790
rect 24320 12238 24348 15914
rect 24688 15502 24716 16050
rect 24872 15570 24900 16050
rect 25688 16040 25740 16046
rect 25688 15982 25740 15988
rect 25700 15706 25728 15982
rect 26068 15706 26096 16118
rect 26516 15904 26568 15910
rect 26516 15846 26568 15852
rect 26528 15706 26556 15846
rect 25688 15700 25740 15706
rect 25688 15642 25740 15648
rect 26056 15700 26108 15706
rect 26056 15642 26108 15648
rect 26516 15700 26568 15706
rect 26516 15642 26568 15648
rect 26988 15570 27016 16118
rect 28080 16040 28132 16046
rect 28080 15982 28132 15988
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 26976 15564 27028 15570
rect 26976 15506 27028 15512
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24872 14958 24900 15506
rect 27436 15496 27488 15502
rect 27488 15456 27568 15484
rect 27436 15438 27488 15444
rect 24860 14952 24912 14958
rect 24860 14894 24912 14900
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24400 14408 24452 14414
rect 24400 14350 24452 14356
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24860 14408 24912 14414
rect 24860 14350 24912 14356
rect 24412 14074 24440 14350
rect 24400 14068 24452 14074
rect 24400 14010 24452 14016
rect 24504 13818 24532 14350
rect 24412 13790 24532 13818
rect 24412 13394 24440 13790
rect 24492 13728 24544 13734
rect 24492 13670 24544 13676
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24504 13530 24532 13670
rect 24492 13524 24544 13530
rect 24492 13466 24544 13472
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24688 13258 24716 13670
rect 24872 13326 24900 14350
rect 25056 13326 25084 14418
rect 26056 14408 26108 14414
rect 26056 14350 26108 14356
rect 25320 14340 25372 14346
rect 25320 14282 25372 14288
rect 25332 14074 25360 14282
rect 25412 14272 25464 14278
rect 25412 14214 25464 14220
rect 25872 14272 25924 14278
rect 25872 14214 25924 14220
rect 25424 14074 25452 14214
rect 25884 14074 25912 14214
rect 25320 14068 25372 14074
rect 25320 14010 25372 14016
rect 25412 14068 25464 14074
rect 25412 14010 25464 14016
rect 25872 14068 25924 14074
rect 25872 14010 25924 14016
rect 25228 13932 25280 13938
rect 25228 13874 25280 13880
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 25240 13258 25268 13874
rect 25780 13864 25832 13870
rect 25780 13806 25832 13812
rect 25412 13728 25464 13734
rect 25412 13670 25464 13676
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 25228 13252 25280 13258
rect 25228 13194 25280 13200
rect 24768 13184 24820 13190
rect 24768 13126 24820 13132
rect 24780 12238 24808 13126
rect 24308 12232 24360 12238
rect 24308 12174 24360 12180
rect 24768 12232 24820 12238
rect 24768 12174 24820 12180
rect 24308 12096 24360 12102
rect 24308 12038 24360 12044
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24860 12096 24912 12102
rect 24860 12038 24912 12044
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24124 9444 24176 9450
rect 24124 9386 24176 9392
rect 24136 9178 24164 9386
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24228 8974 24256 9522
rect 24216 8968 24268 8974
rect 24216 8910 24268 8916
rect 23940 8832 23992 8838
rect 23940 8774 23992 8780
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23952 7886 23980 8434
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23860 7410 23888 7686
rect 23952 7546 23980 7822
rect 23940 7540 23992 7546
rect 23940 7482 23992 7488
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23952 6934 23980 7482
rect 23940 6928 23992 6934
rect 23940 6870 23992 6876
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23756 5908 23808 5914
rect 23756 5850 23808 5856
rect 22468 5772 22520 5778
rect 22468 5714 22520 5720
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 22928 5636 22980 5642
rect 22928 5578 22980 5584
rect 22940 5370 22968 5578
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 23032 5234 23060 5714
rect 22376 5228 22428 5234
rect 22376 5170 22428 5176
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 19984 5024 20036 5030
rect 19984 4966 20036 4972
rect 20812 5024 20864 5030
rect 20812 4966 20864 4972
rect 21364 5024 21416 5030
rect 21364 4966 21416 4972
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 19996 4826 20024 4966
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 16580 4820 16632 4826
rect 16580 4762 16632 4768
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 19984 4820 20036 4826
rect 19984 4762 20036 4768
rect 19432 4752 19484 4758
rect 19432 4694 19484 4700
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 18144 4480 18196 4486
rect 18144 4422 18196 4428
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15672 3738 15700 3878
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15580 2514 15608 3130
rect 16500 2774 16528 3334
rect 16592 3194 16620 3402
rect 16580 3188 16632 3194
rect 16580 3130 16632 3136
rect 16672 3120 16724 3126
rect 16672 3062 16724 3068
rect 16500 2746 16620 2774
rect 16592 2582 16620 2746
rect 16684 2582 16712 3062
rect 16776 2650 16804 4082
rect 16868 2650 16896 4422
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 2774 17264 4014
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 17880 3194 17908 3402
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17144 2746 17264 2774
rect 16764 2644 16816 2650
rect 16764 2586 16816 2592
rect 16856 2644 16908 2650
rect 16856 2586 16908 2592
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 16672 2440 16724 2446
rect 16500 2400 16672 2428
rect 14924 2372 14976 2378
rect 14924 2314 14976 2320
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14936 1306 14964 2314
rect 14936 1278 15148 1306
rect 15120 800 15148 1278
rect 16132 870 16252 898
rect 16132 800 16160 870
rect 938 0 994 800
rect 1950 0 2006 800
rect 2962 0 3018 800
rect 3974 0 4030 800
rect 4986 0 5042 800
rect 5998 0 6054 800
rect 7010 0 7066 800
rect 8022 0 8078 800
rect 9034 0 9090 800
rect 10046 0 10102 800
rect 11058 0 11114 800
rect 12070 0 12126 800
rect 13082 0 13138 800
rect 14094 0 14150 800
rect 15106 0 15162 800
rect 16118 0 16174 800
rect 16224 762 16252 870
rect 16500 762 16528 2400
rect 16672 2382 16724 2388
rect 17144 800 17172 2746
rect 17880 2378 17908 3130
rect 18156 3126 18184 4422
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18248 3738 18276 4082
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18144 3120 18196 3126
rect 18144 3062 18196 3068
rect 17868 2372 17920 2378
rect 17868 2314 17920 2320
rect 18156 870 18276 898
rect 18156 800 18184 870
rect 16224 734 16528 762
rect 17130 0 17186 800
rect 18142 0 18198 800
rect 18248 762 18276 870
rect 18432 762 18460 4014
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18708 2446 18736 3538
rect 19444 2922 19472 4694
rect 20824 4622 20852 4966
rect 21376 4690 21404 4966
rect 22020 4690 22048 4966
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 21364 4684 21416 4690
rect 21364 4626 21416 4632
rect 22008 4684 22060 4690
rect 22008 4626 22060 4632
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19892 3528 19944 3534
rect 19890 3496 19892 3505
rect 21824 3528 21876 3534
rect 19944 3496 19946 3505
rect 21824 3470 21876 3476
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 19890 3431 19946 3440
rect 21088 3460 21140 3466
rect 21088 3402 21140 3408
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 19800 2984 19852 2990
rect 20168 2984 20220 2990
rect 19852 2944 20168 2972
rect 19800 2926 19852 2932
rect 20168 2926 20220 2932
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 18696 2440 18748 2446
rect 18696 2382 18748 2388
rect 19352 1442 19380 2450
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19168 1414 19380 1442
rect 19168 800 19196 1414
rect 20272 1170 20300 2450
rect 21100 1714 21128 3402
rect 21836 2990 21864 3470
rect 21928 3194 21956 3470
rect 21916 3188 21968 3194
rect 21916 3130 21968 3136
rect 22112 3126 22140 4694
rect 22388 4690 22416 5170
rect 22376 4684 22428 4690
rect 22376 4626 22428 4632
rect 22468 4480 22520 4486
rect 22468 4422 22520 4428
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 21824 2984 21876 2990
rect 21824 2926 21876 2932
rect 21824 2848 21876 2854
rect 21824 2790 21876 2796
rect 21836 2446 21864 2790
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21100 1686 21220 1714
rect 20180 1142 20300 1170
rect 20180 800 20208 1142
rect 21192 800 21220 1686
rect 22204 800 22232 4014
rect 22480 3602 22508 4422
rect 23296 4072 23348 4078
rect 23296 4014 23348 4020
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22928 3460 22980 3466
rect 22928 3402 22980 3408
rect 22940 3194 22968 3402
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 23308 2122 23336 4014
rect 23492 3126 23520 5850
rect 23572 5772 23624 5778
rect 23572 5714 23624 5720
rect 23584 5234 23612 5714
rect 23572 5228 23624 5234
rect 23572 5170 23624 5176
rect 23768 5166 23796 5850
rect 24320 5794 24348 12038
rect 24596 11762 24624 12038
rect 24872 11898 24900 12038
rect 24860 11892 24912 11898
rect 24860 11834 24912 11840
rect 24584 11756 24636 11762
rect 24584 11698 24636 11704
rect 24872 11354 24900 11834
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25148 11354 25176 11698
rect 25320 11688 25372 11694
rect 25320 11630 25372 11636
rect 25332 11354 25360 11630
rect 24860 11348 24912 11354
rect 24860 11290 24912 11296
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25320 11076 25372 11082
rect 25320 11018 25372 11024
rect 25332 10810 25360 11018
rect 25320 10804 25372 10810
rect 25320 10746 25372 10752
rect 24676 10600 24728 10606
rect 24676 10542 24728 10548
rect 24492 10056 24544 10062
rect 24492 9998 24544 10004
rect 24584 10056 24636 10062
rect 24584 9998 24636 10004
rect 24504 9654 24532 9998
rect 24596 9722 24624 9998
rect 24584 9716 24636 9722
rect 24584 9658 24636 9664
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24504 8974 24532 9590
rect 24688 9586 24716 10542
rect 24860 10056 24912 10062
rect 24860 9998 24912 10004
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24688 9042 24716 9522
rect 24872 9382 24900 9998
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24676 9036 24728 9042
rect 24676 8978 24728 8984
rect 24492 8968 24544 8974
rect 24492 8910 24544 8916
rect 24584 8832 24636 8838
rect 24584 8774 24636 8780
rect 24596 8294 24624 8774
rect 24872 8498 24900 9318
rect 24964 9178 24992 9998
rect 25424 9450 25452 13670
rect 25792 13530 25820 13806
rect 26068 13530 26096 14350
rect 26976 13864 27028 13870
rect 26976 13806 27028 13812
rect 26424 13796 26476 13802
rect 26424 13738 26476 13744
rect 25780 13524 25832 13530
rect 25780 13466 25832 13472
rect 26056 13524 26108 13530
rect 26056 13466 26108 13472
rect 26332 13388 26384 13394
rect 26332 13330 26384 13336
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 25608 12434 25636 13262
rect 25780 12436 25832 12442
rect 25608 12406 25780 12434
rect 25780 12378 25832 12384
rect 26160 12238 26188 13262
rect 26344 12442 26372 13330
rect 26332 12436 26384 12442
rect 26332 12378 26384 12384
rect 25504 12232 25556 12238
rect 25504 12174 25556 12180
rect 26148 12232 26200 12238
rect 26148 12174 26200 12180
rect 26332 12232 26384 12238
rect 26332 12174 26384 12180
rect 25516 11762 25544 12174
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25608 11762 25636 12038
rect 25504 11756 25556 11762
rect 25504 11698 25556 11704
rect 25596 11756 25648 11762
rect 25596 11698 25648 11704
rect 25516 11150 25544 11698
rect 25608 11150 25636 11698
rect 26056 11688 26108 11694
rect 26056 11630 26108 11636
rect 25504 11144 25556 11150
rect 25504 11086 25556 11092
rect 25596 11144 25648 11150
rect 25596 11086 25648 11092
rect 25504 11008 25556 11014
rect 25504 10950 25556 10956
rect 25516 10266 25544 10950
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 25516 9518 25544 9862
rect 25504 9512 25556 9518
rect 25504 9454 25556 9460
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25780 9376 25832 9382
rect 25780 9318 25832 9324
rect 24952 9172 25004 9178
rect 24952 9114 25004 9120
rect 25240 8974 25268 9318
rect 25792 9178 25820 9318
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25228 8968 25280 8974
rect 25228 8910 25280 8916
rect 25240 8498 25268 8910
rect 25872 8832 25924 8838
rect 25872 8774 25924 8780
rect 24860 8492 24912 8498
rect 24860 8434 24912 8440
rect 25228 8492 25280 8498
rect 25228 8434 25280 8440
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 24584 8288 24636 8294
rect 24584 8230 24636 8236
rect 24596 7886 24624 8230
rect 24872 8022 24900 8434
rect 24952 8424 25004 8430
rect 25240 8378 25268 8434
rect 24952 8366 25004 8372
rect 24860 8016 24912 8022
rect 24860 7958 24912 7964
rect 24964 7886 24992 8366
rect 25148 8350 25268 8378
rect 25320 8356 25372 8362
rect 25148 8090 25176 8350
rect 25320 8298 25372 8304
rect 25228 8288 25280 8294
rect 25228 8230 25280 8236
rect 25136 8084 25188 8090
rect 25136 8026 25188 8032
rect 24584 7880 24636 7886
rect 24584 7822 24636 7828
rect 24952 7880 25004 7886
rect 24952 7822 25004 7828
rect 25240 7410 25268 8230
rect 25332 7818 25360 8298
rect 25688 8084 25740 8090
rect 25688 8026 25740 8032
rect 25700 7818 25728 8026
rect 25792 7886 25820 8434
rect 25884 8106 25912 8774
rect 25884 8090 26004 8106
rect 25884 8084 26016 8090
rect 25884 8078 25964 8084
rect 25780 7880 25832 7886
rect 25780 7822 25832 7828
rect 25320 7812 25372 7818
rect 25320 7754 25372 7760
rect 25688 7812 25740 7818
rect 25688 7754 25740 7760
rect 25884 7750 25912 8078
rect 25964 8026 26016 8032
rect 25964 7948 26016 7954
rect 25964 7890 26016 7896
rect 25872 7744 25924 7750
rect 25872 7686 25924 7692
rect 25976 7546 26004 7890
rect 25964 7540 26016 7546
rect 25964 7482 26016 7488
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24320 5766 24624 5794
rect 24124 5568 24176 5574
rect 24124 5510 24176 5516
rect 24136 5234 24164 5510
rect 24124 5228 24176 5234
rect 24124 5170 24176 5176
rect 24412 5166 24440 5766
rect 24596 5710 24624 5766
rect 24584 5704 24636 5710
rect 24584 5646 24636 5652
rect 25136 5568 25188 5574
rect 25136 5510 25188 5516
rect 25148 5234 25176 5510
rect 26068 5370 26096 11630
rect 26160 11354 26188 12174
rect 26344 11898 26372 12174
rect 26332 11892 26384 11898
rect 26332 11834 26384 11840
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 26436 10674 26464 13738
rect 26988 13530 27016 13806
rect 26976 13524 27028 13530
rect 26976 13466 27028 13472
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26528 12850 26556 13126
rect 26620 12986 26648 13126
rect 26608 12980 26660 12986
rect 26608 12922 26660 12928
rect 26792 12980 26844 12986
rect 26792 12922 26844 12928
rect 26516 12844 26568 12850
rect 26516 12786 26568 12792
rect 26804 10674 26832 12922
rect 26988 12646 27016 13466
rect 27436 13320 27488 13326
rect 27436 13262 27488 13268
rect 27448 12986 27476 13262
rect 27436 12980 27488 12986
rect 27436 12922 27488 12928
rect 26976 12640 27028 12646
rect 26976 12582 27028 12588
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 26424 10668 26476 10674
rect 26424 10610 26476 10616
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 26436 10062 26464 10610
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26424 10056 26476 10062
rect 26424 9998 26476 10004
rect 26528 9994 26556 10406
rect 26804 10130 26832 10610
rect 26792 10124 26844 10130
rect 26792 10066 26844 10072
rect 26516 9988 26568 9994
rect 26516 9930 26568 9936
rect 26528 9654 26556 9930
rect 27344 9920 27396 9926
rect 27344 9862 27396 9868
rect 26516 9648 26568 9654
rect 26516 9590 26568 9596
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 26988 8566 27016 9522
rect 27356 9518 27384 9862
rect 27344 9512 27396 9518
rect 27344 9454 27396 9460
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26976 8560 27028 8566
rect 26976 8502 27028 8508
rect 27068 8560 27120 8566
rect 27068 8502 27120 8508
rect 26528 8090 26556 8502
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26516 7744 26568 7750
rect 26516 7686 26568 7692
rect 26528 7342 26556 7686
rect 27080 7342 27108 8502
rect 27356 8498 27384 9454
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27356 8378 27384 8434
rect 27264 8350 27384 8378
rect 27264 8294 27292 8350
rect 27252 8288 27304 8294
rect 27252 8230 27304 8236
rect 26516 7336 26568 7342
rect 26516 7278 26568 7284
rect 27068 7336 27120 7342
rect 27068 7278 27120 7284
rect 27448 5914 27476 11290
rect 27540 9518 27568 15456
rect 27804 15360 27856 15366
rect 27804 15302 27856 15308
rect 27816 13920 27844 15302
rect 27816 13892 28028 13920
rect 27804 13184 27856 13190
rect 27804 13126 27856 13132
rect 27816 12782 27844 13126
rect 27804 12776 27856 12782
rect 27804 12718 27856 12724
rect 27816 12238 27844 12718
rect 27804 12232 27856 12238
rect 27804 12174 27856 12180
rect 27712 12096 27764 12102
rect 27712 12038 27764 12044
rect 27896 12096 27948 12102
rect 27896 12038 27948 12044
rect 27724 11354 27752 12038
rect 27908 11762 27936 12038
rect 27896 11756 27948 11762
rect 27896 11698 27948 11704
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 27712 11348 27764 11354
rect 27712 11290 27764 11296
rect 27528 9512 27580 9518
rect 27528 9454 27580 9460
rect 27620 9172 27672 9178
rect 27620 9114 27672 9120
rect 27632 8634 27660 9114
rect 27712 9104 27764 9110
rect 27712 9046 27764 9052
rect 27620 8628 27672 8634
rect 27620 8570 27672 8576
rect 27724 8498 27752 9046
rect 27816 8906 27844 11494
rect 28000 11082 28028 13892
rect 28092 12850 28120 15982
rect 28172 15904 28224 15910
rect 28172 15846 28224 15852
rect 28184 15706 28212 15846
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 28172 15700 28224 15706
rect 28172 15642 28224 15648
rect 28172 15428 28224 15434
rect 28172 15370 28224 15376
rect 28080 12844 28132 12850
rect 28080 12786 28132 12792
rect 28080 12232 28132 12238
rect 28080 12174 28132 12180
rect 28092 11898 28120 12174
rect 28184 11898 28212 15370
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 28264 12368 28316 12374
rect 28264 12310 28316 12316
rect 28276 11898 28304 12310
rect 28368 12238 28396 12786
rect 28540 12640 28592 12646
rect 28540 12582 28592 12588
rect 28356 12232 28408 12238
rect 28356 12174 28408 12180
rect 28080 11892 28132 11898
rect 28080 11834 28132 11840
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 28264 11892 28316 11898
rect 28264 11834 28316 11840
rect 28080 11620 28132 11626
rect 28080 11562 28132 11568
rect 27988 11076 28040 11082
rect 27988 11018 28040 11024
rect 28000 9110 28028 11018
rect 27988 9104 28040 9110
rect 27988 9046 28040 9052
rect 27896 8968 27948 8974
rect 27896 8910 27948 8916
rect 27804 8900 27856 8906
rect 27804 8842 27856 8848
rect 27816 8498 27844 8842
rect 27908 8634 27936 8910
rect 27988 8832 28040 8838
rect 27988 8774 28040 8780
rect 27896 8628 27948 8634
rect 27896 8570 27948 8576
rect 27712 8492 27764 8498
rect 27712 8434 27764 8440
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 28000 7410 28028 8774
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 28000 6798 28028 7346
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 27436 5908 27488 5914
rect 27436 5850 27488 5856
rect 27160 5840 27212 5846
rect 27160 5782 27212 5788
rect 26424 5704 26476 5710
rect 26424 5646 26476 5652
rect 26056 5364 26108 5370
rect 26056 5306 26108 5312
rect 26436 5234 26464 5646
rect 26884 5364 26936 5370
rect 26884 5306 26936 5312
rect 25136 5228 25188 5234
rect 25136 5170 25188 5176
rect 26424 5228 26476 5234
rect 26424 5170 26476 5176
rect 23756 5160 23808 5166
rect 23756 5102 23808 5108
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 24952 5092 25004 5098
rect 24952 5034 25004 5040
rect 26240 5092 26292 5098
rect 26240 5034 26292 5040
rect 24308 5024 24360 5030
rect 24308 4966 24360 4972
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23940 4140 23992 4146
rect 23940 4082 23992 4088
rect 23480 3120 23532 3126
rect 23480 3062 23532 3068
rect 23584 3058 23612 4082
rect 23952 3738 23980 4082
rect 24320 3738 24348 4966
rect 24860 4548 24912 4554
rect 24860 4490 24912 4496
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 23940 3732 23992 3738
rect 23940 3674 23992 3680
rect 24308 3732 24360 3738
rect 24308 3674 24360 3680
rect 24400 3732 24452 3738
rect 24400 3674 24452 3680
rect 23676 3058 23704 3674
rect 24412 3534 24440 3674
rect 24400 3528 24452 3534
rect 24400 3470 24452 3476
rect 23572 3052 23624 3058
rect 23572 2994 23624 3000
rect 23664 3052 23716 3058
rect 23664 2994 23716 3000
rect 23676 2514 23704 2994
rect 24872 2774 24900 4490
rect 24780 2746 24900 2774
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 23216 2094 23336 2122
rect 23216 800 23244 2094
rect 24228 870 24348 898
rect 24228 800 24256 870
rect 18248 734 18460 762
rect 19154 0 19210 800
rect 20166 0 20222 800
rect 21178 0 21234 800
rect 22190 0 22246 800
rect 23202 0 23258 800
rect 24214 0 24270 800
rect 24320 762 24348 870
rect 24780 762 24808 2746
rect 24964 2514 24992 5034
rect 25596 4616 25648 4622
rect 25596 4558 25648 4564
rect 25228 4072 25280 4078
rect 25228 4014 25280 4020
rect 24952 2508 25004 2514
rect 24952 2450 25004 2456
rect 25240 800 25268 4014
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 25332 3194 25360 3402
rect 25608 3194 25636 4558
rect 26252 3670 26280 5034
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26700 4140 26752 4146
rect 26700 4082 26752 4088
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 26240 3664 26292 3670
rect 26240 3606 26292 3612
rect 26240 3528 26292 3534
rect 26240 3470 26292 3476
rect 25320 3188 25372 3194
rect 25320 3130 25372 3136
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25332 2310 25360 3130
rect 26252 3058 26280 3470
rect 26240 3052 26292 3058
rect 26240 2994 26292 3000
rect 26436 2774 26464 4014
rect 26528 3738 26556 4082
rect 26516 3732 26568 3738
rect 26516 3674 26568 3680
rect 26252 2746 26464 2774
rect 25320 2304 25372 2310
rect 25320 2246 25372 2252
rect 26252 800 26280 2746
rect 26712 2650 26740 4082
rect 26896 2990 26924 5306
rect 27172 5234 27200 5782
rect 27252 5568 27304 5574
rect 27252 5510 27304 5516
rect 27160 5228 27212 5234
rect 27160 5170 27212 5176
rect 27172 4826 27200 5170
rect 27264 5166 27292 5510
rect 27448 5370 27476 5850
rect 28092 5710 28120 11562
rect 28184 11082 28212 11834
rect 28552 11694 28580 12582
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 28540 11688 28592 11694
rect 28540 11630 28592 11636
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 28172 11076 28224 11082
rect 28172 11018 28224 11024
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28172 7336 28224 7342
rect 28172 7278 28224 7284
rect 28184 6866 28212 7278
rect 28264 7200 28316 7206
rect 28264 7142 28316 7148
rect 28172 6860 28224 6866
rect 28172 6802 28224 6808
rect 28276 5710 28304 7142
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 27528 5704 27580 5710
rect 27528 5646 27580 5652
rect 28080 5704 28132 5710
rect 28080 5646 28132 5652
rect 28264 5704 28316 5710
rect 28264 5646 28316 5652
rect 27436 5364 27488 5370
rect 27436 5306 27488 5312
rect 27252 5160 27304 5166
rect 27252 5102 27304 5108
rect 27160 4820 27212 4826
rect 27160 4762 27212 4768
rect 27264 4690 27292 5102
rect 27252 4684 27304 4690
rect 27252 4626 27304 4632
rect 27448 4622 27476 5306
rect 27540 5166 27568 5646
rect 27712 5568 27764 5574
rect 27712 5510 27764 5516
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 27528 5160 27580 5166
rect 27528 5102 27580 5108
rect 27724 4622 27752 5510
rect 28184 5302 28212 5510
rect 28172 5296 28224 5302
rect 28172 5238 28224 5244
rect 28460 5234 28488 6802
rect 28920 5710 28948 8774
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 28908 5704 28960 5710
rect 28908 5646 28960 5652
rect 28540 5568 28592 5574
rect 28540 5510 28592 5516
rect 27804 5228 27856 5234
rect 27804 5170 27856 5176
rect 28448 5228 28500 5234
rect 28448 5170 28500 5176
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 27712 4616 27764 4622
rect 27712 4558 27764 4564
rect 27816 4486 27844 5170
rect 28552 5166 28580 5510
rect 28920 5234 28948 5646
rect 29552 5568 29604 5574
rect 29552 5510 29604 5516
rect 29564 5302 29592 5510
rect 29552 5296 29604 5302
rect 29552 5238 29604 5244
rect 30840 5296 30892 5302
rect 30840 5238 30892 5244
rect 28908 5228 28960 5234
rect 28908 5170 28960 5176
rect 28540 5160 28592 5166
rect 28540 5102 28592 5108
rect 30104 5160 30156 5166
rect 30104 5102 30156 5108
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 29000 5024 29052 5030
rect 29000 4966 29052 4972
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27988 4480 28040 4486
rect 27988 4422 28040 4428
rect 27712 3936 27764 3942
rect 27712 3878 27764 3884
rect 26976 3460 27028 3466
rect 26976 3402 27028 3408
rect 26988 3126 27016 3402
rect 27528 3188 27580 3194
rect 27528 3130 27580 3136
rect 26976 3120 27028 3126
rect 26976 3062 27028 3068
rect 26884 2984 26936 2990
rect 26884 2926 26936 2932
rect 26976 2984 27028 2990
rect 26976 2926 27028 2932
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 26988 2514 27016 2926
rect 27436 2848 27488 2854
rect 27264 2808 27436 2836
rect 26976 2508 27028 2514
rect 26976 2450 27028 2456
rect 27264 800 27292 2808
rect 27436 2790 27488 2796
rect 27540 2514 27568 3130
rect 27724 3126 27752 3878
rect 27802 3496 27858 3505
rect 27802 3431 27858 3440
rect 27712 3120 27764 3126
rect 27712 3062 27764 3068
rect 27528 2508 27580 2514
rect 27528 2450 27580 2456
rect 27724 2378 27752 3062
rect 27816 2990 27844 3431
rect 27804 2984 27856 2990
rect 27804 2926 27856 2932
rect 28000 2774 28028 4422
rect 28816 3732 28868 3738
rect 28816 3674 28868 3680
rect 28724 3664 28776 3670
rect 28724 3606 28776 3612
rect 28736 2774 28764 3606
rect 28828 3398 28856 3674
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 28828 3058 28856 3334
rect 29012 3126 29040 4966
rect 29104 4078 29132 5034
rect 30116 4282 30144 5102
rect 29184 4276 29236 4282
rect 29184 4218 29236 4224
rect 30104 4276 30156 4282
rect 30104 4218 30156 4224
rect 29092 4072 29144 4078
rect 29092 4014 29144 4020
rect 29196 3738 29224 4218
rect 30852 4214 30880 5238
rect 31852 5024 31904 5030
rect 31852 4966 31904 4972
rect 30380 4208 30432 4214
rect 30380 4150 30432 4156
rect 30840 4208 30892 4214
rect 30840 4150 30892 4156
rect 29184 3732 29236 3738
rect 29184 3674 29236 3680
rect 29276 3664 29328 3670
rect 29276 3606 29328 3612
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 29000 3120 29052 3126
rect 29000 3062 29052 3068
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 27908 2746 28028 2774
rect 28460 2746 28764 2774
rect 27908 2514 27936 2746
rect 27896 2508 27948 2514
rect 27896 2450 27948 2456
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 28460 1714 28488 2746
rect 29104 2446 29132 3538
rect 29184 3528 29236 3534
rect 29184 3470 29236 3476
rect 29196 3194 29224 3470
rect 29184 3188 29236 3194
rect 29184 3130 29236 3136
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 28276 1686 28488 1714
rect 28276 800 28304 1686
rect 29288 800 29316 3606
rect 30392 3126 30420 4150
rect 30564 3936 30616 3942
rect 30564 3878 30616 3884
rect 30576 3194 30604 3878
rect 31864 3534 31892 4966
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 32312 3596 32364 3602
rect 32312 3538 32364 3544
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31852 3528 31904 3534
rect 31852 3470 31904 3476
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30380 3120 30432 3126
rect 30380 3062 30432 3068
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30392 2378 30420 2790
rect 31036 2650 31064 3470
rect 31300 2984 31352 2990
rect 31300 2926 31352 2932
rect 31024 2644 31076 2650
rect 31024 2586 31076 2592
rect 30472 2508 30524 2514
rect 30472 2450 30524 2456
rect 30380 2372 30432 2378
rect 30380 2314 30432 2320
rect 30484 1442 30512 2450
rect 30300 1414 30512 1442
rect 30300 800 30328 1414
rect 31312 800 31340 2926
rect 32128 2848 32180 2854
rect 32128 2790 32180 2796
rect 32140 2446 32168 2790
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32324 800 32352 3538
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 33612 3194 33640 3334
rect 33600 3188 33652 3194
rect 33600 3130 33652 3136
rect 33324 3052 33376 3058
rect 33324 2994 33376 3000
rect 33336 800 33364 2994
rect 34244 2848 34296 2854
rect 34244 2790 34296 2796
rect 34256 2514 34284 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34244 2508 34296 2514
rect 34244 2450 34296 2456
rect 34520 2440 34572 2446
rect 34520 2382 34572 2388
rect 35348 2440 35400 2446
rect 35348 2382 35400 2388
rect 34532 1442 34560 2382
rect 34348 1414 34560 1442
rect 34348 800 34376 1414
rect 35360 800 35388 2382
rect 24320 734 24808 762
rect 25226 0 25282 800
rect 26238 0 26294 800
rect 27250 0 27306 800
rect 28262 0 28318 800
rect 29274 0 29330 800
rect 30286 0 30342 800
rect 31298 0 31354 800
rect 32310 0 32366 800
rect 33322 0 33378 800
rect 34334 0 34390 800
rect 35346 0 35402 800
<< via2 >>
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10230 11500 10232 11520
rect 10232 11500 10284 11520
rect 10284 11500 10286 11520
rect 10230 11464 10286 11500
rect 12714 11464 12770 11520
rect 14370 11056 14426 11112
rect 14370 10920 14426 10976
rect 14370 7792 14426 7848
rect 15014 12708 15070 12744
rect 15014 12688 15016 12708
rect 15016 12688 15068 12708
rect 15068 12688 15070 12708
rect 15934 12688 15990 12744
rect 15842 10920 15898 10976
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19890 3476 19892 3496
rect 19892 3476 19944 3496
rect 19944 3476 19946 3496
rect 19890 3440 19946 3476
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 27802 3440 27858 3496
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
<< metal3 >>
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 15009 12746 15075 12749
rect 15929 12746 15995 12749
rect 15009 12744 15995 12746
rect 15009 12688 15014 12744
rect 15070 12688 15934 12744
rect 15990 12688 15995 12744
rect 15009 12686 15995 12688
rect 15009 12683 15075 12686
rect 15929 12683 15995 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 10225 11522 10291 11525
rect 12709 11522 12775 11525
rect 10225 11520 12775 11522
rect 10225 11464 10230 11520
rect 10286 11464 12714 11520
rect 12770 11464 12775 11520
rect 10225 11462 12775 11464
rect 10225 11459 10291 11462
rect 12709 11459 12775 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 14365 11116 14431 11117
rect 14365 11114 14412 11116
rect 14320 11112 14412 11114
rect 14320 11056 14370 11112
rect 14320 11054 14412 11056
rect 14365 11052 14412 11054
rect 14476 11052 14482 11116
rect 14365 11051 14431 11052
rect 14365 10978 14431 10981
rect 15837 10978 15903 10981
rect 14365 10976 15903 10978
rect 14365 10920 14370 10976
rect 14426 10920 15842 10976
rect 15898 10920 15903 10976
rect 14365 10918 15903 10920
rect 14365 10915 14431 10918
rect 15837 10915 15903 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 14365 7852 14431 7853
rect 14365 7848 14412 7852
rect 14476 7850 14482 7852
rect 14365 7792 14370 7848
rect 14365 7788 14412 7792
rect 14476 7790 14522 7850
rect 14476 7788 14482 7790
rect 14365 7787 14431 7788
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19885 3498 19951 3501
rect 27797 3498 27863 3501
rect 19885 3496 27863 3498
rect 19885 3440 19890 3496
rect 19946 3440 27802 3496
rect 27858 3440 27863 3496
rect 19885 3438 27863 3440
rect 19885 3435 19951 3438
rect 27797 3435 27863 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 14412 11112 14476 11116
rect 14412 11056 14426 11112
rect 14426 11056 14476 11112
rect 14412 11052 14476 11056
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 14412 7848 14476 7852
rect 14412 7792 14426 7848
rect 14426 7792 14476 7848
rect 14412 7788 14476 7792
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 36480 4528 36496
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 19568 35936 19888 36496
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 14411 11116 14477 11117
rect 14411 11052 14412 11116
rect 14476 11052 14477 11116
rect 14411 11051 14477 11052
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 14414 7853 14474 11051
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 14411 7852 14477 7853
rect 14411 7788 14412 7852
rect 14476 7788 14477 7852
rect 14411 7787 14477 7788
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 36480 35248 36496
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _380_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _381_
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _382_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _383_
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _384_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _385_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _386_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _387_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_4  _388_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _389_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _390_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _391_
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__o22a_1  _392_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15456 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _393_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _394_
timestamp 1688980957
transform 1 0 13248 0 -1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _395_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15824 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_4  _396_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_4  _397_
timestamp 1688980957
transform 1 0 8280 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _398_
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _399_
timestamp 1688980957
transform 1 0 14260 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _400_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _401_
timestamp 1688980957
transform 1 0 11592 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _402_
timestamp 1688980957
transform 1 0 11592 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _403_
timestamp 1688980957
transform 1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _404_
timestamp 1688980957
transform -1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _405_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15456 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _406_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _407_
timestamp 1688980957
transform 1 0 15272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _408_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17204 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_4  _409_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_4  _410_
timestamp 1688980957
transform 1 0 6808 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _411_
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_2  _412_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16744 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _413_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_2  _414_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _415_
timestamp 1688980957
transform 1 0 9936 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _416_
timestamp 1688980957
transform 1 0 9936 0 1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_2  _417_
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _418_
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _419_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _420_
timestamp 1688980957
transform 1 0 15824 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _421_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _422_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16100 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _423_
timestamp 1688980957
transform -1 0 16652 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _424_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _425_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _426_
timestamp 1688980957
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _427_
timestamp 1688980957
transform -1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _428_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _429_
timestamp 1688980957
transform -1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _430_
timestamp 1688980957
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _431_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _432_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _433_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12144 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _434_
timestamp 1688980957
transform 1 0 11960 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1688980957
transform -1 0 23920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _436_
timestamp 1688980957
transform -1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _437_
timestamp 1688980957
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _438_
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _439_
timestamp 1688980957
transform 1 0 9936 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _440_
timestamp 1688980957
transform 1 0 13248 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _441_
timestamp 1688980957
transform 1 0 17940 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _443_
timestamp 1688980957
transform 1 0 19228 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _444_
timestamp 1688980957
transform 1 0 18032 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _445_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_2  _446_
timestamp 1688980957
transform -1 0 15456 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _447_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _448_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_1  _449_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16560 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _450_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _451_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _452_
timestamp 1688980957
transform 1 0 19412 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _453_
timestamp 1688980957
transform -1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _454_
timestamp 1688980957
transform -1 0 20424 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _455_
timestamp 1688980957
transform -1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _456_
timestamp 1688980957
transform -1 0 20424 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _457_
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _458_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20332 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _460_
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _461_
timestamp 1688980957
transform 1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _462_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17020 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _463_
timestamp 1688980957
transform -1 0 16652 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _464_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _465_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _466_
timestamp 1688980957
transform -1 0 18400 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _467_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _468_
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _469_
timestamp 1688980957
transform -1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _470_
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _471_
timestamp 1688980957
transform -1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _472_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12880 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _473_
timestamp 1688980957
transform 1 0 12144 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _474_
timestamp 1688980957
transform 1 0 12788 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_1  _475_
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _476_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _477_
timestamp 1688980957
transform 1 0 17204 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _478_
timestamp 1688980957
transform -1 0 11316 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _479_
timestamp 1688980957
transform -1 0 10672 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _480_
timestamp 1688980957
transform -1 0 11408 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_1  _481_
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _482_
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _483_
timestamp 1688980957
transform 1 0 12052 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _484_
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _485_
timestamp 1688980957
transform -1 0 18584 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _486_
timestamp 1688980957
transform 1 0 18952 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _487_
timestamp 1688980957
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _488_
timestamp 1688980957
transform -1 0 20240 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _489_
timestamp 1688980957
transform 1 0 20240 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _490_
timestamp 1688980957
transform -1 0 21528 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _491_
timestamp 1688980957
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _492_
timestamp 1688980957
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _493_
timestamp 1688980957
transform 1 0 20424 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _494_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21528 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _495_
timestamp 1688980957
transform -1 0 20608 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _496_
timestamp 1688980957
transform 1 0 21620 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _497_
timestamp 1688980957
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _498_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18032 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _499_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _500_
timestamp 1688980957
transform -1 0 20608 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _501_
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _502_
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _503_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13340 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _504_
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_2  _505_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16100 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _506_
timestamp 1688980957
transform -1 0 18492 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _507_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16468 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _508_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a2111o_1  _509_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _510_
timestamp 1688980957
transform 1 0 16744 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _511_
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _512_
timestamp 1688980957
transform -1 0 10120 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _513_
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _514_
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _515_
timestamp 1688980957
transform 1 0 10856 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _516_
timestamp 1688980957
transform -1 0 12236 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _517_
timestamp 1688980957
transform 1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _518_
timestamp 1688980957
transform -1 0 12144 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _519_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _520_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _521_
timestamp 1688980957
transform 1 0 18768 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _522_
timestamp 1688980957
transform 1 0 19412 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _523_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _524_
timestamp 1688980957
transform 1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _525_
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1688980957
transform 1 0 21804 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _527_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _528_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23000 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _529_
timestamp 1688980957
transform 1 0 21068 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _530_
timestamp 1688980957
transform 1 0 20148 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _531_
timestamp 1688980957
transform -1 0 19780 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _532_
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_4  _533_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  _534_
timestamp 1688980957
transform 1 0 20700 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_4  _535_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__a2bb2o_1  _536_
timestamp 1688980957
transform -1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _537_
timestamp 1688980957
transform -1 0 15640 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _538_
timestamp 1688980957
transform -1 0 14536 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _539_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14536 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _540_
timestamp 1688980957
transform 1 0 14720 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _541_
timestamp 1688980957
transform 1 0 15364 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _542_
timestamp 1688980957
transform -1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _543_
timestamp 1688980957
transform -1 0 16468 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _544_
timestamp 1688980957
transform -1 0 16744 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _545_
timestamp 1688980957
transform 1 0 15732 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _546_
timestamp 1688980957
transform 1 0 16652 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_4  _547_
timestamp 1688980957
transform -1 0 10948 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _548_
timestamp 1688980957
transform 1 0 9384 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _549_
timestamp 1688980957
transform 1 0 10764 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_4  _550_
timestamp 1688980957
transform -1 0 12880 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__or4b_4  _551_
timestamp 1688980957
transform -1 0 10212 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__a2bb2o_1  _552_
timestamp 1688980957
transform 1 0 9108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _553_
timestamp 1688980957
transform 1 0 9108 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _554_
timestamp 1688980957
transform 1 0 9752 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _555_
timestamp 1688980957
transform 1 0 9108 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _556_
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _557_
timestamp 1688980957
transform -1 0 10304 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _558_
timestamp 1688980957
transform -1 0 11408 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _559_
timestamp 1688980957
transform -1 0 11132 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _560_
timestamp 1688980957
transform -1 0 11500 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _561_
timestamp 1688980957
transform 1 0 10948 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _562_
timestamp 1688980957
transform 1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _563_
timestamp 1688980957
transform -1 0 21252 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _564_
timestamp 1688980957
transform -1 0 20056 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _565_
timestamp 1688980957
transform 1 0 19412 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _566_
timestamp 1688980957
transform -1 0 20240 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _567_
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _568_
timestamp 1688980957
transform 1 0 20240 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _569_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22356 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _570_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _571_
timestamp 1688980957
transform -1 0 22356 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _572_
timestamp 1688980957
transform -1 0 23552 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _573_
timestamp 1688980957
transform 1 0 22172 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _574_
timestamp 1688980957
transform -1 0 21712 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _575_
timestamp 1688980957
transform 1 0 20056 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _576_
timestamp 1688980957
transform -1 0 18308 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _577_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _578_
timestamp 1688980957
transform -1 0 15640 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _579_
timestamp 1688980957
transform 1 0 14536 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _580_
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _581_
timestamp 1688980957
transform -1 0 15548 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _582_
timestamp 1688980957
transform 1 0 14444 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _583_
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _584_
timestamp 1688980957
transform 1 0 18032 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _585_
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _586_
timestamp 1688980957
transform -1 0 13616 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _587_
timestamp 1688980957
transform -1 0 9016 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _588_
timestamp 1688980957
transform 1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _589_
timestamp 1688980957
transform 1 0 9016 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_2  _590_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9476 0 -1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _591_
timestamp 1688980957
transform 1 0 10580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _592_
timestamp 1688980957
transform -1 0 9752 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _593_
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _594_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _595_
timestamp 1688980957
transform 1 0 12696 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _596_
timestamp 1688980957
transform 1 0 12144 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _597_
timestamp 1688980957
transform 1 0 20976 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _598_
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _599_
timestamp 1688980957
transform 1 0 19780 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _600_
timestamp 1688980957
transform 1 0 20516 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__a311o_1  _601_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _602_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _603_
timestamp 1688980957
transform 1 0 23736 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _604_
timestamp 1688980957
transform 1 0 22448 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _605_
timestamp 1688980957
transform 1 0 23000 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _606_
timestamp 1688980957
transform -1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _607_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _608_
timestamp 1688980957
transform -1 0 21712 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _609_
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _610_
timestamp 1688980957
transform 1 0 20424 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _611_
timestamp 1688980957
transform -1 0 18032 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _612_
timestamp 1688980957
transform -1 0 15916 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _613_
timestamp 1688980957
transform 1 0 16744 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _614_
timestamp 1688980957
transform -1 0 16192 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _615_
timestamp 1688980957
transform 1 0 15088 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _616_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15088 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _617_
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _618_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _619_
timestamp 1688980957
transform -1 0 17020 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _620_
timestamp 1688980957
transform 1 0 17204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _621_
timestamp 1688980957
transform -1 0 17572 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _622_
timestamp 1688980957
transform 1 0 18492 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _623_
timestamp 1688980957
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _624_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_2  _625_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__xnor2_1  _626_
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _627_
timestamp 1688980957
transform -1 0 10212 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _628_
timestamp 1688980957
transform -1 0 9936 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _629_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11592 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _630_
timestamp 1688980957
transform -1 0 10856 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _631_
timestamp 1688980957
transform 1 0 12236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _632_
timestamp 1688980957
transform -1 0 12604 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _633_
timestamp 1688980957
transform 1 0 12972 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _634_
timestamp 1688980957
transform -1 0 13984 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _635_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_1  _636_
timestamp 1688980957
transform -1 0 19136 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _637_
timestamp 1688980957
transform -1 0 21528 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _638_
timestamp 1688980957
transform 1 0 20608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _639_
timestamp 1688980957
transform -1 0 21620 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _640_
timestamp 1688980957
transform 1 0 21160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _641_
timestamp 1688980957
transform 1 0 21896 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _642_
timestamp 1688980957
transform -1 0 21896 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _643_
timestamp 1688980957
transform 1 0 21896 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _644_
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ba_1  _645_
timestamp 1688980957
transform -1 0 25208 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _646_
timestamp 1688980957
transform 1 0 21896 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _647_
timestamp 1688980957
transform -1 0 16468 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _648_
timestamp 1688980957
transform -1 0 16376 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _649_
timestamp 1688980957
transform 1 0 16652 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _650_
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _651_
timestamp 1688980957
transform 1 0 18216 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _652_
timestamp 1688980957
transform 1 0 10212 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _653_
timestamp 1688980957
transform -1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _654_
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_1  _655_
timestamp 1688980957
transform 1 0 12696 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _656_
timestamp 1688980957
transform -1 0 13800 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _657_
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _658_
timestamp 1688980957
transform -1 0 21528 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _659_
timestamp 1688980957
transform 1 0 20884 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a21boi_2  _660_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _661_
timestamp 1688980957
transform 1 0 21988 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _662_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23736 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _663_
timestamp 1688980957
transform 1 0 23092 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _664_
timestamp 1688980957
transform -1 0 23552 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _665_
timestamp 1688980957
transform -1 0 24380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _666_
timestamp 1688980957
transform -1 0 23276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _667_
timestamp 1688980957
transform 1 0 22724 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _668_
timestamp 1688980957
transform 1 0 24380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _669_
timestamp 1688980957
transform -1 0 24104 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _670_
timestamp 1688980957
transform -1 0 24932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _671_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _672_
timestamp 1688980957
transform -1 0 25300 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _673_
timestamp 1688980957
transform -1 0 24840 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _674_
timestamp 1688980957
transform 1 0 24840 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _675_
timestamp 1688980957
transform 1 0 24932 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_2  _676_
timestamp 1688980957
transform -1 0 26496 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _677_
timestamp 1688980957
transform -1 0 24932 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _678_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_2  _679_
timestamp 1688980957
transform 1 0 17388 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _680_
timestamp 1688980957
transform -1 0 12696 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _681_
timestamp 1688980957
transform -1 0 13432 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _682_
timestamp 1688980957
transform -1 0 25208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _683_
timestamp 1688980957
transform 1 0 24564 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_2  _684_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22724 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _685_
timestamp 1688980957
transform 1 0 26036 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _686_
timestamp 1688980957
transform 1 0 25392 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _687_
timestamp 1688980957
transform 1 0 28152 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _688_
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_1  _689_
timestamp 1688980957
transform 1 0 23368 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _690_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23736 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _691_
timestamp 1688980957
transform 1 0 24380 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _692_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _693_
timestamp 1688980957
transform -1 0 24104 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _694_
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _695_
timestamp 1688980957
transform -1 0 25668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _696_
timestamp 1688980957
transform -1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _697_
timestamp 1688980957
transform 1 0 26128 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _698_
timestamp 1688980957
transform 1 0 26128 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _699_
timestamp 1688980957
transform 1 0 26036 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _700_
timestamp 1688980957
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _701_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _702_
timestamp 1688980957
transform 1 0 27416 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _703_
timestamp 1688980957
transform -1 0 29164 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _704_
timestamp 1688980957
transform -1 0 28704 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _705_
timestamp 1688980957
transform 1 0 27692 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _706_
timestamp 1688980957
transform -1 0 28888 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _707_
timestamp 1688980957
transform -1 0 26772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _708_
timestamp 1688980957
transform 1 0 23828 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _709_
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _710_
timestamp 1688980957
transform 1 0 23460 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _711_
timestamp 1688980957
transform 1 0 24932 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _712_
timestamp 1688980957
transform -1 0 25852 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _713_
timestamp 1688980957
transform 1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _714_
timestamp 1688980957
transform -1 0 26128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _715_
timestamp 1688980957
transform -1 0 26036 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _716_
timestamp 1688980957
transform 1 0 25484 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _717_
timestamp 1688980957
transform 1 0 26496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _718_
timestamp 1688980957
transform 1 0 26772 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _719_
timestamp 1688980957
transform 1 0 27232 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _720_
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _721_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26864 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _722_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 27968 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _723_
timestamp 1688980957
transform 1 0 27968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _724_
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _725_
timestamp 1688980957
transform -1 0 27968 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _726_
timestamp 1688980957
transform -1 0 28244 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _727_
timestamp 1688980957
transform -1 0 25576 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _728_
timestamp 1688980957
transform -1 0 24012 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _729_
timestamp 1688980957
transform 1 0 23184 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _730_
timestamp 1688980957
transform -1 0 25116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _731_
timestamp 1688980957
transform 1 0 24564 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _732_
timestamp 1688980957
transform 1 0 24932 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _733_
timestamp 1688980957
transform -1 0 25484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _734_
timestamp 1688980957
transform 1 0 25208 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _735_
timestamp 1688980957
transform 1 0 25760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _736_
timestamp 1688980957
transform -1 0 25484 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _737_
timestamp 1688980957
transform 1 0 25668 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _738_
timestamp 1688980957
transform -1 0 26496 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _739_
timestamp 1688980957
transform 1 0 26496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _740_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _741_
timestamp 1688980957
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _742_
timestamp 1688980957
transform -1 0 27692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _743_
timestamp 1688980957
transform 1 0 27600 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _744_
timestamp 1688980957
transform 1 0 27692 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _745_
timestamp 1688980957
transform 1 0 27140 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _746_
timestamp 1688980957
transform 1 0 27784 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _747_
timestamp 1688980957
transform -1 0 25300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _748_
timestamp 1688980957
transform -1 0 24380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _749_
timestamp 1688980957
transform 1 0 24840 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _750_
timestamp 1688980957
transform -1 0 27508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _751_
timestamp 1688980957
transform -1 0 26864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _752_
timestamp 1688980957
transform 1 0 28336 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _753_
timestamp 1688980957
transform -1 0 25208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _754_
timestamp 1688980957
transform -1 0 28336 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _755_
timestamp 1688980957
transform -1 0 28796 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _756_
timestamp 1688980957
transform 1 0 27876 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _757_
timestamp 1688980957
transform -1 0 28980 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _758_
timestamp 1688980957
transform -1 0 29624 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _759_
timestamp 1688980957
transform 1 0 27140 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _760_
timestamp 1688980957
transform 1 0 27048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _761_
timestamp 1688980957
transform 1 0 27600 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _762_
timestamp 1688980957
transform -1 0 27600 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _763_
timestamp 1688980957
transform 1 0 25208 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _764_
timestamp 1688980957
transform 1 0 24104 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _765_
timestamp 1688980957
transform 1 0 23368 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _766_
timestamp 1688980957
transform 1 0 22356 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _767_
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _768_
timestamp 1688980957
transform 1 0 20608 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _769_
timestamp 1688980957
transform 1 0 19320 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _770_
timestamp 1688980957
transform 1 0 17572 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _771_
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _772_
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _773_
timestamp 1688980957
transform -1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _774_
timestamp 1688980957
transform -1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _775_
timestamp 1688980957
transform 1 0 15180 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dfrtp_1  _776_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _777_
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _778_
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp 1688980957
transform 1 0 17940 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _780_
timestamp 1688980957
transform 1 0 19780 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _781_
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _782_
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _783_
timestamp 1688980957
transform 1 0 23644 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _784_
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _785_
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _786_
timestamp 1688980957
transform 1 0 26220 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _787_
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _788_
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _789_
timestamp 1688980957
transform 1 0 28796 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _790_
timestamp 1688980957
transform 1 0 28796 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _791_
timestamp 1688980957
transform 1 0 30084 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _792_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _793_
timestamp 1688980957
transform 1 0 4140 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _794_
timestamp 1688980957
transform 1 0 5152 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _795_
timestamp 1688980957
transform 1 0 6716 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _796_
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _797_
timestamp 1688980957
transform -1 0 11132 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _798_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8464 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _799_
timestamp 1688980957
transform -1 0 12972 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _800_
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _801_
timestamp 1688980957
transform 1 0 5152 0 1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _802_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _803_
timestamp 1688980957
transform 1 0 6900 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _804_
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _805_
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _806_
timestamp 1688980957
transform -1 0 13984 0 1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _807_
timestamp 1688980957
transform -1 0 15640 0 -1 3264
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _808_
timestamp 1688980957
transform -1 0 14076 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__515__B pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__C
timestamp 1688980957
transform 1 0 10304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__551__D_N
timestamp 1688980957
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__A2_N
timestamp 1688980957
transform 1 0 9200 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__552__B1
timestamp 1688980957
transform 1 0 11592 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__B
timestamp 1688980957
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__A2
timestamp 1688980957
transform -1 0 9292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__588__B1
timestamp 1688980957
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__590__A3
timestamp 1688980957
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A2_N
timestamp 1688980957
transform 1 0 12144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__B1
timestamp 1688980957
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__625__A2
timestamp 1688980957
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__A2
timestamp 1688980957
transform -1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__653__B1
timestamp 1688980957
transform 1 0 11316 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__665__B
timestamp 1688980957
transform 1 0 23920 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__680__C1
timestamp 1688980957
transform -1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__692__C
timestamp 1688980957
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__692__D_N
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__A2_N
timestamp 1688980957
transform 1 0 23184 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__693__B1
timestamp 1688980957
transform 1 0 23000 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__708__B
timestamp 1688980957
transform 1 0 23644 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__710__C_N
timestamp 1688980957
transform 1 0 23276 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__727__B
timestamp 1688980957
transform -1 0 25668 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__728__B
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__729__A1
timestamp 1688980957
transform 1 0 23000 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__748__A2
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__748__C1
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__753__B1
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__808__D
timestamp 1688980957
transform -1 0 14444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__buf_6  fanout36 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20056 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  fanout37 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout38
timestamp 1688980957
transform -1 0 18676 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout39 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28704 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_13 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_24
timestamp 1688980957
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_35
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_46
timestamp 1688980957
transform 1 0 5336 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_60
timestamp 1688980957
transform 1 0 6624 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_64 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6992 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_68
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_79
timestamp 1688980957
transform 1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_90
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_136
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_172
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_213
timestamp 1688980957
transform 1 0 20700 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_241
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_276
timestamp 1688980957
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_281 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_325
timestamp 1688980957
transform 1 0 31004 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_353
timestamp 1688980957
transform 1 0 33580 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_109
timestamp 1688980957
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_119
timestamp 1688980957
transform 1 0 12052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_134
timestamp 1688980957
transform 1 0 13432 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_158
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_265
timestamp 1688980957
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 1688980957
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_327
timestamp 1688980957
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_356
timestamp 1688980957
transform 1 0 33856 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_37
timestamp 1688980957
transform 1 0 4508 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_93
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_191
timestamp 1688980957
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_206
timestamp 1688980957
transform 1 0 20056 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_212
timestamp 1688980957
transform 1 0 20608 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_293
timestamp 1688980957
transform 1 0 28060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_299
timestamp 1688980957
transform 1 0 28612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_304
timestamp 1688980957
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_109
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_117
timestamp 1688980957
transform 1 0 11868 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_145
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_163
timestamp 1688980957
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_202
timestamp 1688980957
transform 1 0 19688 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_214
timestamp 1688980957
transform 1 0 20792 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_222
timestamp 1688980957
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_229
timestamp 1688980957
transform 1 0 22172 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_262
timestamp 1688980957
transform 1 0 25208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_297
timestamp 1688980957
transform 1 0 28428 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_321
timestamp 1688980957
transform 1 0 30636 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_333
timestamp 1688980957
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_367
timestamp 1688980957
transform 1 0 34868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_67
timestamp 1688980957
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1688980957
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_129
timestamp 1688980957
transform 1 0 12972 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_163
timestamp 1688980957
transform 1 0 16100 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_172
timestamp 1688980957
transform 1 0 16928 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_178
timestamp 1688980957
transform 1 0 17480 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_219
timestamp 1688980957
transform 1 0 21252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_225
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_269
timestamp 1688980957
transform 1 0 25852 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_281
timestamp 1688980957
transform 1 0 26956 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_293
timestamp 1688980957
transform 1 0 28060 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_305
timestamp 1688980957
transform 1 0 29164 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_120
timestamp 1688980957
transform 1 0 12144 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_128
timestamp 1688980957
transform 1 0 12880 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_163
timestamp 1688980957
transform 1 0 16100 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_175
timestamp 1688980957
transform 1 0 17204 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_187
timestamp 1688980957
transform 1 0 18308 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_199
timestamp 1688980957
transform 1 0 19412 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_208
timestamp 1688980957
transform 1 0 20240 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_216
timestamp 1688980957
transform 1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_229
timestamp 1688980957
transform 1 0 22172 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_238
timestamp 1688980957
transform 1 0 23000 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_257
timestamp 1688980957
transform 1 0 24748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_276
timestamp 1688980957
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_295
timestamp 1688980957
transform 1 0 28244 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_310
timestamp 1688980957
transform 1 0 29624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_314
timestamp 1688980957
transform 1 0 29992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_367
timestamp 1688980957
transform 1 0 34868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_67
timestamp 1688980957
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_79
timestamp 1688980957
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_94
timestamp 1688980957
transform 1 0 9752 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_111
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_147
timestamp 1688980957
transform 1 0 14628 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_151
timestamp 1688980957
transform 1 0 14996 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_156
timestamp 1688980957
transform 1 0 15456 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_168
timestamp 1688980957
transform 1 0 16560 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_179
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_188
timestamp 1688980957
transform 1 0 18400 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_201
timestamp 1688980957
transform 1 0 19596 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_217
timestamp 1688980957
transform 1 0 21068 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_229
timestamp 1688980957
transform 1 0 22172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_248
timestamp 1688980957
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_262
timestamp 1688980957
transform 1 0 25208 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_274
timestamp 1688980957
transform 1 0 26312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_279
timestamp 1688980957
transform 1 0 26772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_286
timestamp 1688980957
transform 1 0 27416 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_141
timestamp 1688980957
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_145
timestamp 1688980957
transform 1 0 14444 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_153
timestamp 1688980957
transform 1 0 15180 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_157
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_189
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_197
timestamp 1688980957
transform 1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_202
timestamp 1688980957
transform 1 0 19688 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_214
timestamp 1688980957
transform 1 0 20792 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_222
timestamp 1688980957
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_367
timestamp 1688980957
transform 1 0 34868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_169
timestamp 1688980957
transform 1 0 16652 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_182
timestamp 1688980957
transform 1 0 17848 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_204
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_210
timestamp 1688980957
transform 1 0 20424 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_216
timestamp 1688980957
transform 1 0 20976 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_241
timestamp 1688980957
transform 1 0 23276 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_298
timestamp 1688980957
transform 1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_306
timestamp 1688980957
transform 1 0 29256 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_95
timestamp 1688980957
transform 1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_146
timestamp 1688980957
transform 1 0 14536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_155
timestamp 1688980957
transform 1 0 15364 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_182
timestamp 1688980957
transform 1 0 17848 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_190
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_202
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_211
timestamp 1688980957
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_222
timestamp 1688980957
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_233
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_240
timestamp 1688980957
transform 1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_244
timestamp 1688980957
transform 1 0 23552 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_253
timestamp 1688980957
transform 1 0 24380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_257
timestamp 1688980957
transform 1 0 24748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_265
timestamp 1688980957
transform 1 0 25484 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_287
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_299
timestamp 1688980957
transform 1 0 28612 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_311
timestamp 1688980957
transform 1 0 29716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_323
timestamp 1688980957
transform 1 0 30820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_367
timestamp 1688980957
transform 1 0 34868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_99
timestamp 1688980957
transform 1 0 10212 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_105
timestamp 1688980957
transform 1 0 10764 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_117
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_138
timestamp 1688980957
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_149
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_157
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_169
timestamp 1688980957
transform 1 0 16652 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_181
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_226
timestamp 1688980957
transform 1 0 21896 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_249
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_266
timestamp 1688980957
transform 1 0 25576 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_279
timestamp 1688980957
transform 1 0 26772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_291
timestamp 1688980957
transform 1 0 27876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_303
timestamp 1688980957
transform 1 0 28980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_100
timestamp 1688980957
transform 1 0 10304 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_121
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_156
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_182
timestamp 1688980957
transform 1 0 17848 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_199
timestamp 1688980957
transform 1 0 19412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_212
timestamp 1688980957
transform 1 0 20608 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_252
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_256
timestamp 1688980957
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_263
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_267
timestamp 1688980957
transform 1 0 25668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_275
timestamp 1688980957
transform 1 0 26404 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_294
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_306
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_318
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_330
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_367
timestamp 1688980957
transform 1 0 34868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_118
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_130
timestamp 1688980957
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_181
timestamp 1688980957
transform 1 0 17756 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_193
timestamp 1688980957
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_213
timestamp 1688980957
transform 1 0 20700 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_224
timestamp 1688980957
transform 1 0 21712 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_230
timestamp 1688980957
transform 1 0 22264 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_238
timestamp 1688980957
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_242
timestamp 1688980957
transform 1 0 23368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_248
timestamp 1688980957
transform 1 0 23920 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_260
timestamp 1688980957
transform 1 0 25024 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_303
timestamp 1688980957
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_77
timestamp 1688980957
transform 1 0 8188 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_100
timestamp 1688980957
transform 1 0 10304 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_136
timestamp 1688980957
transform 1 0 13616 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_148
timestamp 1688980957
transform 1 0 14720 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_160
timestamp 1688980957
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_187
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_199
timestamp 1688980957
transform 1 0 19412 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_212
timestamp 1688980957
transform 1 0 20608 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_231
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_240
timestamp 1688980957
transform 1 0 23184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_272
timestamp 1688980957
transform 1 0 26128 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_288
timestamp 1688980957
transform 1 0 27600 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_300
timestamp 1688980957
transform 1 0 28704 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_312
timestamp 1688980957
transform 1 0 29808 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_324
timestamp 1688980957
transform 1 0 30912 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_367
timestamp 1688980957
transform 1 0 34868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_61
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_107
timestamp 1688980957
transform 1 0 10948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_113
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_127
timestamp 1688980957
transform 1 0 12788 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_148
timestamp 1688980957
transform 1 0 14720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_156
timestamp 1688980957
transform 1 0 15456 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_168
timestamp 1688980957
transform 1 0 16560 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_176
timestamp 1688980957
transform 1 0 17296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_215
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_237
timestamp 1688980957
transform 1 0 22908 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_241
timestamp 1688980957
transform 1 0 23276 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_248
timestamp 1688980957
transform 1 0 23920 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_258
timestamp 1688980957
transform 1 0 24840 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_262
timestamp 1688980957
transform 1 0 25208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_274
timestamp 1688980957
transform 1 0 26312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_278
timestamp 1688980957
transform 1 0 26680 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_287
timestamp 1688980957
transform 1 0 27508 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_299
timestamp 1688980957
transform 1 0 28612 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_87
timestamp 1688980957
transform 1 0 9108 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_119
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_156
timestamp 1688980957
transform 1 0 15456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_180
timestamp 1688980957
transform 1 0 17664 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_192
timestamp 1688980957
transform 1 0 18768 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_204
timestamp 1688980957
transform 1 0 19872 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_216
timestamp 1688980957
transform 1 0 20976 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_233
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_246
timestamp 1688980957
transform 1 0 23736 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_252
timestamp 1688980957
transform 1 0 24288 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_258
timestamp 1688980957
transform 1 0 24840 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_270
timestamp 1688980957
transform 1 0 25944 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_367
timestamp 1688980957
transform 1 0 34868 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_95
timestamp 1688980957
transform 1 0 9844 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_112
timestamp 1688980957
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_116
timestamp 1688980957
transform 1 0 11776 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_127
timestamp 1688980957
transform 1 0 12788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_170
timestamp 1688980957
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_182
timestamp 1688980957
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_203
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_215
timestamp 1688980957
transform 1 0 20884 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_227
timestamp 1688980957
transform 1 0 21988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_239
timestamp 1688980957
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_257
timestamp 1688980957
transform 1 0 24748 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_267
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_279
timestamp 1688980957
transform 1 0 26772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 1688980957
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_104
timestamp 1688980957
transform 1 0 10672 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_108
timestamp 1688980957
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_124
timestamp 1688980957
transform 1 0 12512 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_136
timestamp 1688980957
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_146
timestamp 1688980957
transform 1 0 14536 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_150
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_154
timestamp 1688980957
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_172
timestamp 1688980957
transform 1 0 16928 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_184
timestamp 1688980957
transform 1 0 18032 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_190
timestamp 1688980957
transform 1 0 18584 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_196
timestamp 1688980957
transform 1 0 19136 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_200
timestamp 1688980957
transform 1 0 19504 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_215
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_243
timestamp 1688980957
transform 1 0 23460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_251
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_277
timestamp 1688980957
transform 1 0 26588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_287
timestamp 1688980957
transform 1 0 27508 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_302
timestamp 1688980957
transform 1 0 28888 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_314
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_326
timestamp 1688980957
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_334
timestamp 1688980957
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_367
timestamp 1688980957
transform 1 0 34868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_99
timestamp 1688980957
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_103
timestamp 1688980957
transform 1 0 10580 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_120
timestamp 1688980957
transform 1 0 12144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_152
timestamp 1688980957
transform 1 0 15088 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_180
timestamp 1688980957
transform 1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_201
timestamp 1688980957
transform 1 0 19596 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_213
timestamp 1688980957
transform 1 0 20700 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_225
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_232
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_249
timestamp 1688980957
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_263
timestamp 1688980957
transform 1 0 25300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_269
timestamp 1688980957
transform 1 0 25852 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_104
timestamp 1688980957
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_140
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_146
timestamp 1688980957
transform 1 0 14536 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_163
timestamp 1688980957
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_178
timestamp 1688980957
transform 1 0 17480 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_190
timestamp 1688980957
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_197
timestamp 1688980957
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_232
timestamp 1688980957
transform 1 0 22448 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_244
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_256
timestamp 1688980957
transform 1 0 24656 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_268
timestamp 1688980957
transform 1 0 25760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_296
timestamp 1688980957
transform 1 0 28336 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_308
timestamp 1688980957
transform 1 0 29440 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_320
timestamp 1688980957
transform 1 0 30544 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_332
timestamp 1688980957
transform 1 0 31648 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_367
timestamp 1688980957
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_98
timestamp 1688980957
transform 1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_102
timestamp 1688980957
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_106
timestamp 1688980957
transform 1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_118
timestamp 1688980957
transform 1 0 11960 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_130
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_158
timestamp 1688980957
transform 1 0 15640 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_164
timestamp 1688980957
transform 1 0 16192 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_176
timestamp 1688980957
transform 1 0 17296 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_192
timestamp 1688980957
transform 1 0 18768 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_237
timestamp 1688980957
transform 1 0 22908 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_244
timestamp 1688980957
transform 1 0 23552 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1688980957
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_261
timestamp 1688980957
transform 1 0 25116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_278
timestamp 1688980957
transform 1 0 26680 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_291
timestamp 1688980957
transform 1 0 27876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_303
timestamp 1688980957
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_89
timestamp 1688980957
transform 1 0 9292 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_119
timestamp 1688980957
transform 1 0 12052 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_129
timestamp 1688980957
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_133
timestamp 1688980957
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_187
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_196
timestamp 1688980957
transform 1 0 19136 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_203
timestamp 1688980957
transform 1 0 19780 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_211
timestamp 1688980957
transform 1 0 20516 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_216
timestamp 1688980957
transform 1 0 20976 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_228
timestamp 1688980957
transform 1 0 22080 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_234
timestamp 1688980957
transform 1 0 22632 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_259
timestamp 1688980957
transform 1 0 24932 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_272
timestamp 1688980957
transform 1 0 26128 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_367
timestamp 1688980957
transform 1 0 34868 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_99
timestamp 1688980957
transform 1 0 10212 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_136
timestamp 1688980957
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_149
timestamp 1688980957
transform 1 0 14812 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_166
timestamp 1688980957
transform 1 0 16376 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_187
timestamp 1688980957
transform 1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_217
timestamp 1688980957
transform 1 0 21068 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_231
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_239
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_250
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_258
timestamp 1688980957
transform 1 0 24840 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_272
timestamp 1688980957
transform 1 0 26128 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_284
timestamp 1688980957
transform 1 0 27232 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_296
timestamp 1688980957
transform 1 0 28336 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_104
timestamp 1688980957
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_117
timestamp 1688980957
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_126
timestamp 1688980957
transform 1 0 12696 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_134
timestamp 1688980957
transform 1 0 13432 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_146
timestamp 1688980957
transform 1 0 14536 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_184
timestamp 1688980957
transform 1 0 18032 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_196
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_206
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_222
timestamp 1688980957
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_367
timestamp 1688980957
transform 1 0 34868 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_89
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_94
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_102
timestamp 1688980957
transform 1 0 10488 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_113
timestamp 1688980957
transform 1 0 11500 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_128
timestamp 1688980957
transform 1 0 12880 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_138
timestamp 1688980957
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_147
timestamp 1688980957
transform 1 0 14628 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_155
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_167
timestamp 1688980957
transform 1 0 16468 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_182
timestamp 1688980957
transform 1 0 17848 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_223
timestamp 1688980957
transform 1 0 21620 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_235
timestamp 1688980957
transform 1 0 22724 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_262
timestamp 1688980957
transform 1 0 25208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_292
timestamp 1688980957
transform 1 0 27968 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_304
timestamp 1688980957
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_106
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1688980957
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1688980957
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_234
timestamp 1688980957
transform 1 0 22632 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_238
timestamp 1688980957
transform 1 0 23000 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_251
timestamp 1688980957
transform 1 0 24196 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_268
timestamp 1688980957
transform 1 0 25760 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_297
timestamp 1688980957
transform 1 0 28428 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_309
timestamp 1688980957
transform 1 0 29532 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_321
timestamp 1688980957
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_333
timestamp 1688980957
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_367
timestamp 1688980957
transform 1 0 34868 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_99
timestamp 1688980957
transform 1 0 10212 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_111
timestamp 1688980957
transform 1 0 11316 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_123
timestamp 1688980957
transform 1 0 12420 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_135
timestamp 1688980957
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_151
timestamp 1688980957
transform 1 0 14996 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_155
timestamp 1688980957
transform 1 0 15364 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_167
timestamp 1688980957
transform 1 0 16468 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_182
timestamp 1688980957
transform 1 0 17848 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_194
timestamp 1688980957
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_235
timestamp 1688980957
transform 1 0 22724 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_247
timestamp 1688980957
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_89
timestamp 1688980957
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_106
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_133
timestamp 1688980957
transform 1 0 13340 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_145
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_153
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_160
timestamp 1688980957
transform 1 0 15824 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_179
timestamp 1688980957
transform 1 0 17572 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_187
timestamp 1688980957
transform 1 0 18308 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_194
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_206
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_222
timestamp 1688980957
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_234
timestamp 1688980957
transform 1 0 22632 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_246
timestamp 1688980957
transform 1 0 23736 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_258
timestamp 1688980957
transform 1 0 24840 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_270
timestamp 1688980957
transform 1 0 25944 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_278
timestamp 1688980957
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_114
timestamp 1688980957
transform 1 0 11592 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_118
timestamp 1688980957
transform 1 0 11960 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_125
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_157
timestamp 1688980957
transform 1 0 15548 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_179
timestamp 1688980957
transform 1 0 17572 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_207
timestamp 1688980957
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_219
timestamp 1688980957
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_231
timestamp 1688980957
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_243
timestamp 1688980957
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_131
timestamp 1688980957
transform 1 0 13156 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_143
timestamp 1688980957
transform 1 0 14260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_162
timestamp 1688980957
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_187
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_192
timestamp 1688980957
transform 1 0 18768 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_204
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_210
timestamp 1688980957
transform 1 0 20424 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_367
timestamp 1688980957
transform 1 0 34868 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_117
timestamp 1688980957
transform 1 0 11868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_172
timestamp 1688980957
transform 1 0 16928 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_191
timestamp 1688980957
transform 1 0 18676 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_203
timestamp 1688980957
transform 1 0 19780 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_215
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_367
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 1688980957
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_367
timestamp 1688980957
transform 1 0 34868 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 1688980957
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1688980957
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_367
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1688980957
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_367
timestamp 1688980957
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_367
timestamp 1688980957
transform 1 0 34868 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_367
timestamp 1688980957
transform 1 0 34868 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_367
timestamp 1688980957
transform 1 0 34868 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 1688980957
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 1688980957
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 1688980957
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_367
timestamp 1688980957
transform 1 0 34868 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_367
timestamp 1688980957
transform 1 0 34868 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_367
timestamp 1688980957
transform 1 0 34868 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_367
timestamp 1688980957
transform 1 0 34868 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_367
timestamp 1688980957
transform 1 0 34868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_367
timestamp 1688980957
transform 1 0 34868 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_367
timestamp 1688980957
transform 1 0 34868 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_367
timestamp 1688980957
transform 1 0 34868 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_69
timestamp 1688980957
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_81
timestamp 1688980957
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_113
timestamp 1688980957
transform 1 0 11500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_125
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_169
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_181
timestamp 1688980957
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_237
timestamp 1688980957
transform 1 0 22908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_249
timestamp 1688980957
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_281
timestamp 1688980957
transform 1 0 26956 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_293
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_305
timestamp 1688980957
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_337
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_349
timestamp 1688980957
transform 1 0 33212 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_361
timestamp 1688980957
transform 1 0 34316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1688980957
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 2300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 14168 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform -1 0 34960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34592 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_12  output20 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16744 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 1688980957
transform 1 0 31004 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 1688980957
transform 1 0 32476 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 1688980957
transform 1 0 18216 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 1688980957
transform -1 0 22172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 1688980957
transform -1 0 23736 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 1688980957
transform 1 0 23736 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 1688980957
transform -1 0 25852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 1688980957
transform -1 0 26772 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output35
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 35236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 35236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 35236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 35236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 35236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 35236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 35236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 35236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 35236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 35236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 35236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 35236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 35236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 35236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 35236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 35236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 35236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 35236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 35236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 35236 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 35236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 35236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 35236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 35236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 35236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 35236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 35236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 35236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 35236 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 35236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 35236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 35236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 35236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 35236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 35236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 35236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 35236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 35236 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 35236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 35236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 35236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 35236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 35236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 35236 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 35236 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 35236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 35236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 35236 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 11408 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 21712 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 32016 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
<< labels >>
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 a[0]
port 0 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 a[1]
port 1 nsew signal input
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 a[2]
port 2 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 a[3]
port 3 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 a[4]
port 4 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 a[5]
port 5 nsew signal input
flabel metal2 s 13082 0 13138 800 0 FreeSans 224 90 0 0 a[6]
port 6 nsew signal input
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 a[7]
port 7 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 b[0]
port 8 nsew signal input
flabel metal2 s 3974 0 4030 800 0 FreeSans 224 90 0 0 b[1]
port 9 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 b[2]
port 10 nsew signal input
flabel metal2 s 8022 0 8078 800 0 FreeSans 224 90 0 0 b[3]
port 11 nsew signal input
flabel metal2 s 10046 0 10102 800 0 FreeSans 224 90 0 0 b[4]
port 12 nsew signal input
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 b[5]
port 13 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 b[6]
port 14 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 b[7]
port 15 nsew signal input
flabel metal2 s 33322 0 33378 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 control
port 17 nsew signal input
flabel metal2 s 17130 0 17186 800 0 FreeSans 224 90 0 0 p[0]
port 18 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 p[10]
port 19 nsew signal tristate
flabel metal2 s 28262 0 28318 800 0 FreeSans 224 90 0 0 p[11]
port 20 nsew signal tristate
flabel metal2 s 29274 0 29330 800 0 FreeSans 224 90 0 0 p[12]
port 21 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 p[13]
port 22 nsew signal tristate
flabel metal2 s 31298 0 31354 800 0 FreeSans 224 90 0 0 p[14]
port 23 nsew signal tristate
flabel metal2 s 32310 0 32366 800 0 FreeSans 224 90 0 0 p[15]
port 24 nsew signal tristate
flabel metal2 s 18142 0 18198 800 0 FreeSans 224 90 0 0 p[1]
port 25 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 p[2]
port 26 nsew signal tristate
flabel metal2 s 20166 0 20222 800 0 FreeSans 224 90 0 0 p[3]
port 27 nsew signal tristate
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 p[4]
port 28 nsew signal tristate
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 p[5]
port 29 nsew signal tristate
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 p[6]
port 30 nsew signal tristate
flabel metal2 s 24214 0 24270 800 0 FreeSans 224 90 0 0 p[7]
port 31 nsew signal tristate
flabel metal2 s 25226 0 25282 800 0 FreeSans 224 90 0 0 p[8]
port 32 nsew signal tristate
flabel metal2 s 26238 0 26294 800 0 FreeSans 224 90 0 0 p[9]
port 33 nsew signal tristate
flabel metal2 s 34334 0 34390 800 0 FreeSans 224 90 0 0 rst
port 34 nsew signal input
flabel metal4 s 4208 2128 4528 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 34928 2128 35248 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 19568 2128 19888 36496 0 FreeSans 1920 90 0 0 vssd1
port 36 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36400 38800
<< end >>
