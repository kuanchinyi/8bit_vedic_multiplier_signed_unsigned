magic
tech sky130A
magscale 1 2
timestamp 1726925974
<< viali >>
rect 1409 36125 1443 36159
rect 33149 36125 33183 36159
rect 34345 36057 34379 36091
rect 1593 35989 1627 36023
rect 1409 35037 1443 35071
rect 1593 34901 1627 34935
rect 33149 33949 33183 33983
rect 34345 33881 34379 33915
rect 1409 32861 1443 32895
rect 1593 32725 1627 32759
rect 33149 31773 33183 31807
rect 34345 31705 34379 31739
rect 1409 30685 1443 30719
rect 1593 30549 1627 30583
rect 33149 29597 33183 29631
rect 34345 29529 34379 29563
rect 1409 28509 1443 28543
rect 1593 28373 1627 28407
rect 23673 28373 23707 28407
rect 23673 28169 23707 28203
rect 25605 28169 25639 28203
rect 5917 28033 5951 28067
rect 6561 28033 6595 28067
rect 21649 28033 21683 28067
rect 21925 28033 21959 28067
rect 23857 28033 23891 28067
rect 22201 27965 22235 27999
rect 24133 27965 24167 27999
rect 6009 27829 6043 27863
rect 5162 27625 5196 27659
rect 12817 27625 12851 27659
rect 22017 27625 22051 27659
rect 22661 27625 22695 27659
rect 23857 27625 23891 27659
rect 21373 27557 21407 27591
rect 23029 27557 23063 27591
rect 4905 27489 4939 27523
rect 12449 27489 12483 27523
rect 18429 27489 18463 27523
rect 19349 27489 19383 27523
rect 19809 27489 19843 27523
rect 24409 27489 24443 27523
rect 4537 27421 4571 27455
rect 4629 27421 4663 27455
rect 12541 27421 12575 27455
rect 13001 27421 13035 27455
rect 13185 27421 13219 27455
rect 14105 27421 14139 27455
rect 14289 27421 14323 27455
rect 14657 27421 14691 27455
rect 14841 27421 14875 27455
rect 18337 27421 18371 27455
rect 18521 27421 18555 27455
rect 19441 27421 19475 27455
rect 21465 27421 21499 27455
rect 21557 27421 21591 27455
rect 21741 27421 21775 27455
rect 21833 27421 21867 27455
rect 22099 27431 22133 27465
rect 22201 27421 22235 27455
rect 22385 27421 22419 27455
rect 22477 27421 22511 27455
rect 22937 27421 22971 27455
rect 24041 27421 24075 27455
rect 33241 27421 33275 27455
rect 6929 27353 6963 27387
rect 14197 27353 14231 27387
rect 23489 27353 23523 27387
rect 24685 27353 24719 27387
rect 34345 27353 34379 27387
rect 4721 27285 4755 27319
rect 7205 27285 7239 27319
rect 13001 27285 13035 27319
rect 14749 27285 14783 27319
rect 24133 27285 24167 27319
rect 26157 27285 26191 27319
rect 12081 27081 12115 27115
rect 14933 27081 14967 27115
rect 16313 27081 16347 27115
rect 19165 27081 19199 27115
rect 19257 27081 19291 27115
rect 19441 27081 19475 27115
rect 25513 27081 25547 27115
rect 12817 27013 12851 27047
rect 13369 27013 13403 27047
rect 16681 27013 16715 27047
rect 16881 27013 16915 27047
rect 18213 27013 18247 27047
rect 18429 27013 18463 27047
rect 21465 27013 21499 27047
rect 3893 26945 3927 26979
rect 11897 26945 11931 26979
rect 12081 26945 12115 26979
rect 12357 26945 12391 26979
rect 12541 26945 12575 26979
rect 13001 26945 13035 26979
rect 13093 26945 13127 26979
rect 13185 26945 13219 26979
rect 14013 26945 14047 26979
rect 14105 26945 14139 26979
rect 14381 26945 14415 26979
rect 14657 26945 14691 26979
rect 14841 26945 14875 26979
rect 15117 26945 15151 26979
rect 15393 26945 15427 26979
rect 15577 26945 15611 26979
rect 15945 26945 15979 26979
rect 17417 26945 17451 26979
rect 17785 26945 17819 26979
rect 17969 26945 18003 26979
rect 18613 26945 18647 26979
rect 18705 26945 18739 26979
rect 18889 26945 18923 26979
rect 18981 26945 19015 26979
rect 20177 26945 20211 26979
rect 20637 26945 20671 26979
rect 21097 26945 21131 26979
rect 21251 26945 21285 26979
rect 22017 26945 22051 26979
rect 24409 26945 24443 26979
rect 25145 26945 25179 26979
rect 25421 26945 25455 26979
rect 4169 26877 4203 26911
rect 5917 26877 5951 26911
rect 12173 26877 12207 26911
rect 12633 26877 12667 26911
rect 14289 26877 14323 26911
rect 15301 26877 15335 26911
rect 15853 26877 15887 26911
rect 17141 26877 17175 26911
rect 17509 26877 17543 26911
rect 21005 26877 21039 26911
rect 21925 26877 21959 26911
rect 22385 26877 22419 26911
rect 13369 26809 13403 26843
rect 14473 26809 14507 26843
rect 17049 26809 17083 26843
rect 17325 26809 17359 26843
rect 17601 26809 17635 26843
rect 18061 26809 18095 26843
rect 19809 26809 19843 26843
rect 6561 26741 6595 26775
rect 14197 26741 14231 26775
rect 15393 26741 15427 26775
rect 16865 26741 16899 26775
rect 17417 26741 17451 26775
rect 18245 26741 18279 26775
rect 19441 26741 19475 26775
rect 22661 26741 22695 26775
rect 25237 26741 25271 26775
rect 25973 26741 26007 26775
rect 26249 26741 26283 26775
rect 6009 26537 6043 26571
rect 6377 26537 6411 26571
rect 12541 26537 12575 26571
rect 14197 26537 14231 26571
rect 15761 26537 15795 26571
rect 24133 26537 24167 26571
rect 15485 26469 15519 26503
rect 16221 26469 16255 26503
rect 17509 26469 17543 26503
rect 22937 26469 22971 26503
rect 11805 26401 11839 26435
rect 12173 26401 12207 26435
rect 15393 26401 15427 26435
rect 22753 26401 22787 26435
rect 24409 26401 24443 26435
rect 26157 26401 26191 26435
rect 1409 26333 1443 26367
rect 5273 26333 5307 26367
rect 5733 26333 5767 26367
rect 11713 26333 11747 26367
rect 11897 26333 11931 26367
rect 12081 26333 12115 26367
rect 12357 26333 12391 26367
rect 14197 26333 14231 26367
rect 14381 26333 14415 26367
rect 15117 26333 15151 26367
rect 15301 26333 15335 26367
rect 15577 26333 15611 26367
rect 15945 26333 15979 26367
rect 16037 26333 16071 26367
rect 16957 26333 16991 26367
rect 17141 26333 17175 26367
rect 17233 26333 17267 26367
rect 17877 26333 17911 26367
rect 18061 26333 18095 26367
rect 23029 26333 23063 26367
rect 5365 26265 5399 26299
rect 16221 26265 16255 26299
rect 17049 26265 17083 26299
rect 17509 26265 17543 26299
rect 17969 26265 18003 26299
rect 22753 26265 22787 26299
rect 24685 26265 24719 26299
rect 1593 26197 1627 26231
rect 5641 26197 5675 26231
rect 15025 26197 15059 26231
rect 17325 26197 17359 26231
rect 14013 25993 14047 26027
rect 15485 25993 15519 26027
rect 22201 25993 22235 26027
rect 23673 25993 23707 26027
rect 4537 25925 4571 25959
rect 10977 25925 11011 25959
rect 11621 25925 11655 25959
rect 16221 25925 16255 25959
rect 26065 25925 26099 25959
rect 10701 25857 10735 25891
rect 10793 25857 10827 25891
rect 11161 25857 11195 25891
rect 11345 25857 11379 25891
rect 11805 25857 11839 25891
rect 11989 25857 12023 25891
rect 12357 25857 12391 25891
rect 13001 25857 13035 25891
rect 13829 25857 13863 25891
rect 14105 25857 14139 25891
rect 14289 25857 14323 25891
rect 15393 25857 15427 25891
rect 15577 25857 15611 25891
rect 15669 25857 15703 25891
rect 15761 25857 15795 25891
rect 15945 25857 15979 25891
rect 17325 25857 17359 25891
rect 20085 25857 20119 25891
rect 20269 25857 20303 25891
rect 20453 25857 20487 25891
rect 20913 25857 20947 25891
rect 22385 25857 22419 25891
rect 22477 25857 22511 25891
rect 22661 25857 22695 25891
rect 22753 25857 22787 25891
rect 22845 25857 22879 25891
rect 23489 25857 23523 25891
rect 23949 25857 23983 25891
rect 24133 25857 24167 25891
rect 26157 25857 26191 25891
rect 4261 25789 4295 25823
rect 11253 25789 11287 25823
rect 12173 25789 12207 25823
rect 12541 25789 12575 25823
rect 12909 25789 12943 25823
rect 13645 25789 13679 25823
rect 14197 25789 14231 25823
rect 17233 25789 17267 25823
rect 21005 25789 21039 25823
rect 22937 25789 22971 25823
rect 23305 25789 23339 25823
rect 24409 25789 24443 25823
rect 25881 25789 25915 25823
rect 6009 25721 6043 25755
rect 13369 25721 13403 25755
rect 15853 25721 15887 25755
rect 21281 25721 21315 25755
rect 23213 25721 23247 25755
rect 6561 25653 6595 25687
rect 10057 25653 10091 25687
rect 17693 25653 17727 25687
rect 22109 25653 22143 25687
rect 23029 25653 23063 25687
rect 26433 25653 26467 25687
rect 8033 25449 8067 25483
rect 10149 25449 10183 25483
rect 10609 25449 10643 25483
rect 11069 25449 11103 25483
rect 11805 25449 11839 25483
rect 12633 25449 12667 25483
rect 12817 25449 12851 25483
rect 15945 25449 15979 25483
rect 17969 25449 18003 25483
rect 20177 25449 20211 25483
rect 21281 25449 21315 25483
rect 23305 25449 23339 25483
rect 7209 25381 7243 25415
rect 10977 25381 11011 25415
rect 16313 25381 16347 25415
rect 18245 25381 18279 25415
rect 18613 25381 18647 25415
rect 18889 25381 18923 25415
rect 21925 25381 21959 25415
rect 23489 25381 23523 25415
rect 4445 25313 4479 25347
rect 7941 25313 7975 25347
rect 11253 25313 11287 25347
rect 11713 25313 11747 25347
rect 12173 25313 12207 25347
rect 14749 25313 14783 25347
rect 18061 25313 18095 25347
rect 18521 25313 18555 25347
rect 21465 25313 21499 25347
rect 22937 25313 22971 25347
rect 4169 25245 4203 25279
rect 7113 25245 7147 25279
rect 7297 25245 7331 25279
rect 7389 25245 7423 25279
rect 7849 25245 7883 25279
rect 10609 25245 10643 25279
rect 10793 25245 10827 25279
rect 11345 25245 11379 25279
rect 11989 25245 12023 25279
rect 12265 25245 12299 25279
rect 12541 25245 12575 25279
rect 15301 25245 15335 25279
rect 15485 25245 15519 25279
rect 15577 25245 15611 25279
rect 15669 25245 15703 25279
rect 16037 25245 16071 25279
rect 16221 25245 16255 25279
rect 16681 25245 16715 25279
rect 18245 25245 18279 25279
rect 18429 25245 18463 25279
rect 18705 25245 18739 25279
rect 20085 25245 20119 25279
rect 20361 25245 20395 25279
rect 20453 25245 20487 25279
rect 20637 25245 20671 25279
rect 20729 25245 20763 25279
rect 20821 25245 20855 25279
rect 21097 25245 21131 25279
rect 21557 25245 21591 25279
rect 23029 25245 23063 25279
rect 23489 25245 23523 25279
rect 23673 25245 23707 25279
rect 23949 25245 23983 25279
rect 33149 25245 33183 25279
rect 6193 25177 6227 25211
rect 8125 25177 8159 25211
rect 10333 25177 10367 25211
rect 11621 25177 11655 25211
rect 17877 25177 17911 25211
rect 19717 25177 19751 25211
rect 19901 25177 19935 25211
rect 34345 25177 34379 25211
rect 6469 25109 6503 25143
rect 6929 25109 6963 25143
rect 7665 25109 7699 25143
rect 9781 25109 9815 25143
rect 15117 25109 15151 25143
rect 20913 25109 20947 25143
rect 11161 24905 11195 24939
rect 12081 24905 12115 24939
rect 12725 24905 12759 24939
rect 13921 24905 13955 24939
rect 15301 24905 15335 24939
rect 19809 24905 19843 24939
rect 21005 24905 21039 24939
rect 12449 24837 12483 24871
rect 5181 24769 5215 24803
rect 5641 24769 5675 24803
rect 6929 24769 6963 24803
rect 7481 24769 7515 24803
rect 8493 24769 8527 24803
rect 9229 24769 9263 24803
rect 10609 24769 10643 24803
rect 12633 24769 12667 24803
rect 12817 24769 12851 24803
rect 13645 24769 13679 24803
rect 14013 24769 14047 24803
rect 14565 24769 14599 24803
rect 14657 24769 14691 24803
rect 15485 24769 15519 24803
rect 15639 24769 15673 24803
rect 16221 24769 16255 24803
rect 19257 24769 19291 24803
rect 19717 24769 19751 24803
rect 19901 24769 19935 24803
rect 20545 24769 20579 24803
rect 21189 24769 21223 24803
rect 10701 24701 10735 24735
rect 13921 24701 13955 24735
rect 14105 24701 14139 24735
rect 14841 24701 14875 24735
rect 15853 24701 15887 24735
rect 15945 24701 15979 24735
rect 19165 24701 19199 24735
rect 20453 24701 20487 24735
rect 20913 24701 20947 24735
rect 21373 24701 21407 24735
rect 8309 24633 8343 24667
rect 13737 24633 13771 24667
rect 14381 24633 14415 24667
rect 16037 24633 16071 24667
rect 19625 24633 19659 24667
rect 5273 24565 5307 24599
rect 6101 24565 6135 24599
rect 14197 24565 14231 24599
rect 16129 24565 16163 24599
rect 11161 24361 11195 24395
rect 11621 24361 11655 24395
rect 11897 24361 11931 24395
rect 12173 24361 12207 24395
rect 12541 24361 12575 24395
rect 13645 24361 13679 24395
rect 14289 24361 14323 24395
rect 15301 24361 15335 24395
rect 17601 24361 17635 24395
rect 18521 24361 18555 24395
rect 18613 24361 18647 24395
rect 24133 24361 24167 24395
rect 6653 24293 6687 24327
rect 13829 24293 13863 24327
rect 15669 24293 15703 24327
rect 18705 24293 18739 24327
rect 6193 24225 6227 24259
rect 9229 24225 9263 24259
rect 11805 24225 11839 24259
rect 11897 24225 11931 24259
rect 12081 24225 12115 24259
rect 12449 24225 12483 24259
rect 17049 24225 17083 24259
rect 17325 24225 17359 24259
rect 18245 24225 18279 24259
rect 24409 24225 24443 24259
rect 1409 24157 1443 24191
rect 4169 24157 4203 24191
rect 6561 24157 6595 24191
rect 6745 24157 6779 24191
rect 7481 24157 7515 24191
rect 8033 24157 8067 24191
rect 9137 24157 9171 24191
rect 11345 24157 11379 24191
rect 11437 24157 11471 24191
rect 11713 24157 11747 24191
rect 12541 24157 12575 24191
rect 12633 24157 12667 24191
rect 12817 24157 12851 24191
rect 13001 24157 13035 24191
rect 13185 24157 13219 24191
rect 13277 24157 13311 24191
rect 13369 24157 13403 24191
rect 13737 24157 13771 24191
rect 13921 24157 13955 24191
rect 15209 24157 15243 24191
rect 16957 24157 16991 24191
rect 17417 24157 17451 24191
rect 17601 24157 17635 24191
rect 18153 24157 18187 24191
rect 4445 24089 4479 24123
rect 11161 24089 11195 24123
rect 12725 24089 12759 24123
rect 14105 24089 14139 24123
rect 19073 24089 19107 24123
rect 24685 24089 24719 24123
rect 1593 24021 1627 24055
rect 9505 24021 9539 24055
rect 14305 24021 14339 24055
rect 14473 24021 14507 24055
rect 26157 24021 26191 24055
rect 13829 23817 13863 23851
rect 20913 23817 20947 23851
rect 24961 23817 24995 23851
rect 9137 23749 9171 23783
rect 12357 23749 12391 23783
rect 23121 23749 23155 23783
rect 6653 23681 6687 23715
rect 7389 23681 7423 23715
rect 7665 23681 7699 23715
rect 8033 23681 8067 23715
rect 8401 23681 8435 23715
rect 8953 23681 8987 23715
rect 9873 23681 9907 23715
rect 10517 23681 10551 23715
rect 12265 23681 12299 23715
rect 12449 23681 12483 23715
rect 12817 23681 12851 23715
rect 12909 23681 12943 23715
rect 13093 23681 13127 23715
rect 13185 23681 13219 23715
rect 13737 23681 13771 23715
rect 20637 23681 20671 23715
rect 21097 23681 21131 23715
rect 22017 23681 22051 23715
rect 22845 23681 22879 23715
rect 23029 23681 23063 23715
rect 23213 23681 23247 23715
rect 23489 23681 23523 23715
rect 24869 23681 24903 23715
rect 3985 23613 4019 23647
rect 4261 23613 4295 23647
rect 6009 23613 6043 23647
rect 13369 23613 13403 23647
rect 20453 23613 20487 23647
rect 21373 23613 21407 23647
rect 21925 23613 21959 23647
rect 23581 23613 23615 23647
rect 23857 23613 23891 23647
rect 7113 23545 7147 23579
rect 20821 23545 20855 23579
rect 21281 23545 21315 23579
rect 22385 23545 22419 23579
rect 11345 23477 11379 23511
rect 25421 23477 25455 23511
rect 5089 23273 5123 23307
rect 7113 23273 7147 23307
rect 13093 23273 13127 23307
rect 16221 23273 16255 23307
rect 20085 23273 20119 23307
rect 21649 23273 21683 23307
rect 22569 23273 22603 23307
rect 4905 23205 4939 23239
rect 12173 23205 12207 23239
rect 21005 23205 21039 23239
rect 21465 23205 21499 23239
rect 6837 23137 6871 23171
rect 8033 23137 8067 23171
rect 15301 23137 15335 23171
rect 16681 23137 16715 23171
rect 19717 23137 19751 23171
rect 21189 23137 21223 23171
rect 4997 23069 5031 23103
rect 6929 23069 6963 23103
rect 7941 23069 7975 23103
rect 9781 23069 9815 23103
rect 10425 23069 10459 23103
rect 12081 23069 12115 23103
rect 12357 23069 12391 23103
rect 12466 23069 12500 23103
rect 12633 23069 12667 23103
rect 13185 23069 13219 23103
rect 13369 23069 13403 23103
rect 15393 23069 15427 23103
rect 16037 23069 16071 23103
rect 16497 23069 16531 23103
rect 16773 23069 16807 23103
rect 19809 23069 19843 23103
rect 20821 23069 20855 23103
rect 33149 23069 33183 23103
rect 12725 23001 12759 23035
rect 12909 23001 12943 23035
rect 16405 23001 16439 23035
rect 20637 23001 20671 23035
rect 34345 23001 34379 23035
rect 5641 22933 5675 22967
rect 6101 22933 6135 22967
rect 8309 22933 8343 22967
rect 13277 22933 13311 22967
rect 15761 22933 15795 22967
rect 17141 22933 17175 22967
rect 6009 22729 6043 22763
rect 10241 22729 10275 22763
rect 14841 22729 14875 22763
rect 15669 22729 15703 22763
rect 19349 22729 19383 22763
rect 22661 22729 22695 22763
rect 23397 22729 23431 22763
rect 23857 22729 23891 22763
rect 3893 22661 3927 22695
rect 5641 22661 5675 22695
rect 9781 22661 9815 22695
rect 25881 22661 25915 22695
rect 5733 22593 5767 22627
rect 6561 22593 6595 22627
rect 7021 22593 7055 22627
rect 7941 22593 7975 22627
rect 8585 22593 8619 22627
rect 10517 22593 10551 22627
rect 14381 22593 14415 22627
rect 14657 22593 14691 22627
rect 14933 22593 14967 22627
rect 15301 22593 15335 22627
rect 15393 22593 15427 22627
rect 15761 22593 15795 22627
rect 15945 22593 15979 22627
rect 17785 22593 17819 22627
rect 18245 22593 18279 22627
rect 18429 22593 18463 22627
rect 18705 22593 18739 22627
rect 19563 22593 19597 22627
rect 19717 22593 19751 22627
rect 22753 22593 22787 22627
rect 22937 22593 22971 22627
rect 23213 22593 23247 22627
rect 23949 22593 23983 22627
rect 25973 22593 26007 22627
rect 26249 22593 26283 22627
rect 3617 22525 3651 22559
rect 5365 22525 5399 22559
rect 6469 22525 6503 22559
rect 10333 22525 10367 22559
rect 14473 22525 14507 22559
rect 15117 22525 15151 22559
rect 15209 22525 15243 22559
rect 15853 22525 15887 22559
rect 17693 22525 17727 22559
rect 18153 22525 18187 22559
rect 18797 22525 18831 22559
rect 19073 22525 19107 22559
rect 24225 22525 24259 22559
rect 25697 22525 25731 22559
rect 9781 22457 9815 22491
rect 14381 22389 14415 22423
rect 18245 22389 18279 22423
rect 5825 22185 5859 22219
rect 10333 22185 10367 22219
rect 11529 22185 11563 22219
rect 15393 22185 15427 22219
rect 18245 22185 18279 22219
rect 20637 22185 20671 22219
rect 21465 22185 21499 22219
rect 23305 22185 23339 22219
rect 7849 22117 7883 22151
rect 9137 22117 9171 22151
rect 10885 22117 10919 22151
rect 13001 22117 13035 22151
rect 20821 22117 20855 22151
rect 21097 22117 21131 22151
rect 22201 22117 22235 22151
rect 10241 22049 10275 22083
rect 11161 22049 11195 22083
rect 20361 22049 20395 22083
rect 21741 22049 21775 22083
rect 23121 22049 23155 22083
rect 1409 21981 1443 22015
rect 5549 21981 5583 22015
rect 5641 21981 5675 22015
rect 6009 21981 6043 22015
rect 6377 21981 6411 22015
rect 7941 21981 7975 22015
rect 8125 21981 8159 22015
rect 8309 21981 8343 22015
rect 9137 21981 9171 22015
rect 9505 21981 9539 22015
rect 9873 21981 9907 22015
rect 10149 21981 10183 22015
rect 10425 21981 10459 22015
rect 10793 21981 10827 22015
rect 10977 21981 11011 22015
rect 11069 21981 11103 22015
rect 11345 21981 11379 22015
rect 12725 21981 12759 22015
rect 13553 21981 13587 22015
rect 13737 21981 13771 22015
rect 14749 21981 14783 22015
rect 14933 21981 14967 22015
rect 15025 21981 15059 22015
rect 15117 21981 15151 22015
rect 16405 21981 16439 22015
rect 18245 21981 18279 22015
rect 18429 21981 18463 22015
rect 18521 21981 18555 22015
rect 19901 21981 19935 22015
rect 20177 21981 20211 22015
rect 21005 21981 21039 22015
rect 21281 21981 21315 22015
rect 21833 21981 21867 22015
rect 23029 21981 23063 22015
rect 5825 21913 5859 21947
rect 13011 21913 13045 21947
rect 16129 21913 16163 21947
rect 16313 21913 16347 21947
rect 20453 21913 20487 21947
rect 1593 21845 1627 21879
rect 5365 21845 5399 21879
rect 10609 21845 10643 21879
rect 12817 21845 12851 21879
rect 13645 21845 13679 21879
rect 16405 21845 16439 21879
rect 19993 21845 20027 21879
rect 20653 21845 20687 21879
rect 6469 21641 6503 21675
rect 10241 21641 10275 21675
rect 11253 21641 11287 21675
rect 16037 21641 16071 21675
rect 16773 21641 16807 21675
rect 17417 21641 17451 21675
rect 18061 21641 18095 21675
rect 21005 21641 21039 21675
rect 21649 21641 21683 21675
rect 23029 21641 23063 21675
rect 4077 21573 4111 21607
rect 9413 21573 9447 21607
rect 10885 21573 10919 21607
rect 12633 21573 12667 21607
rect 15761 21573 15795 21607
rect 17509 21573 17543 21607
rect 17709 21573 17743 21607
rect 21189 21573 21223 21607
rect 22477 21573 22511 21607
rect 6101 21505 6135 21539
rect 6644 21505 6678 21539
rect 6745 21505 6779 21539
rect 6929 21505 6963 21539
rect 7941 21505 7975 21539
rect 8677 21505 8711 21539
rect 9965 21505 9999 21539
rect 10701 21505 10735 21539
rect 10977 21505 11011 21539
rect 11069 21505 11103 21539
rect 12725 21505 12759 21539
rect 13645 21505 13679 21539
rect 13737 21505 13771 21539
rect 14473 21505 14507 21539
rect 15393 21505 15427 21539
rect 15577 21505 15611 21539
rect 15945 21505 15979 21539
rect 16221 21505 16255 21539
rect 17049 21505 17083 21539
rect 17969 21505 18003 21539
rect 18245 21505 18279 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 22017 21505 22051 21539
rect 22201 21505 22235 21539
rect 22293 21505 22327 21539
rect 22753 21505 22787 21539
rect 23305 21505 23339 21539
rect 3801 21437 3835 21471
rect 5825 21437 5859 21471
rect 10057 21437 10091 21471
rect 10333 21437 10367 21471
rect 10425 21437 10459 21471
rect 10609 21437 10643 21471
rect 11805 21437 11839 21471
rect 12909 21437 12943 21471
rect 13001 21437 13035 21471
rect 13369 21437 13403 21471
rect 13829 21437 13863 21471
rect 13921 21437 13955 21471
rect 14381 21437 14415 21471
rect 15301 21437 15335 21471
rect 16405 21437 16439 21471
rect 16957 21437 16991 21471
rect 21833 21437 21867 21471
rect 23029 21437 23063 21471
rect 6837 21369 6871 21403
rect 9781 21369 9815 21403
rect 9873 21369 9907 21403
rect 14105 21369 14139 21403
rect 21465 21369 21499 21403
rect 17693 21301 17727 21335
rect 17877 21301 17911 21335
rect 18245 21301 18279 21335
rect 22661 21301 22695 21335
rect 22845 21301 22879 21335
rect 4905 21097 4939 21131
rect 5365 21097 5399 21131
rect 10149 21097 10183 21131
rect 10885 21097 10919 21131
rect 13093 21097 13127 21131
rect 13553 21097 13587 21131
rect 13737 21097 13771 21131
rect 14565 21097 14599 21131
rect 15577 21097 15611 21131
rect 16405 21097 16439 21131
rect 18429 21097 18463 21131
rect 20269 21097 20303 21131
rect 20545 21097 20579 21131
rect 24133 21097 24167 21131
rect 6561 21029 6595 21063
rect 7297 20961 7331 20995
rect 8953 20961 8987 20995
rect 14933 20961 14967 20995
rect 15393 20961 15427 20995
rect 16037 20961 16071 20995
rect 22753 20961 22787 20995
rect 23213 20961 23247 20995
rect 24685 20961 24719 20995
rect 4813 20893 4847 20927
rect 6285 20893 6319 20927
rect 7021 20893 7055 20927
rect 9321 20893 9355 20927
rect 9413 20893 9447 20927
rect 9873 20893 9907 20927
rect 10241 20893 10275 20927
rect 10333 20893 10367 20927
rect 10517 20893 10551 20927
rect 10701 20893 10735 20927
rect 13093 20893 13127 20927
rect 13461 20893 13495 20927
rect 14197 20893 14231 20927
rect 14289 20893 14323 20927
rect 14381 20893 14415 20927
rect 15301 20893 15335 20927
rect 16221 20893 16255 20927
rect 17969 20893 18003 20927
rect 18061 20893 18095 20927
rect 18429 20893 18463 20927
rect 19260 20871 19294 20905
rect 19533 20893 19567 20927
rect 19809 20893 19843 20927
rect 20085 20893 20119 20927
rect 20361 20893 20395 20927
rect 20637 20893 20671 20927
rect 22845 20893 22879 20927
rect 24409 20893 24443 20927
rect 33149 20893 33183 20927
rect 9045 20825 9079 20859
rect 10609 20825 10643 20859
rect 10977 20825 11011 20859
rect 11161 20825 11195 20859
rect 11345 20825 11379 20859
rect 13721 20825 13755 20859
rect 13921 20825 13955 20859
rect 15025 20825 15059 20859
rect 20453 20825 20487 20859
rect 34345 20825 34379 20859
rect 9597 20757 9631 20791
rect 9965 20757 9999 20791
rect 10057 20757 10091 20791
rect 13277 20757 13311 20791
rect 18613 20757 18647 20791
rect 19349 20757 19383 20791
rect 19717 20757 19751 20791
rect 19901 20757 19935 20791
rect 26157 20757 26191 20791
rect 10241 20553 10275 20587
rect 10333 20553 10367 20587
rect 10609 20553 10643 20587
rect 18889 20553 18923 20587
rect 18981 20553 19015 20587
rect 19717 20553 19751 20587
rect 25053 20553 25087 20587
rect 25421 20553 25455 20587
rect 8861 20485 8895 20519
rect 12725 20485 12759 20519
rect 19625 20485 19659 20519
rect 6837 20417 6871 20451
rect 7297 20417 7331 20451
rect 9229 20417 9263 20451
rect 9781 20417 9815 20451
rect 10517 20417 10551 20451
rect 10701 20417 10735 20451
rect 12541 20417 12575 20451
rect 13001 20417 13035 20451
rect 13185 20417 13219 20451
rect 15485 20417 15519 20451
rect 15853 20417 15887 20451
rect 18061 20417 18095 20451
rect 19073 20417 19107 20451
rect 19441 20417 19475 20451
rect 19717 20417 19751 20451
rect 24961 20417 24995 20451
rect 8953 20349 8987 20383
rect 9321 20349 9355 20383
rect 9873 20349 9907 20383
rect 9965 20349 9999 20383
rect 10057 20349 10091 20383
rect 16497 20349 16531 20383
rect 17693 20349 17727 20383
rect 17785 20349 17819 20383
rect 18153 20349 18187 20383
rect 18613 20349 18647 20383
rect 10885 20281 10919 20315
rect 12909 20281 12943 20315
rect 18337 20281 18371 20315
rect 9505 20213 9539 20247
rect 13185 20213 13219 20247
rect 9781 20009 9815 20043
rect 10793 20009 10827 20043
rect 11069 20009 11103 20043
rect 11621 20009 11655 20043
rect 13001 20009 13035 20043
rect 12449 19941 12483 19975
rect 12541 19941 12575 19975
rect 12909 19941 12943 19975
rect 16957 19941 16991 19975
rect 5825 19873 5859 19907
rect 10149 19873 10183 19907
rect 13093 19873 13127 19907
rect 13645 19873 13679 19907
rect 14289 19873 14323 19907
rect 1409 19805 1443 19839
rect 5733 19805 5767 19839
rect 6101 19805 6135 19839
rect 6285 19805 6319 19839
rect 7113 19805 7147 19839
rect 7481 19805 7515 19839
rect 9137 19805 9171 19839
rect 9321 19805 9355 19839
rect 9413 19805 9447 19839
rect 9505 19805 9539 19839
rect 10517 19805 10551 19839
rect 10609 19805 10643 19839
rect 10885 19805 10919 19839
rect 11161 19805 11195 19839
rect 11529 19805 11563 19839
rect 11989 19805 12023 19839
rect 12173 19805 12207 19839
rect 12633 19805 12667 19839
rect 13001 19805 13035 19839
rect 13277 19805 13311 19839
rect 13553 19805 13587 19839
rect 13737 19805 13771 19839
rect 14381 19805 14415 19839
rect 15209 19805 15243 19839
rect 19441 19805 19475 19839
rect 5089 19737 5123 19771
rect 8309 19737 8343 19771
rect 10241 19737 10275 19771
rect 11805 19737 11839 19771
rect 16589 19737 16623 19771
rect 19257 19737 19291 19771
rect 1593 19669 1627 19703
rect 11345 19669 11379 19703
rect 12265 19669 12299 19703
rect 13461 19669 13495 19703
rect 17049 19669 17083 19703
rect 19625 19669 19659 19703
rect 5917 19465 5951 19499
rect 12081 19465 12115 19499
rect 18245 19465 18279 19499
rect 19993 19465 20027 19499
rect 5733 19397 5767 19431
rect 7481 19397 7515 19431
rect 18797 19397 18831 19431
rect 6193 19329 6227 19363
rect 7665 19329 7699 19363
rect 8033 19329 8067 19363
rect 11069 19329 11103 19363
rect 11161 19329 11195 19363
rect 11805 19329 11839 19363
rect 11989 19329 12023 19363
rect 12265 19329 12299 19363
rect 12449 19329 12483 19363
rect 12541 19329 12575 19363
rect 12725 19329 12759 19363
rect 13553 19329 13587 19363
rect 13737 19329 13771 19363
rect 13921 19329 13955 19363
rect 16773 19329 16807 19363
rect 16957 19329 16991 19363
rect 17325 19329 17359 19363
rect 17785 19329 17819 19363
rect 17877 19329 17911 19363
rect 18061 19329 18095 19363
rect 18429 19329 18463 19363
rect 18613 19329 18647 19363
rect 19073 19329 19107 19363
rect 19533 19329 19567 19363
rect 19625 19329 19659 19363
rect 19809 19329 19843 19363
rect 6653 19261 6687 19295
rect 9505 19261 9539 19295
rect 12909 19261 12943 19295
rect 13001 19261 13035 19295
rect 17233 19261 17267 19295
rect 17693 19261 17727 19295
rect 18981 19261 19015 19295
rect 12633 19193 12667 19227
rect 13277 19193 13311 19227
rect 16773 19193 16807 19227
rect 17049 19193 17083 19227
rect 5917 19125 5951 19159
rect 13461 19125 13495 19159
rect 19349 19125 19383 19159
rect 8033 18921 8067 18955
rect 8401 18921 8435 18955
rect 15485 18921 15519 18955
rect 17233 18921 17267 18955
rect 17693 18921 17727 18955
rect 20085 18853 20119 18887
rect 21005 18853 21039 18887
rect 3893 18785 3927 18819
rect 4169 18785 4203 18819
rect 5917 18785 5951 18819
rect 8125 18785 8159 18819
rect 14381 18785 14415 18819
rect 16957 18785 16991 18819
rect 19625 18785 19659 18819
rect 20545 18785 20579 18819
rect 6653 18717 6687 18751
rect 6837 18717 6871 18751
rect 7113 18717 7147 18751
rect 7481 18717 7515 18751
rect 7573 18717 7607 18751
rect 7904 18717 7938 18751
rect 15025 18717 15059 18751
rect 15301 18717 15335 18751
rect 15853 18717 15887 18751
rect 16865 18717 16899 18751
rect 17877 18717 17911 18751
rect 19717 18717 19751 18751
rect 20637 18717 20671 18751
rect 33149 18717 33183 18751
rect 6285 18649 6319 18683
rect 7757 18649 7791 18683
rect 15577 18649 15611 18683
rect 15761 18649 15795 18683
rect 17601 18649 17635 18683
rect 17785 18649 17819 18683
rect 34345 18649 34379 18683
rect 15117 18581 15151 18615
rect 15853 18581 15887 18615
rect 4997 18377 5031 18411
rect 5457 18377 5491 18411
rect 6009 18377 6043 18411
rect 14473 18377 14507 18411
rect 15209 18377 15243 18411
rect 15945 18377 15979 18411
rect 17877 18377 17911 18411
rect 8309 18309 8343 18343
rect 10057 18309 10091 18343
rect 13093 18309 13127 18343
rect 14105 18309 14139 18343
rect 16221 18309 16255 18343
rect 4905 18241 4939 18275
rect 6929 18241 6963 18275
rect 7481 18241 7515 18275
rect 8953 18241 8987 18275
rect 9505 18241 9539 18275
rect 9689 18241 9723 18275
rect 10609 18241 10643 18275
rect 11345 18241 11379 18275
rect 12633 18241 12667 18275
rect 12817 18241 12851 18275
rect 13185 18241 13219 18275
rect 13553 18241 13587 18275
rect 14013 18241 14047 18275
rect 14289 18241 14323 18275
rect 14565 18241 14599 18275
rect 14749 18241 14783 18275
rect 14841 18241 14875 18275
rect 14933 18241 14967 18275
rect 15301 18241 15335 18275
rect 15485 18241 15519 18275
rect 15577 18241 15611 18275
rect 15669 18241 15703 18275
rect 17049 18241 17083 18275
rect 17509 18241 17543 18275
rect 17693 18241 17727 18275
rect 9045 18173 9079 18207
rect 10701 18173 10735 18207
rect 13461 18173 13495 18207
rect 16957 18173 16991 18207
rect 9321 18105 9355 18139
rect 9965 18105 9999 18139
rect 17417 18105 17451 18139
rect 13921 18037 13955 18071
rect 6193 17833 6227 17867
rect 10609 17833 10643 17867
rect 10977 17833 11011 17867
rect 14657 17833 14691 17867
rect 18705 17833 18739 17867
rect 20085 17833 20119 17867
rect 20821 17833 20855 17867
rect 23213 17833 23247 17867
rect 24133 17833 24167 17867
rect 9873 17765 9907 17799
rect 10333 17765 10367 17799
rect 12541 17765 12575 17799
rect 15853 17765 15887 17799
rect 18429 17765 18463 17799
rect 18613 17765 18647 17799
rect 23581 17765 23615 17799
rect 3893 17697 3927 17731
rect 10517 17697 10551 17731
rect 11805 17697 11839 17731
rect 14841 17697 14875 17731
rect 15393 17697 15427 17731
rect 18797 17697 18831 17731
rect 18981 17697 19015 17731
rect 21097 17697 21131 17731
rect 21189 17697 21223 17731
rect 22845 17697 22879 17731
rect 23121 17697 23155 17731
rect 24685 17697 24719 17731
rect 1409 17629 1443 17663
rect 7021 17629 7055 17663
rect 7757 17629 7791 17663
rect 9689 17629 9723 17663
rect 9873 17629 9907 17663
rect 10333 17629 10367 17663
rect 10885 17629 10919 17663
rect 10977 17629 11011 17663
rect 11161 17629 11195 17663
rect 11345 17629 11379 17663
rect 11621 17629 11655 17663
rect 12173 17629 12207 17663
rect 12265 17629 12299 17663
rect 14657 17629 14691 17663
rect 15025 17629 15059 17663
rect 15485 17629 15519 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 18521 17629 18555 17663
rect 18889 17629 18923 17663
rect 19073 17629 19107 17663
rect 20269 17629 20303 17663
rect 20361 17629 20395 17663
rect 20453 17629 20487 17663
rect 20610 17629 20644 17663
rect 20729 17629 20763 17663
rect 21005 17629 21039 17663
rect 21281 17629 21315 17663
rect 22753 17629 22787 17663
rect 23397 17629 23431 17663
rect 23673 17629 23707 17663
rect 24409 17629 24443 17663
rect 4169 17561 4203 17595
rect 5917 17561 5951 17595
rect 8953 17561 8987 17595
rect 9137 17561 9171 17595
rect 9505 17561 9539 17595
rect 9965 17561 9999 17595
rect 10609 17561 10643 17595
rect 11897 17561 11931 17595
rect 12081 17561 12115 17595
rect 12541 17561 12575 17595
rect 1593 17493 1627 17527
rect 9229 17493 9263 17527
rect 9321 17493 9355 17527
rect 10793 17493 10827 17527
rect 11437 17493 11471 17527
rect 12173 17493 12207 17527
rect 12357 17493 12391 17527
rect 14473 17493 14507 17527
rect 14933 17493 14967 17527
rect 26157 17493 26191 17527
rect 4997 17289 5031 17323
rect 5457 17289 5491 17323
rect 6009 17289 6043 17323
rect 9689 17289 9723 17323
rect 9873 17289 9907 17323
rect 14841 17289 14875 17323
rect 15117 17289 15151 17323
rect 21465 17289 21499 17323
rect 22017 17289 22051 17323
rect 23121 17289 23155 17323
rect 24869 17289 24903 17323
rect 25329 17289 25363 17323
rect 8033 17221 8067 17255
rect 9137 17221 9171 17255
rect 12265 17221 12299 17255
rect 12481 17221 12515 17255
rect 21281 17221 21315 17255
rect 4905 17153 4939 17187
rect 8769 17153 8803 17187
rect 8861 17153 8895 17187
rect 9045 17153 9079 17187
rect 9229 17153 9263 17187
rect 9505 17153 9539 17187
rect 9597 17153 9631 17187
rect 9873 17153 9907 17187
rect 13185 17153 13219 17187
rect 13369 17153 13403 17187
rect 13645 17153 13679 17187
rect 15025 17153 15059 17187
rect 15209 17153 15243 17187
rect 17969 17153 18003 17187
rect 18613 17153 18647 17187
rect 20729 17153 20763 17187
rect 20821 17153 20855 17187
rect 21005 17153 21039 17187
rect 21097 17153 21131 17187
rect 21373 17153 21407 17187
rect 21833 17153 21867 17187
rect 22017 17153 22051 17187
rect 24777 17153 24811 17187
rect 8401 17085 8435 17119
rect 13553 17085 13587 17119
rect 18061 17085 18095 17119
rect 18337 17085 18371 17119
rect 18521 17085 18555 17119
rect 9413 17017 9447 17051
rect 12633 17017 12667 17051
rect 14565 17017 14599 17051
rect 8493 16949 8527 16983
rect 8622 16949 8656 16983
rect 12449 16949 12483 16983
rect 13737 16949 13771 16983
rect 18889 16949 18923 16983
rect 10149 16745 10183 16779
rect 10333 16745 10367 16779
rect 12633 16745 12667 16779
rect 13461 16745 13495 16779
rect 13737 16745 13771 16779
rect 14289 16745 14323 16779
rect 14841 16745 14875 16779
rect 15669 16745 15703 16779
rect 21189 16745 21223 16779
rect 8033 16677 8067 16711
rect 14197 16677 14231 16711
rect 16497 16677 16531 16711
rect 17325 16677 17359 16711
rect 3893 16609 3927 16643
rect 4169 16609 4203 16643
rect 8953 16609 8987 16643
rect 9965 16609 9999 16643
rect 12541 16609 12575 16643
rect 13921 16609 13955 16643
rect 16681 16609 16715 16643
rect 16865 16609 16899 16643
rect 18613 16609 18647 16643
rect 21097 16609 21131 16643
rect 6377 16541 6411 16575
rect 6837 16541 6871 16575
rect 9321 16541 9355 16575
rect 9413 16541 9447 16575
rect 10615 16541 10649 16575
rect 10787 16541 10821 16575
rect 12357 16541 12391 16575
rect 12633 16541 12667 16575
rect 13645 16541 13679 16575
rect 14105 16541 14139 16575
rect 14381 16541 14415 16575
rect 14565 16541 14599 16575
rect 14933 16541 14967 16575
rect 15117 16541 15151 16575
rect 15853 16541 15887 16575
rect 16037 16541 16071 16575
rect 16129 16541 16163 16575
rect 16957 16541 16991 16575
rect 18705 16541 18739 16575
rect 18797 16541 18831 16575
rect 18889 16541 18923 16575
rect 19533 16541 19567 16575
rect 19625 16541 19659 16575
rect 19809 16541 19843 16575
rect 20729 16541 20763 16575
rect 20821 16541 20855 16575
rect 21005 16541 21039 16575
rect 33149 16541 33183 16575
rect 5917 16473 5951 16507
rect 9045 16473 9079 16507
rect 10317 16473 10351 16507
rect 10517 16473 10551 16507
rect 13921 16473 13955 16507
rect 16221 16473 16255 16507
rect 19257 16473 19291 16507
rect 34345 16473 34379 16507
rect 9597 16405 9631 16439
rect 10701 16405 10735 16439
rect 12817 16405 12851 16439
rect 14657 16405 14691 16439
rect 19073 16405 19107 16439
rect 19441 16405 19475 16439
rect 4537 16201 4571 16235
rect 9229 16201 9263 16235
rect 14473 16201 14507 16235
rect 16405 16201 16439 16235
rect 21189 16201 21223 16235
rect 23121 16201 23155 16235
rect 23765 16201 23799 16235
rect 25605 16201 25639 16235
rect 4353 16133 4387 16167
rect 4813 16133 4847 16167
rect 8585 16133 8619 16167
rect 9321 16133 9355 16167
rect 15669 16133 15703 16167
rect 16221 16133 16255 16167
rect 20821 16133 20855 16167
rect 21005 16133 21039 16167
rect 24133 16133 24167 16167
rect 25789 16133 25823 16167
rect 4445 16065 4479 16099
rect 5273 16065 5307 16099
rect 5457 16065 5491 16099
rect 5825 16065 5859 16099
rect 6009 16065 6043 16099
rect 6193 16065 6227 16099
rect 6837 16065 6871 16099
rect 7113 16065 7147 16099
rect 8677 16065 8711 16099
rect 8953 16065 8987 16099
rect 11529 16065 11563 16099
rect 11713 16065 11747 16099
rect 11805 16065 11839 16099
rect 11989 16065 12023 16099
rect 12633 16065 12667 16099
rect 12817 16065 12851 16099
rect 13093 16065 13127 16099
rect 13369 16065 13403 16099
rect 13553 16065 13587 16099
rect 13737 16065 13771 16099
rect 15301 16065 15335 16099
rect 15485 16065 15519 16099
rect 15577 16065 15611 16099
rect 15761 16065 15795 16099
rect 16497 16065 16531 16099
rect 16681 16065 16715 16099
rect 19901 16065 19935 16099
rect 20085 16065 20119 16099
rect 20177 16065 20211 16099
rect 20361 16065 20395 16099
rect 20453 16065 20487 16099
rect 20545 16065 20579 16099
rect 21465 16065 21499 16099
rect 22017 16065 22051 16099
rect 22477 16065 22511 16099
rect 22661 16065 22695 16099
rect 22937 16065 22971 16099
rect 23397 16065 23431 16099
rect 25881 16065 25915 16099
rect 26157 16065 26191 16099
rect 9045 15997 9079 16031
rect 9689 15997 9723 16031
rect 12265 15997 12299 16031
rect 12909 15997 12943 16031
rect 19993 15997 20027 16031
rect 21281 15997 21315 16031
rect 21649 15997 21683 16031
rect 21925 15997 21959 16031
rect 23305 15997 23339 16031
rect 23857 15997 23891 16031
rect 9781 15929 9815 15963
rect 10241 15929 10275 15963
rect 10609 15929 10643 15963
rect 12173 15929 12207 15963
rect 13001 15929 13035 15963
rect 15393 15929 15427 15963
rect 20729 15929 20763 15963
rect 22385 15929 22419 15963
rect 9873 15861 9907 15895
rect 11529 15861 11563 15895
rect 12081 15861 12115 15895
rect 12541 15861 12575 15895
rect 13277 15861 13311 15895
rect 16221 15861 16255 15895
rect 16773 15861 16807 15895
rect 6193 15657 6227 15691
rect 7021 15657 7055 15691
rect 8493 15657 8527 15691
rect 10149 15657 10183 15691
rect 12357 15657 12391 15691
rect 12817 15657 12851 15691
rect 15301 15657 15335 15691
rect 15577 15657 15611 15691
rect 16221 15657 16255 15691
rect 20913 15657 20947 15691
rect 22385 15657 22419 15691
rect 23765 15657 23799 15691
rect 6653 15589 6687 15623
rect 10609 15589 10643 15623
rect 12909 15589 12943 15623
rect 6745 15521 6779 15555
rect 7757 15521 7791 15555
rect 12541 15521 12575 15555
rect 15209 15521 15243 15555
rect 1409 15453 1443 15487
rect 6377 15453 6411 15487
rect 6524 15453 6558 15487
rect 7941 15453 7975 15487
rect 8217 15453 8251 15487
rect 8309 15453 8343 15487
rect 9505 15453 9539 15487
rect 9689 15453 9723 15487
rect 9781 15453 9815 15487
rect 9873 15453 9907 15487
rect 10425 15453 10459 15487
rect 10793 15453 10827 15487
rect 11069 15453 11103 15487
rect 11437 15453 11471 15487
rect 11897 15453 11931 15487
rect 12265 15453 12299 15487
rect 12909 15453 12943 15487
rect 13093 15453 13127 15487
rect 13185 15453 13219 15487
rect 13369 15453 13403 15487
rect 15393 15453 15427 15487
rect 15669 15453 15703 15487
rect 16129 15453 16163 15487
rect 16313 15453 16347 15487
rect 16681 15453 16715 15487
rect 16865 15453 16899 15487
rect 20821 15453 20855 15487
rect 21005 15453 21039 15487
rect 7849 15385 7883 15419
rect 9321 15385 9355 15419
rect 15117 15385 15151 15419
rect 15853 15385 15887 15419
rect 1593 15317 1627 15351
rect 13277 15317 13311 15351
rect 16037 15317 16071 15351
rect 16773 15317 16807 15351
rect 16865 15113 16899 15147
rect 19717 15113 19751 15147
rect 4353 15045 4387 15079
rect 8493 15045 8527 15079
rect 9689 15045 9723 15079
rect 10241 15045 10275 15079
rect 10425 15045 10459 15079
rect 10793 15045 10827 15079
rect 11253 15045 11287 15079
rect 19533 15045 19567 15079
rect 4077 14977 4111 15011
rect 6653 14977 6687 15011
rect 6837 14977 6871 15011
rect 6930 14999 6964 15033
rect 7022 14983 7056 15017
rect 10609 14977 10643 15011
rect 10885 14977 10919 15011
rect 11069 14977 11103 15011
rect 15393 14977 15427 15011
rect 15577 14977 15611 15011
rect 16681 14977 16715 15011
rect 16865 14977 16899 15011
rect 17325 14977 17359 15011
rect 17969 14977 18003 15011
rect 18889 14977 18923 15011
rect 19349 14977 19383 15011
rect 6101 14909 6135 14943
rect 7665 14909 7699 14943
rect 9321 14909 9355 14943
rect 17233 14909 17267 14943
rect 17877 14909 17911 14943
rect 18981 14909 19015 14943
rect 19257 14909 19291 14943
rect 7297 14841 7331 14875
rect 17693 14841 17727 14875
rect 15577 14773 15611 14807
rect 18245 14773 18279 14807
rect 4905 14569 4939 14603
rect 5181 14569 5215 14603
rect 6837 14569 6871 14603
rect 10057 14569 10091 14603
rect 12725 14569 12759 14603
rect 13369 14569 13403 14603
rect 13829 14569 13863 14603
rect 15393 14569 15427 14603
rect 15945 14569 15979 14603
rect 19533 14569 19567 14603
rect 19993 14569 20027 14603
rect 20637 14569 20671 14603
rect 22293 14569 22327 14603
rect 22569 14569 22603 14603
rect 6193 14501 6227 14535
rect 20729 14501 20763 14535
rect 12081 14433 12115 14467
rect 12817 14433 12851 14467
rect 13461 14433 13495 14467
rect 19625 14433 19659 14467
rect 22661 14433 22695 14467
rect 5089 14365 5123 14399
rect 5549 14365 5583 14399
rect 5825 14365 5859 14399
rect 7113 14365 7147 14399
rect 9965 14365 9999 14399
rect 10517 14365 10551 14399
rect 10885 14365 10919 14399
rect 11161 14365 11195 14399
rect 11345 14365 11379 14399
rect 11437 14365 11471 14399
rect 11529 14365 11563 14399
rect 11989 14365 12023 14399
rect 12265 14365 12299 14399
rect 12357 14365 12391 14399
rect 13001 14365 13035 14399
rect 13645 14365 13679 14399
rect 14657 14365 14691 14399
rect 14841 14365 14875 14399
rect 15025 14365 15059 14399
rect 15301 14365 15335 14399
rect 15820 14365 15854 14399
rect 16221 14365 16255 14399
rect 16405 14365 16439 14399
rect 19257 14365 19291 14399
rect 19717 14365 19751 14399
rect 20177 14365 20211 14399
rect 20453 14365 20487 14399
rect 20729 14365 20763 14399
rect 21005 14365 21039 14399
rect 21097 14365 21131 14399
rect 21281 14365 21315 14399
rect 22385 14365 22419 14399
rect 22477 14365 22511 14399
rect 33149 14365 33183 14399
rect 7021 14297 7055 14331
rect 7573 14297 7607 14331
rect 10701 14297 10735 14331
rect 10793 14297 10827 14331
rect 12725 14297 12759 14331
rect 13369 14297 13403 14331
rect 14933 14297 14967 14331
rect 20840 14297 20874 14331
rect 34345 14297 34379 14331
rect 5457 14229 5491 14263
rect 11069 14229 11103 14263
rect 11713 14229 11747 14263
rect 12541 14229 12575 14263
rect 13185 14229 13219 14263
rect 15209 14229 15243 14263
rect 15761 14229 15795 14263
rect 16405 14229 16439 14263
rect 19349 14229 19383 14263
rect 20269 14229 20303 14263
rect 21281 14229 21315 14263
rect 6561 14025 6595 14059
rect 18889 14025 18923 14059
rect 19073 14025 19107 14059
rect 20269 14025 20303 14059
rect 23673 14025 23707 14059
rect 25513 14025 25547 14059
rect 6101 13957 6135 13991
rect 14565 13957 14599 13991
rect 14657 13957 14691 13991
rect 15209 13957 15243 13991
rect 19717 13957 19751 13991
rect 19901 13957 19935 13991
rect 20545 13957 20579 13991
rect 24041 13957 24075 13991
rect 25697 13957 25731 13991
rect 26065 13957 26099 13991
rect 4077 13889 4111 13923
rect 7481 13889 7515 13923
rect 7849 13889 7883 13923
rect 10609 13889 10643 13923
rect 10793 13889 10827 13923
rect 10891 13889 10925 13923
rect 11069 13889 11103 13923
rect 13185 13889 13219 13923
rect 13461 13889 13495 13923
rect 13645 13889 13679 13923
rect 13921 13889 13955 13923
rect 14289 13889 14323 13923
rect 14381 13889 14415 13923
rect 14749 13889 14783 13923
rect 15301 13889 15335 13923
rect 15577 13889 15611 13923
rect 15669 13889 15703 13923
rect 18797 13889 18831 13923
rect 18981 13889 19015 13923
rect 19809 13889 19843 13923
rect 20085 13889 20119 13923
rect 20361 13889 20395 13923
rect 20821 13889 20855 13923
rect 21005 13889 21039 13923
rect 21189 13889 21223 13923
rect 21281 13889 21315 13923
rect 22017 13889 22051 13923
rect 22753 13889 22787 13923
rect 25789 13889 25823 13923
rect 13093 13821 13127 13855
rect 19257 13821 19291 13855
rect 19349 13821 19383 13855
rect 20729 13821 20763 13855
rect 21925 13821 21959 13855
rect 22385 13821 22419 13855
rect 22661 13821 22695 13855
rect 23121 13821 23155 13855
rect 23765 13821 23799 13855
rect 8677 13753 8711 13787
rect 15393 13753 15427 13787
rect 21005 13753 21039 13787
rect 4340 13685 4374 13719
rect 10701 13685 10735 13719
rect 10977 13685 11011 13719
rect 12357 13685 12391 13719
rect 12909 13685 12943 13719
rect 13921 13685 13955 13719
rect 14933 13685 14967 13719
rect 21465 13685 21499 13719
rect 6377 13481 6411 13515
rect 8401 13481 8435 13515
rect 11805 13481 11839 13515
rect 12725 13481 12759 13515
rect 13185 13481 13219 13515
rect 18981 13481 19015 13515
rect 19625 13481 19659 13515
rect 19993 13481 20027 13515
rect 22385 13481 22419 13515
rect 22661 13481 22695 13515
rect 11713 13413 11747 13447
rect 11897 13413 11931 13447
rect 13001 13413 13035 13447
rect 18245 13413 18279 13447
rect 4077 13345 4111 13379
rect 19257 13345 19291 13379
rect 21649 13345 21683 13379
rect 1409 13277 1443 13311
rect 6101 13277 6135 13311
rect 7297 13277 7331 13311
rect 7941 13277 7975 13311
rect 11989 13277 12023 13311
rect 12173 13277 12207 13311
rect 12449 13277 12483 13311
rect 12725 13277 12759 13311
rect 13093 13277 13127 13311
rect 13369 13277 13403 13311
rect 14105 13277 14139 13311
rect 14289 13277 14323 13311
rect 14381 13277 14415 13311
rect 17601 13277 17635 13311
rect 17785 13277 17819 13311
rect 17969 13277 18003 13311
rect 18797 13277 18831 13311
rect 18981 13277 19015 13311
rect 19441 13277 19475 13311
rect 19717 13277 19751 13311
rect 19993 13277 20027 13311
rect 21557 13277 21591 13311
rect 21741 13277 21775 13311
rect 22109 13277 22143 13311
rect 22201 13277 22235 13311
rect 4353 13209 4387 13243
rect 19901 13209 19935 13243
rect 22385 13209 22419 13243
rect 1593 13141 1627 13175
rect 11437 13141 11471 13175
rect 13645 13141 13679 13175
rect 5181 12937 5215 12971
rect 5549 12937 5583 12971
rect 10425 12937 10459 12971
rect 11253 12937 11287 12971
rect 14657 12937 14691 12971
rect 17325 12937 17359 12971
rect 17969 12937 18003 12971
rect 10333 12869 10367 12903
rect 13001 12869 13035 12903
rect 13093 12869 13127 12903
rect 16037 12869 16071 12903
rect 17141 12869 17175 12903
rect 5089 12801 5123 12835
rect 7297 12801 7331 12835
rect 7849 12801 7883 12835
rect 10241 12801 10275 12835
rect 11529 12801 11563 12835
rect 11713 12801 11747 12835
rect 12081 12801 12115 12835
rect 12265 12801 12299 12835
rect 13369 12801 13403 12835
rect 13645 12801 13679 12835
rect 13829 12801 13863 12835
rect 14565 12801 14599 12835
rect 14841 12801 14875 12835
rect 15669 12801 15703 12835
rect 16221 12801 16255 12835
rect 16313 12801 16347 12835
rect 16681 12801 16715 12835
rect 16865 12801 16899 12835
rect 16957 12801 16991 12835
rect 17233 12801 17267 12835
rect 18245 12801 18279 12835
rect 22293 12801 22327 12835
rect 10793 12733 10827 12767
rect 10885 12733 10919 12767
rect 10977 12733 11011 12767
rect 11069 12733 11103 12767
rect 13553 12733 13587 12767
rect 14105 12733 14139 12767
rect 15025 12733 15059 12767
rect 17693 12733 17727 12767
rect 17785 12733 17819 12767
rect 18337 12733 18371 12767
rect 18613 12733 18647 12767
rect 22201 12733 22235 12767
rect 10057 12665 10091 12699
rect 11621 12665 11655 12699
rect 16129 12665 16163 12699
rect 17233 12665 17267 12699
rect 10609 12597 10643 12631
rect 12265 12597 12299 12631
rect 14013 12597 14047 12631
rect 15761 12597 15795 12631
rect 16681 12597 16715 12631
rect 22661 12597 22695 12631
rect 6469 12393 6503 12427
rect 10793 12393 10827 12427
rect 11345 12393 11379 12427
rect 16313 12393 16347 12427
rect 17049 12393 17083 12427
rect 17877 12393 17911 12427
rect 22477 12393 22511 12427
rect 13921 12325 13955 12359
rect 16865 12325 16899 12359
rect 20637 12325 20671 12359
rect 4169 12257 4203 12291
rect 13645 12257 13679 12291
rect 14289 12257 14323 12291
rect 14841 12257 14875 12291
rect 20177 12257 20211 12291
rect 20821 12257 20855 12291
rect 21281 12257 21315 12291
rect 21741 12257 21775 12291
rect 22201 12257 22235 12291
rect 10701 12189 10735 12223
rect 10885 12189 10919 12223
rect 11437 12189 11471 12223
rect 11621 12189 11655 12223
rect 11713 12189 11747 12223
rect 11805 12189 11839 12223
rect 11989 12189 12023 12223
rect 12265 12189 12299 12223
rect 12541 12189 12575 12223
rect 12725 12189 12759 12223
rect 13553 12189 13587 12223
rect 14105 12189 14139 12223
rect 14565 12189 14599 12223
rect 14933 12189 14967 12223
rect 15945 12189 15979 12223
rect 16589 12189 16623 12223
rect 17417 12189 17451 12223
rect 17509 12189 17543 12223
rect 17693 12189 17727 12223
rect 20269 12189 20303 12223
rect 20729 12189 20763 12223
rect 20913 12189 20947 12223
rect 22293 12189 22327 12223
rect 24409 12189 24443 12223
rect 33149 12189 33183 12223
rect 4445 12121 4479 12155
rect 6193 12121 6227 12155
rect 12633 12121 12667 12155
rect 16313 12121 16347 12155
rect 34345 12121 34379 12155
rect 11621 12053 11655 12087
rect 12173 12053 12207 12087
rect 12357 12053 12391 12087
rect 14473 12053 14507 12087
rect 15761 12053 15795 12087
rect 16497 12053 16531 12087
rect 21833 12053 21867 12087
rect 24501 12053 24535 12087
rect 24961 12053 24995 12087
rect 5273 11849 5307 11883
rect 5641 11849 5675 11883
rect 11805 11849 11839 11883
rect 15669 11849 15703 11883
rect 16313 11849 16347 11883
rect 15301 11781 15335 11815
rect 15501 11781 15535 11815
rect 23673 11781 23707 11815
rect 5181 11713 5215 11747
rect 11989 11713 12023 11747
rect 12173 11713 12207 11747
rect 12449 11713 12483 11747
rect 12633 11713 12667 11747
rect 16129 11713 16163 11747
rect 16313 11713 16347 11747
rect 17325 11713 17359 11747
rect 17509 11713 17543 11747
rect 22109 11713 22143 11747
rect 11897 11645 11931 11679
rect 17417 11645 17451 11679
rect 22017 11645 22051 11679
rect 23397 11645 23431 11679
rect 12357 11577 12391 11611
rect 22477 11577 22511 11611
rect 12633 11509 12667 11543
rect 15485 11509 15519 11543
rect 20637 11509 20671 11543
rect 23305 11509 23339 11543
rect 25145 11509 25179 11543
rect 6561 11305 6595 11339
rect 1593 11237 1627 11271
rect 4537 11169 4571 11203
rect 6285 11169 6319 11203
rect 12357 11169 12391 11203
rect 1409 11101 1443 11135
rect 4261 11101 4295 11135
rect 12265 11101 12299 11135
rect 24501 11101 24535 11135
rect 24961 11101 24995 11135
rect 24593 11033 24627 11067
rect 12633 10965 12667 10999
rect 5273 10761 5307 10795
rect 5641 10761 5675 10795
rect 13737 10693 13771 10727
rect 23765 10693 23799 10727
rect 5181 10625 5215 10659
rect 13461 10557 13495 10591
rect 23489 10557 23523 10591
rect 25237 10489 25271 10523
rect 13277 10421 13311 10455
rect 15209 10421 15243 10455
rect 23305 10421 23339 10455
rect 14473 10217 14507 10251
rect 14381 10013 14415 10047
rect 14841 10013 14875 10047
rect 33149 10013 33183 10047
rect 34345 9945 34379 9979
rect 1593 9129 1627 9163
rect 6285 9129 6319 9163
rect 3985 8993 4019 9027
rect 1409 8925 1443 8959
rect 4261 8857 4295 8891
rect 6009 8857 6043 8891
rect 5089 8585 5123 8619
rect 5549 8585 5583 8619
rect 4997 8449 5031 8483
rect 32965 8041 32999 8075
rect 33149 7837 33183 7871
rect 34345 7769 34379 7803
rect 1409 6749 1443 6783
rect 1593 6613 1627 6647
rect 21649 5729 21683 5763
rect 21373 5661 21407 5695
rect 23397 5661 23431 5695
rect 23673 5661 23707 5695
rect 33149 5661 33183 5695
rect 23305 5593 23339 5627
rect 34345 5593 34379 5627
rect 21189 5525 21223 5559
rect 23121 5525 23155 5559
rect 1593 4777 1627 4811
rect 1409 4573 1443 4607
rect 21097 3553 21131 3587
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 33149 3485 33183 3519
rect 22753 3417 22787 3451
rect 34345 3417 34379 3451
rect 20453 3349 20487 3383
rect 22569 3349 22603 3383
rect 23213 3349 23247 3383
rect 20729 3145 20763 3179
rect 1593 2601 1627 2635
rect 9965 2465 9999 2499
rect 27813 2465 27847 2499
rect 1409 2397 1443 2431
rect 9137 2397 9171 2431
rect 27353 2397 27387 2431
<< metal1 >>
rect 1104 36474 35248 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 35248 36474
rect 1104 36400 35248 36422
rect 934 36116 940 36168
rect 992 36156 998 36168
rect 1397 36159 1455 36165
rect 1397 36156 1409 36159
rect 992 36128 1409 36156
rect 992 36116 998 36128
rect 1397 36125 1409 36128
rect 1443 36125 1455 36159
rect 1397 36119 1455 36125
rect 25590 36116 25596 36168
rect 25648 36156 25654 36168
rect 33137 36159 33195 36165
rect 33137 36156 33149 36159
rect 25648 36128 33149 36156
rect 25648 36116 25654 36128
rect 33137 36125 33149 36128
rect 33183 36125 33195 36159
rect 33137 36119 33195 36125
rect 34330 36048 34336 36100
rect 34388 36048 34394 36100
rect 1581 36023 1639 36029
rect 1581 35989 1593 36023
rect 1627 36020 1639 36023
rect 4614 36020 4620 36032
rect 1627 35992 4620 36020
rect 1627 35989 1639 35992
rect 1581 35983 1639 35989
rect 4614 35980 4620 35992
rect 4672 35980 4678 36032
rect 1104 35930 35236 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 35236 35930
rect 1104 35856 35236 35878
rect 1104 35386 35248 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 35248 35386
rect 1104 35312 35248 35334
rect 934 35028 940 35080
rect 992 35068 998 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 992 35040 1409 35068
rect 992 35028 998 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 3878 34932 3884 34944
rect 1627 34904 3884 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 3878 34892 3884 34904
rect 3936 34892 3942 34944
rect 1104 34842 35236 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 35236 34842
rect 1104 34768 35236 34790
rect 1104 34298 35248 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 35248 34298
rect 1104 34224 35248 34246
rect 23658 33940 23664 33992
rect 23716 33980 23722 33992
rect 33137 33983 33195 33989
rect 33137 33980 33149 33983
rect 23716 33952 33149 33980
rect 23716 33940 23722 33952
rect 33137 33949 33149 33952
rect 33183 33949 33195 33983
rect 33137 33943 33195 33949
rect 34333 33915 34391 33921
rect 34333 33881 34345 33915
rect 34379 33912 34391 33915
rect 34882 33912 34888 33924
rect 34379 33884 34888 33912
rect 34379 33881 34391 33884
rect 34333 33875 34391 33881
rect 34882 33872 34888 33884
rect 34940 33872 34946 33924
rect 1104 33754 35236 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 35236 33754
rect 1104 33680 35236 33702
rect 1104 33210 35248 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 35248 33210
rect 1104 33136 35248 33158
rect 934 32852 940 32904
rect 992 32892 998 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 992 32864 1409 32892
rect 992 32852 998 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32756 1639 32759
rect 4706 32756 4712 32768
rect 1627 32728 4712 32756
rect 1627 32725 1639 32728
rect 1581 32719 1639 32725
rect 4706 32716 4712 32728
rect 4764 32716 4770 32768
rect 1104 32666 35236 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 35236 32666
rect 1104 32592 35236 32614
rect 1104 32122 35248 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 35248 32122
rect 1104 32048 35248 32070
rect 33134 31764 33140 31816
rect 33192 31764 33198 31816
rect 34330 31696 34336 31748
rect 34388 31696 34394 31748
rect 1104 31578 35236 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 35236 31578
rect 1104 31504 35236 31526
rect 1104 31034 35248 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 35248 31034
rect 1104 30960 35248 30982
rect 1394 30676 1400 30728
rect 1452 30676 1458 30728
rect 1581 30583 1639 30589
rect 1581 30549 1593 30583
rect 1627 30580 1639 30583
rect 4798 30580 4804 30592
rect 1627 30552 4804 30580
rect 1627 30549 1639 30552
rect 1581 30543 1639 30549
rect 4798 30540 4804 30552
rect 4856 30540 4862 30592
rect 1104 30490 35236 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 35236 30490
rect 1104 30416 35236 30438
rect 1104 29946 35248 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 35248 29946
rect 1104 29872 35248 29894
rect 33137 29631 33195 29637
rect 33137 29597 33149 29631
rect 33183 29628 33195 29631
rect 33318 29628 33324 29640
rect 33183 29600 33324 29628
rect 33183 29597 33195 29600
rect 33137 29591 33195 29597
rect 33318 29588 33324 29600
rect 33376 29588 33382 29640
rect 34333 29563 34391 29569
rect 34333 29529 34345 29563
rect 34379 29560 34391 29563
rect 34882 29560 34888 29572
rect 34379 29532 34888 29560
rect 34379 29529 34391 29532
rect 34333 29523 34391 29529
rect 34882 29520 34888 29532
rect 34940 29520 34946 29572
rect 1104 29402 35236 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 35236 29402
rect 1104 29328 35236 29350
rect 1104 28858 35248 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 35248 28858
rect 1104 28784 35248 28806
rect 934 28500 940 28552
rect 992 28540 998 28552
rect 1397 28543 1455 28549
rect 1397 28540 1409 28543
rect 992 28512 1409 28540
rect 992 28500 998 28512
rect 1397 28509 1409 28512
rect 1443 28509 1455 28543
rect 1397 28503 1455 28509
rect 1578 28364 1584 28416
rect 1636 28364 1642 28416
rect 23566 28364 23572 28416
rect 23624 28404 23630 28416
rect 23661 28407 23719 28413
rect 23661 28404 23673 28407
rect 23624 28376 23673 28404
rect 23624 28364 23630 28376
rect 23661 28373 23673 28376
rect 23707 28373 23719 28407
rect 23661 28367 23719 28373
rect 1104 28314 35236 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 35236 28314
rect 1104 28240 35236 28262
rect 23566 28200 23572 28212
rect 22066 28172 23572 28200
rect 22066 28132 22094 28172
rect 23566 28160 23572 28172
rect 23624 28160 23630 28212
rect 23658 28160 23664 28212
rect 23716 28160 23722 28212
rect 25590 28160 25596 28212
rect 25648 28160 25654 28212
rect 21928 28104 22094 28132
rect 5905 28067 5963 28073
rect 5905 28033 5917 28067
rect 5951 28064 5963 28067
rect 5994 28064 6000 28076
rect 5951 28036 6000 28064
rect 5951 28033 5963 28036
rect 5905 28027 5963 28033
rect 5994 28024 6000 28036
rect 6052 28064 6058 28076
rect 21928 28073 21956 28104
rect 22922 28092 22928 28144
rect 22980 28092 22986 28144
rect 6549 28067 6607 28073
rect 6549 28064 6561 28067
rect 6052 28036 6561 28064
rect 6052 28024 6058 28036
rect 6549 28033 6561 28036
rect 6595 28033 6607 28067
rect 6549 28027 6607 28033
rect 21637 28067 21695 28073
rect 21637 28033 21649 28067
rect 21683 28064 21695 28067
rect 21913 28067 21971 28073
rect 21913 28064 21925 28067
rect 21683 28036 21925 28064
rect 21683 28033 21695 28036
rect 21637 28027 21695 28033
rect 21913 28033 21925 28036
rect 21959 28033 21971 28067
rect 23584 28064 23612 28160
rect 24854 28092 24860 28144
rect 24912 28092 24918 28144
rect 23842 28064 23848 28076
rect 23584 28036 23848 28064
rect 21913 28027 21971 28033
rect 23842 28024 23848 28036
rect 23900 28024 23906 28076
rect 22186 27956 22192 28008
rect 22244 27956 22250 28008
rect 24121 27999 24179 28005
rect 24121 27996 24133 27999
rect 23952 27968 24133 27996
rect 5902 27820 5908 27872
rect 5960 27860 5966 27872
rect 5997 27863 6055 27869
rect 5997 27860 6009 27863
rect 5960 27832 6009 27860
rect 5960 27820 5966 27832
rect 5997 27829 6009 27832
rect 6043 27829 6055 27863
rect 5997 27823 6055 27829
rect 22646 27820 22652 27872
rect 22704 27860 22710 27872
rect 23952 27860 23980 27968
rect 24121 27965 24133 27968
rect 24167 27965 24179 27999
rect 24121 27959 24179 27965
rect 22704 27832 23980 27860
rect 22704 27820 22710 27832
rect 1104 27770 35248 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 35248 27770
rect 1104 27696 35248 27718
rect 1578 27616 1584 27668
rect 1636 27656 1642 27668
rect 5150 27659 5208 27665
rect 5150 27656 5162 27659
rect 1636 27628 5162 27656
rect 1636 27616 1642 27628
rect 5150 27625 5162 27628
rect 5196 27625 5208 27659
rect 5150 27619 5208 27625
rect 12805 27659 12863 27665
rect 12805 27625 12817 27659
rect 12851 27656 12863 27659
rect 22005 27659 22063 27665
rect 12851 27628 13124 27656
rect 12851 27625 12863 27628
rect 12805 27619 12863 27625
rect 11974 27548 11980 27600
rect 12032 27588 12038 27600
rect 12032 27560 13032 27588
rect 12032 27548 12038 27560
rect 4893 27523 4951 27529
rect 4893 27520 4905 27523
rect 4080 27492 4905 27520
rect 4080 27464 4108 27492
rect 4893 27489 4905 27492
rect 4939 27489 4951 27523
rect 4893 27483 4951 27489
rect 12434 27480 12440 27532
rect 12492 27480 12498 27532
rect 13004 27464 13032 27560
rect 13096 27520 13124 27628
rect 22005 27625 22017 27659
rect 22051 27656 22063 27659
rect 22186 27656 22192 27668
rect 22051 27628 22192 27656
rect 22051 27625 22063 27628
rect 22005 27619 22063 27625
rect 22186 27616 22192 27628
rect 22244 27616 22250 27668
rect 22646 27616 22652 27668
rect 22704 27616 22710 27668
rect 22922 27616 22928 27668
rect 22980 27616 22986 27668
rect 23842 27616 23848 27668
rect 23900 27616 23906 27668
rect 21361 27591 21419 27597
rect 21361 27557 21373 27591
rect 21407 27588 21419 27591
rect 22370 27588 22376 27600
rect 21407 27560 22376 27588
rect 21407 27557 21419 27560
rect 21361 27551 21419 27557
rect 14918 27520 14924 27532
rect 13096 27492 14924 27520
rect 4062 27412 4068 27464
rect 4120 27412 4126 27464
rect 4525 27455 4583 27461
rect 4525 27421 4537 27455
rect 4571 27452 4583 27455
rect 4617 27455 4675 27461
rect 4617 27452 4629 27455
rect 4571 27424 4629 27452
rect 4571 27421 4583 27424
rect 4525 27415 4583 27421
rect 4617 27421 4629 27424
rect 4663 27452 4675 27455
rect 4663 27424 4844 27452
rect 4663 27421 4675 27424
rect 4617 27415 4675 27421
rect 4706 27276 4712 27328
rect 4764 27276 4770 27328
rect 4816 27316 4844 27424
rect 12526 27412 12532 27464
rect 12584 27412 12590 27464
rect 12986 27412 12992 27464
rect 13044 27412 13050 27464
rect 14292 27461 14320 27492
rect 14918 27480 14924 27492
rect 14976 27480 14982 27532
rect 18417 27523 18475 27529
rect 18417 27489 18429 27523
rect 18463 27520 18475 27523
rect 18966 27520 18972 27532
rect 18463 27492 18972 27520
rect 18463 27489 18475 27492
rect 18417 27483 18475 27489
rect 18966 27480 18972 27492
rect 19024 27520 19030 27532
rect 19337 27523 19395 27529
rect 19337 27520 19349 27523
rect 19024 27492 19349 27520
rect 19024 27480 19030 27492
rect 19337 27489 19349 27492
rect 19383 27489 19395 27523
rect 19337 27483 19395 27489
rect 19797 27523 19855 27529
rect 19797 27489 19809 27523
rect 19843 27520 19855 27523
rect 19843 27492 21588 27520
rect 19843 27489 19855 27492
rect 19797 27483 19855 27489
rect 13173 27455 13231 27461
rect 13173 27452 13185 27455
rect 13096 27424 13185 27452
rect 5902 27344 5908 27396
rect 5960 27344 5966 27396
rect 6917 27387 6975 27393
rect 6917 27353 6929 27387
rect 6963 27384 6975 27387
rect 7006 27384 7012 27396
rect 6963 27356 7012 27384
rect 6963 27353 6975 27356
rect 6917 27347 6975 27353
rect 7006 27344 7012 27356
rect 7064 27344 7070 27396
rect 12406 27356 13032 27384
rect 5994 27316 6000 27328
rect 4816 27288 6000 27316
rect 5994 27276 6000 27288
rect 6052 27276 6058 27328
rect 6546 27276 6552 27328
rect 6604 27316 6610 27328
rect 7193 27319 7251 27325
rect 7193 27316 7205 27319
rect 6604 27288 7205 27316
rect 6604 27276 6610 27288
rect 7193 27285 7205 27288
rect 7239 27285 7251 27319
rect 7193 27279 7251 27285
rect 11882 27276 11888 27328
rect 11940 27316 11946 27328
rect 12406 27316 12434 27356
rect 13004 27325 13032 27356
rect 13096 27328 13124 27424
rect 13173 27421 13185 27424
rect 13219 27421 13231 27455
rect 13173 27415 13231 27421
rect 14093 27455 14151 27461
rect 14093 27421 14105 27455
rect 14139 27421 14151 27455
rect 14093 27415 14151 27421
rect 14277 27455 14335 27461
rect 14277 27421 14289 27455
rect 14323 27421 14335 27455
rect 14277 27415 14335 27421
rect 14645 27455 14703 27461
rect 14645 27421 14657 27455
rect 14691 27421 14703 27455
rect 14645 27415 14703 27421
rect 11940 27288 12434 27316
rect 12989 27319 13047 27325
rect 11940 27276 11946 27288
rect 12989 27285 13001 27319
rect 13035 27285 13047 27319
rect 12989 27279 13047 27285
rect 13078 27276 13084 27328
rect 13136 27276 13142 27328
rect 14108 27316 14136 27415
rect 14185 27387 14243 27393
rect 14185 27353 14197 27387
rect 14231 27384 14243 27387
rect 14458 27384 14464 27396
rect 14231 27356 14464 27384
rect 14231 27353 14243 27356
rect 14185 27347 14243 27353
rect 14458 27344 14464 27356
rect 14516 27384 14522 27396
rect 14660 27384 14688 27415
rect 14826 27412 14832 27464
rect 14884 27412 14890 27464
rect 18138 27412 18144 27464
rect 18196 27452 18202 27464
rect 18325 27455 18383 27461
rect 18325 27452 18337 27455
rect 18196 27424 18337 27452
rect 18196 27412 18202 27424
rect 18325 27421 18337 27424
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18509 27455 18567 27461
rect 18509 27421 18521 27455
rect 18555 27421 18567 27455
rect 18509 27415 18567 27421
rect 14516 27356 14688 27384
rect 14516 27344 14522 27356
rect 18524 27328 18552 27415
rect 19242 27412 19248 27464
rect 19300 27452 19306 27464
rect 21560 27461 21588 27492
rect 21744 27461 21772 27560
rect 22370 27548 22376 27560
rect 22428 27548 22434 27600
rect 22940 27588 22968 27616
rect 23017 27591 23075 27597
rect 23017 27588 23029 27591
rect 22940 27560 23029 27588
rect 23017 27557 23029 27560
rect 23063 27557 23075 27591
rect 23017 27551 23075 27557
rect 23860 27520 23888 27616
rect 24118 27520 24124 27532
rect 23860 27492 24124 27520
rect 24118 27480 24124 27492
rect 24176 27520 24182 27532
rect 24397 27523 24455 27529
rect 24397 27520 24409 27523
rect 24176 27492 24409 27520
rect 24176 27480 24182 27492
rect 24397 27489 24409 27492
rect 24443 27489 24455 27523
rect 24397 27483 24455 27489
rect 22087 27465 22145 27471
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19300 27424 19441 27452
rect 19300 27412 19306 27424
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 21453 27455 21511 27461
rect 21453 27421 21465 27455
rect 21499 27421 21511 27455
rect 21453 27415 21511 27421
rect 21545 27455 21603 27461
rect 21545 27421 21557 27455
rect 21591 27421 21603 27455
rect 21545 27415 21603 27421
rect 21729 27455 21787 27461
rect 21729 27421 21741 27455
rect 21775 27421 21787 27455
rect 21729 27415 21787 27421
rect 21468 27384 21496 27415
rect 21818 27412 21824 27464
rect 21876 27412 21882 27464
rect 22087 27462 22099 27465
rect 22020 27434 22099 27462
rect 22020 27396 22048 27434
rect 22087 27431 22099 27434
rect 22133 27431 22145 27465
rect 22087 27425 22145 27431
rect 22186 27412 22192 27464
rect 22244 27412 22250 27464
rect 22370 27412 22376 27464
rect 22428 27412 22434 27464
rect 22465 27455 22523 27461
rect 22465 27421 22477 27455
rect 22511 27421 22523 27455
rect 22465 27415 22523 27421
rect 22925 27455 22983 27461
rect 22925 27421 22937 27455
rect 22971 27452 22983 27455
rect 24029 27455 24087 27461
rect 22971 27424 23520 27452
rect 22971 27421 22983 27424
rect 22925 27415 22983 27421
rect 22002 27384 22008 27396
rect 21468 27356 22008 27384
rect 22002 27344 22008 27356
rect 22060 27344 22066 27396
rect 22480 27384 22508 27415
rect 23492 27393 23520 27424
rect 24029 27421 24041 27455
rect 24075 27421 24087 27455
rect 24029 27415 24087 27421
rect 22296 27356 22508 27384
rect 23477 27387 23535 27393
rect 22296 27328 22324 27356
rect 23477 27353 23489 27387
rect 23523 27384 23535 27387
rect 24044 27384 24072 27415
rect 33226 27412 33232 27464
rect 33284 27412 33290 27464
rect 23523 27356 24072 27384
rect 23523 27353 23535 27356
rect 23477 27347 23535 27353
rect 24044 27328 24072 27356
rect 24670 27344 24676 27396
rect 24728 27344 24734 27396
rect 25406 27344 25412 27396
rect 25464 27344 25470 27396
rect 34333 27387 34391 27393
rect 34333 27353 34345 27387
rect 34379 27384 34391 27387
rect 34882 27384 34888 27396
rect 34379 27356 34888 27384
rect 34379 27353 34391 27356
rect 34333 27347 34391 27353
rect 34882 27344 34888 27356
rect 34940 27344 34946 27396
rect 14550 27316 14556 27328
rect 14108 27288 14556 27316
rect 14550 27276 14556 27288
rect 14608 27276 14614 27328
rect 14737 27319 14795 27325
rect 14737 27285 14749 27319
rect 14783 27316 14795 27319
rect 17126 27316 17132 27328
rect 14783 27288 17132 27316
rect 14783 27285 14795 27288
rect 14737 27279 14795 27285
rect 17126 27276 17132 27288
rect 17184 27316 17190 27328
rect 17678 27316 17684 27328
rect 17184 27288 17684 27316
rect 17184 27276 17190 27288
rect 17678 27276 17684 27288
rect 17736 27276 17742 27328
rect 18506 27276 18512 27328
rect 18564 27276 18570 27328
rect 19150 27276 19156 27328
rect 19208 27316 19214 27328
rect 22186 27316 22192 27328
rect 19208 27288 22192 27316
rect 19208 27276 19214 27288
rect 22186 27276 22192 27288
rect 22244 27276 22250 27328
rect 22278 27276 22284 27328
rect 22336 27276 22342 27328
rect 24026 27276 24032 27328
rect 24084 27276 24090 27328
rect 24121 27319 24179 27325
rect 24121 27285 24133 27319
rect 24167 27316 24179 27319
rect 24854 27316 24860 27328
rect 24167 27288 24860 27316
rect 24167 27285 24179 27288
rect 24121 27279 24179 27285
rect 24854 27276 24860 27288
rect 24912 27276 24918 27328
rect 26145 27319 26203 27325
rect 26145 27285 26157 27319
rect 26191 27316 26203 27319
rect 33134 27316 33140 27328
rect 26191 27288 33140 27316
rect 26191 27285 26203 27288
rect 26145 27279 26203 27285
rect 33134 27276 33140 27288
rect 33192 27276 33198 27328
rect 1104 27226 35236 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 35236 27226
rect 1104 27152 35236 27174
rect 12069 27115 12127 27121
rect 12069 27081 12081 27115
rect 12115 27112 12127 27115
rect 12526 27112 12532 27124
rect 12115 27084 12532 27112
rect 12115 27081 12127 27084
rect 12069 27075 12127 27081
rect 12526 27072 12532 27084
rect 12584 27072 12590 27124
rect 12986 27112 12992 27124
rect 12820 27084 12992 27112
rect 4062 27044 4068 27056
rect 3896 27016 4068 27044
rect 3896 26985 3924 27016
rect 4062 27004 4068 27016
rect 4120 27004 4126 27056
rect 4706 27004 4712 27056
rect 4764 27004 4770 27056
rect 12820 27053 12848 27084
rect 12986 27072 12992 27084
rect 13044 27072 13050 27124
rect 14458 27072 14464 27124
rect 14516 27072 14522 27124
rect 14826 27072 14832 27124
rect 14884 27112 14890 27124
rect 14921 27115 14979 27121
rect 14921 27112 14933 27115
rect 14884 27084 14933 27112
rect 14884 27072 14890 27084
rect 14921 27081 14933 27084
rect 14967 27081 14979 27115
rect 14921 27075 14979 27081
rect 16301 27115 16359 27121
rect 16301 27081 16313 27115
rect 16347 27112 16359 27115
rect 16347 27084 17448 27112
rect 16347 27081 16359 27084
rect 16301 27075 16359 27081
rect 12805 27047 12863 27053
rect 12084 27016 12480 27044
rect 3881 26979 3939 26985
rect 3881 26945 3893 26979
rect 3927 26945 3939 26979
rect 3881 26939 3939 26945
rect 11882 26936 11888 26988
rect 11940 26936 11946 26988
rect 12084 26985 12112 27016
rect 12069 26979 12127 26985
rect 12069 26945 12081 26979
rect 12115 26945 12127 26979
rect 12069 26939 12127 26945
rect 12345 26979 12403 26985
rect 12345 26945 12357 26979
rect 12391 26945 12403 26979
rect 12345 26939 12403 26945
rect 4157 26911 4215 26917
rect 4157 26877 4169 26911
rect 4203 26908 4215 26911
rect 4798 26908 4804 26920
rect 4203 26880 4804 26908
rect 4203 26877 4215 26880
rect 4157 26871 4215 26877
rect 4798 26868 4804 26880
rect 4856 26868 4862 26920
rect 5902 26868 5908 26920
rect 5960 26868 5966 26920
rect 11974 26868 11980 26920
rect 12032 26908 12038 26920
rect 12161 26911 12219 26917
rect 12161 26908 12173 26911
rect 12032 26880 12173 26908
rect 12032 26868 12038 26880
rect 12161 26877 12173 26880
rect 12207 26877 12219 26911
rect 12360 26908 12388 26939
rect 12161 26871 12219 26877
rect 12268 26880 12388 26908
rect 12452 26908 12480 27016
rect 12805 27013 12817 27047
rect 12851 27013 12863 27047
rect 13357 27047 13415 27053
rect 13357 27044 13369 27047
rect 12805 27007 12863 27013
rect 12926 27016 13369 27044
rect 12529 26979 12587 26985
rect 12529 26945 12541 26979
rect 12575 26976 12587 26979
rect 12926 26976 12954 27016
rect 13357 27013 13369 27016
rect 13403 27013 13415 27047
rect 13357 27007 13415 27013
rect 12575 26948 12954 26976
rect 12575 26945 12587 26948
rect 12529 26939 12587 26945
rect 12986 26936 12992 26988
rect 13044 26936 13050 26988
rect 13081 26979 13139 26985
rect 13081 26945 13093 26979
rect 13127 26945 13139 26979
rect 13081 26939 13139 26945
rect 12621 26911 12679 26917
rect 12621 26908 12633 26911
rect 12452 26880 12633 26908
rect 6546 26732 6552 26784
rect 6604 26732 6610 26784
rect 12268 26772 12296 26880
rect 12621 26877 12633 26880
rect 12667 26908 12679 26911
rect 13096 26908 13124 26939
rect 13170 26936 13176 26988
rect 13228 26936 13234 26988
rect 14001 26979 14059 26985
rect 14001 26976 14013 26979
rect 13372 26948 14013 26976
rect 12667 26880 13124 26908
rect 12667 26877 12679 26880
rect 12621 26871 12679 26877
rect 13372 26849 13400 26948
rect 14001 26945 14013 26948
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14093 26979 14151 26985
rect 14093 26945 14105 26979
rect 14139 26976 14151 26979
rect 14182 26976 14188 26988
rect 14139 26948 14188 26976
rect 14139 26945 14151 26948
rect 14093 26939 14151 26945
rect 13357 26843 13415 26849
rect 13357 26809 13369 26843
rect 13403 26809 13415 26843
rect 14016 26840 14044 26939
rect 14182 26936 14188 26948
rect 14240 26976 14246 26988
rect 14369 26979 14427 26985
rect 14369 26976 14381 26979
rect 14240 26948 14381 26976
rect 14240 26936 14246 26948
rect 14369 26945 14381 26948
rect 14415 26945 14427 26979
rect 14369 26939 14427 26945
rect 14476 26976 14504 27072
rect 14844 27016 15608 27044
rect 14844 26985 14872 27016
rect 15580 26988 15608 27016
rect 16022 27004 16028 27056
rect 16080 27044 16086 27056
rect 16669 27047 16727 27053
rect 16669 27044 16681 27047
rect 16080 27016 16681 27044
rect 16080 27004 16086 27016
rect 16669 27013 16681 27016
rect 16715 27013 16727 27047
rect 16669 27007 16727 27013
rect 16758 27004 16764 27056
rect 16816 27044 16822 27056
rect 16869 27047 16927 27053
rect 16869 27044 16881 27047
rect 16816 27016 16881 27044
rect 16816 27004 16822 27016
rect 16869 27013 16881 27016
rect 16915 27013 16927 27047
rect 16869 27007 16927 27013
rect 14645 26979 14703 26985
rect 14645 26976 14657 26979
rect 14476 26948 14657 26976
rect 14277 26911 14335 26917
rect 14277 26877 14289 26911
rect 14323 26908 14335 26911
rect 14476 26908 14504 26948
rect 14645 26945 14657 26948
rect 14691 26945 14703 26979
rect 14645 26939 14703 26945
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 14918 26936 14924 26988
rect 14976 26976 14982 26988
rect 15105 26979 15163 26985
rect 15105 26976 15117 26979
rect 14976 26948 15117 26976
rect 14976 26936 14982 26948
rect 15105 26945 15117 26948
rect 15151 26945 15163 26979
rect 15105 26939 15163 26945
rect 15381 26979 15439 26985
rect 15381 26945 15393 26979
rect 15427 26945 15439 26979
rect 15381 26939 15439 26945
rect 14323 26880 14504 26908
rect 14323 26877 14335 26880
rect 14277 26871 14335 26877
rect 14550 26868 14556 26920
rect 14608 26908 14614 26920
rect 15289 26911 15347 26917
rect 15289 26908 15301 26911
rect 14608 26880 15301 26908
rect 14608 26868 14614 26880
rect 15289 26877 15301 26880
rect 15335 26877 15347 26911
rect 15289 26871 15347 26877
rect 14461 26843 14519 26849
rect 14461 26840 14473 26843
rect 14016 26812 14473 26840
rect 13357 26803 13415 26809
rect 14461 26809 14473 26812
rect 14507 26809 14519 26843
rect 15396 26840 15424 26939
rect 15562 26936 15568 26988
rect 15620 26936 15626 26988
rect 15930 26936 15936 26988
rect 15988 26936 15994 26988
rect 17420 26985 17448 27084
rect 17770 27072 17776 27124
rect 17828 27112 17834 27124
rect 17828 27084 18460 27112
rect 17828 27072 17834 27084
rect 17586 27004 17592 27056
rect 17644 27044 17650 27056
rect 18432 27053 18460 27084
rect 19150 27072 19156 27124
rect 19208 27072 19214 27124
rect 19242 27072 19248 27124
rect 19300 27072 19306 27124
rect 19429 27115 19487 27121
rect 19429 27081 19441 27115
rect 19475 27112 19487 27115
rect 20162 27112 20168 27124
rect 19475 27084 20168 27112
rect 19475 27081 19487 27084
rect 19429 27075 19487 27081
rect 20162 27072 20168 27084
rect 20220 27112 20226 27124
rect 20220 27084 21588 27112
rect 20220 27072 20226 27084
rect 18201 27047 18259 27053
rect 18201 27044 18213 27047
rect 17644 27016 18213 27044
rect 17644 27004 17650 27016
rect 18201 27013 18213 27016
rect 18247 27013 18259 27047
rect 18201 27007 18259 27013
rect 18417 27047 18475 27053
rect 18417 27013 18429 27047
rect 18463 27013 18475 27047
rect 19260 27044 19288 27072
rect 21453 27047 21511 27053
rect 21453 27044 21465 27047
rect 18417 27007 18475 27013
rect 18892 27016 19288 27044
rect 20640 27016 21465 27044
rect 17405 26979 17463 26985
rect 17405 26945 17417 26979
rect 17451 26976 17463 26979
rect 17773 26979 17831 26985
rect 17773 26976 17785 26979
rect 17451 26948 17785 26976
rect 17451 26945 17463 26948
rect 17405 26939 17463 26945
rect 17773 26945 17785 26948
rect 17819 26945 17831 26979
rect 17773 26939 17831 26945
rect 17957 26979 18015 26985
rect 17957 26945 17969 26979
rect 18003 26976 18015 26979
rect 18506 26976 18512 26988
rect 18003 26948 18512 26976
rect 18003 26945 18015 26948
rect 17957 26939 18015 26945
rect 18506 26936 18512 26948
rect 18564 26976 18570 26988
rect 18601 26979 18659 26985
rect 18601 26976 18613 26979
rect 18564 26948 18613 26976
rect 18564 26936 18570 26948
rect 18601 26945 18613 26948
rect 18647 26945 18659 26979
rect 18601 26939 18659 26945
rect 18690 26936 18696 26988
rect 18748 26936 18754 26988
rect 18892 26985 18920 27016
rect 18877 26979 18935 26985
rect 18877 26945 18889 26979
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 18966 26936 18972 26988
rect 19024 26936 19030 26988
rect 20640 26985 20668 27016
rect 21453 27013 21465 27016
rect 21499 27013 21511 27047
rect 21453 27007 21511 27013
rect 20165 26979 20223 26985
rect 20165 26976 20177 26979
rect 19444 26948 20177 26976
rect 15838 26868 15844 26920
rect 15896 26868 15902 26920
rect 17129 26911 17187 26917
rect 17129 26908 17141 26911
rect 17052 26880 17141 26908
rect 17052 26852 17080 26880
rect 17129 26877 17141 26880
rect 17175 26908 17187 26911
rect 17497 26911 17555 26917
rect 17497 26908 17509 26911
rect 17175 26880 17509 26908
rect 17175 26877 17187 26880
rect 17129 26871 17187 26877
rect 17497 26877 17509 26880
rect 17543 26877 17555 26911
rect 17497 26871 17555 26877
rect 17678 26868 17684 26920
rect 17736 26908 17742 26920
rect 17736 26880 18276 26908
rect 17736 26868 17742 26880
rect 14461 26803 14519 26809
rect 14752 26812 15424 26840
rect 12986 26772 12992 26784
rect 12268 26744 12992 26772
rect 12986 26732 12992 26744
rect 13044 26732 13050 26784
rect 14185 26775 14243 26781
rect 14185 26741 14197 26775
rect 14231 26772 14243 26775
rect 14752 26772 14780 26812
rect 16114 26800 16120 26852
rect 16172 26840 16178 26852
rect 16172 26812 16896 26840
rect 16172 26800 16178 26812
rect 14231 26744 14780 26772
rect 15381 26775 15439 26781
rect 14231 26741 14243 26744
rect 14185 26735 14243 26741
rect 15381 26741 15393 26775
rect 15427 26772 15439 26775
rect 16758 26772 16764 26784
rect 15427 26744 16764 26772
rect 15427 26741 15439 26744
rect 15381 26735 15439 26741
rect 16758 26732 16764 26744
rect 16816 26732 16822 26784
rect 16868 26781 16896 26812
rect 17034 26800 17040 26852
rect 17092 26800 17098 26852
rect 17313 26843 17371 26849
rect 17313 26809 17325 26843
rect 17359 26840 17371 26843
rect 17589 26843 17647 26849
rect 17589 26840 17601 26843
rect 17359 26812 17601 26840
rect 17359 26809 17371 26812
rect 17313 26803 17371 26809
rect 17589 26809 17601 26812
rect 17635 26840 17647 26843
rect 18046 26840 18052 26852
rect 17635 26812 18052 26840
rect 17635 26809 17647 26812
rect 17589 26803 17647 26809
rect 18046 26800 18052 26812
rect 18104 26800 18110 26852
rect 18138 26800 18144 26852
rect 18196 26800 18202 26852
rect 16853 26775 16911 26781
rect 16853 26741 16865 26775
rect 16899 26741 16911 26775
rect 16853 26735 16911 26741
rect 17405 26775 17463 26781
rect 17405 26741 17417 26775
rect 17451 26772 17463 26775
rect 18156 26772 18184 26800
rect 18248 26781 18276 26880
rect 17451 26744 18184 26772
rect 18233 26775 18291 26781
rect 17451 26741 17463 26744
rect 17405 26735 17463 26741
rect 18233 26741 18245 26775
rect 18279 26741 18291 26775
rect 18233 26735 18291 26741
rect 19242 26732 19248 26784
rect 19300 26772 19306 26784
rect 19444 26781 19472 26948
rect 20165 26945 20177 26948
rect 20211 26945 20223 26979
rect 20165 26939 20223 26945
rect 20625 26979 20683 26985
rect 20625 26945 20637 26979
rect 20671 26945 20683 26979
rect 21085 26979 21143 26985
rect 21085 26976 21097 26979
rect 20625 26939 20683 26945
rect 20916 26948 21097 26976
rect 19797 26843 19855 26849
rect 19797 26809 19809 26843
rect 19843 26840 19855 26843
rect 19978 26840 19984 26852
rect 19843 26812 19984 26840
rect 19843 26809 19855 26812
rect 19797 26803 19855 26809
rect 19978 26800 19984 26812
rect 20036 26840 20042 26852
rect 20916 26840 20944 26948
rect 21085 26945 21097 26948
rect 21131 26945 21143 26979
rect 21085 26939 21143 26945
rect 21239 26979 21297 26985
rect 21239 26945 21251 26979
rect 21285 26976 21297 26979
rect 21560 26976 21588 27084
rect 25406 27072 25412 27124
rect 25464 27112 25470 27124
rect 25501 27115 25559 27121
rect 25501 27112 25513 27115
rect 25464 27084 25513 27112
rect 25464 27072 25470 27084
rect 25501 27081 25513 27084
rect 25547 27081 25559 27115
rect 25501 27075 25559 27081
rect 21285 26948 21588 26976
rect 21285 26945 21297 26948
rect 21239 26939 21297 26945
rect 22002 26936 22008 26988
rect 22060 26976 22066 26988
rect 22186 26976 22192 26988
rect 22060 26948 22192 26976
rect 22060 26936 22066 26948
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 24026 26936 24032 26988
rect 24084 26976 24090 26988
rect 24397 26979 24455 26985
rect 24397 26976 24409 26979
rect 24084 26948 24409 26976
rect 24084 26936 24090 26948
rect 24397 26945 24409 26948
rect 24443 26976 24455 26979
rect 25133 26979 25191 26985
rect 25133 26976 25145 26979
rect 24443 26948 25145 26976
rect 24443 26945 24455 26948
rect 24397 26939 24455 26945
rect 25133 26945 25145 26948
rect 25179 26976 25191 26979
rect 25409 26979 25467 26985
rect 25409 26976 25421 26979
rect 25179 26948 25421 26976
rect 25179 26945 25191 26948
rect 25133 26939 25191 26945
rect 25409 26945 25421 26948
rect 25455 26976 25467 26979
rect 25455 26948 26004 26976
rect 25455 26945 25467 26948
rect 25409 26939 25467 26945
rect 20993 26911 21051 26917
rect 20993 26877 21005 26911
rect 21039 26908 21051 26911
rect 21818 26908 21824 26920
rect 21039 26880 21824 26908
rect 21039 26877 21051 26880
rect 20993 26871 21051 26877
rect 21818 26868 21824 26880
rect 21876 26908 21882 26920
rect 21913 26911 21971 26917
rect 21913 26908 21925 26911
rect 21876 26880 21925 26908
rect 21876 26868 21882 26880
rect 21913 26877 21925 26880
rect 21959 26908 21971 26911
rect 22278 26908 22284 26920
rect 21959 26880 22284 26908
rect 21959 26877 21971 26880
rect 21913 26871 21971 26877
rect 22278 26868 22284 26880
rect 22336 26868 22342 26920
rect 22373 26911 22431 26917
rect 22373 26877 22385 26911
rect 22419 26908 22431 26911
rect 24670 26908 24676 26920
rect 22419 26880 24676 26908
rect 22419 26877 22431 26880
rect 22373 26871 22431 26877
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 20036 26812 20944 26840
rect 20036 26800 20042 26812
rect 25976 26784 26004 26948
rect 19429 26775 19487 26781
rect 19429 26772 19441 26775
rect 19300 26744 19441 26772
rect 19300 26732 19306 26744
rect 19429 26741 19441 26744
rect 19475 26741 19487 26775
rect 19429 26735 19487 26741
rect 22094 26732 22100 26784
rect 22152 26772 22158 26784
rect 22370 26772 22376 26784
rect 22152 26744 22376 26772
rect 22152 26732 22158 26744
rect 22370 26732 22376 26744
rect 22428 26772 22434 26784
rect 22649 26775 22707 26781
rect 22649 26772 22661 26775
rect 22428 26744 22661 26772
rect 22428 26732 22434 26744
rect 22649 26741 22661 26744
rect 22695 26741 22707 26775
rect 22649 26735 22707 26741
rect 25222 26732 25228 26784
rect 25280 26732 25286 26784
rect 25958 26732 25964 26784
rect 26016 26772 26022 26784
rect 26237 26775 26295 26781
rect 26237 26772 26249 26775
rect 26016 26744 26249 26772
rect 26016 26732 26022 26744
rect 26237 26741 26249 26744
rect 26283 26741 26295 26775
rect 26237 26735 26295 26741
rect 1104 26682 35248 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 35248 26682
rect 1104 26608 35248 26630
rect 5994 26528 6000 26580
rect 6052 26568 6058 26580
rect 6365 26571 6423 26577
rect 6365 26568 6377 26571
rect 6052 26540 6377 26568
rect 6052 26528 6058 26540
rect 6365 26537 6377 26540
rect 6411 26537 6423 26571
rect 6365 26531 6423 26537
rect 12434 26528 12440 26580
rect 12492 26568 12498 26580
rect 12529 26571 12587 26577
rect 12529 26568 12541 26571
rect 12492 26540 12541 26568
rect 12492 26528 12498 26540
rect 12529 26537 12541 26540
rect 12575 26537 12587 26571
rect 12529 26531 12587 26537
rect 13170 26528 13176 26580
rect 13228 26528 13234 26580
rect 14182 26528 14188 26580
rect 14240 26528 14246 26580
rect 15749 26571 15807 26577
rect 15749 26537 15761 26571
rect 15795 26568 15807 26571
rect 18690 26568 18696 26580
rect 15795 26540 18696 26568
rect 15795 26537 15807 26540
rect 15749 26531 15807 26537
rect 18690 26528 18696 26540
rect 18748 26528 18754 26580
rect 24118 26528 24124 26580
rect 24176 26528 24182 26580
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 5261 26367 5319 26373
rect 5261 26333 5273 26367
rect 5307 26364 5319 26367
rect 5442 26364 5448 26376
rect 5307 26336 5448 26364
rect 5307 26333 5319 26336
rect 5261 26327 5319 26333
rect 5442 26324 5448 26336
rect 5500 26364 5506 26376
rect 5721 26367 5779 26373
rect 5721 26364 5733 26367
rect 5500 26336 5733 26364
rect 5500 26324 5506 26336
rect 5721 26333 5733 26336
rect 5767 26364 5779 26367
rect 6012 26364 6040 26528
rect 11793 26435 11851 26441
rect 11793 26401 11805 26435
rect 11839 26432 11851 26435
rect 12161 26435 12219 26441
rect 12161 26432 12173 26435
rect 11839 26404 12173 26432
rect 11839 26401 11851 26404
rect 11793 26395 11851 26401
rect 12161 26401 12173 26404
rect 12207 26401 12219 26435
rect 12161 26395 12219 26401
rect 5767 26336 6040 26364
rect 5767 26333 5779 26336
rect 5721 26327 5779 26333
rect 11698 26324 11704 26376
rect 11756 26324 11762 26376
rect 11885 26367 11943 26373
rect 11885 26364 11897 26367
rect 11808 26336 11897 26364
rect 4614 26296 4620 26308
rect 1596 26268 4620 26296
rect 1596 26237 1624 26268
rect 4614 26256 4620 26268
rect 4672 26256 4678 26308
rect 5353 26299 5411 26305
rect 5353 26265 5365 26299
rect 5399 26296 5411 26299
rect 5534 26296 5540 26308
rect 5399 26268 5540 26296
rect 5399 26265 5411 26268
rect 5353 26259 5411 26265
rect 5534 26256 5540 26268
rect 5592 26256 5598 26308
rect 11808 26240 11836 26336
rect 11885 26333 11897 26336
rect 11931 26333 11943 26367
rect 11885 26327 11943 26333
rect 12069 26367 12127 26373
rect 12069 26333 12081 26367
rect 12115 26333 12127 26367
rect 12069 26327 12127 26333
rect 12084 26296 12112 26327
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12345 26367 12403 26373
rect 12345 26364 12357 26367
rect 12308 26336 12357 26364
rect 12308 26324 12314 26336
rect 12345 26333 12357 26336
rect 12391 26364 12403 26367
rect 13188 26364 13216 26528
rect 15102 26460 15108 26512
rect 15160 26500 15166 26512
rect 15473 26503 15531 26509
rect 15473 26500 15485 26503
rect 15160 26472 15485 26500
rect 15160 26460 15166 26472
rect 15473 26469 15485 26472
rect 15519 26469 15531 26503
rect 15473 26463 15531 26469
rect 15562 26460 15568 26512
rect 15620 26460 15626 26512
rect 16209 26503 16267 26509
rect 16209 26469 16221 26503
rect 16255 26469 16267 26503
rect 16209 26463 16267 26469
rect 15120 26432 15148 26460
rect 14384 26404 15148 26432
rect 15381 26435 15439 26441
rect 12391 26336 13216 26364
rect 12391 26333 12403 26336
rect 12345 26327 12403 26333
rect 14182 26324 14188 26376
rect 14240 26324 14246 26376
rect 14384 26373 14412 26404
rect 15381 26401 15393 26435
rect 15427 26432 15439 26435
rect 15580 26432 15608 26460
rect 15427 26404 15608 26432
rect 15427 26401 15439 26404
rect 15381 26395 15439 26401
rect 14369 26367 14427 26373
rect 14369 26333 14381 26367
rect 14415 26333 14427 26367
rect 14369 26327 14427 26333
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15289 26367 15347 26373
rect 15151 26336 15240 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 15212 26308 15240 26336
rect 15289 26333 15301 26367
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 15565 26367 15623 26373
rect 15565 26333 15577 26367
rect 15611 26333 15623 26367
rect 15565 26327 15623 26333
rect 15933 26367 15991 26373
rect 15933 26333 15945 26367
rect 15979 26333 15991 26367
rect 15933 26327 15991 26333
rect 12802 26296 12808 26308
rect 12084 26268 12808 26296
rect 12802 26256 12808 26268
rect 12860 26256 12866 26308
rect 15194 26256 15200 26308
rect 15252 26256 15258 26308
rect 1581 26231 1639 26237
rect 1581 26197 1593 26231
rect 1627 26228 1639 26231
rect 1627 26200 1661 26228
rect 1627 26197 1639 26200
rect 1581 26191 1639 26197
rect 5626 26188 5632 26240
rect 5684 26188 5690 26240
rect 11790 26188 11796 26240
rect 11848 26188 11854 26240
rect 15013 26231 15071 26237
rect 15013 26197 15025 26231
rect 15059 26228 15071 26231
rect 15304 26228 15332 26327
rect 15378 26228 15384 26240
rect 15059 26200 15384 26228
rect 15059 26197 15071 26200
rect 15013 26191 15071 26197
rect 15378 26188 15384 26200
rect 15436 26188 15442 26240
rect 15580 26228 15608 26327
rect 15948 26296 15976 26327
rect 16022 26324 16028 26376
rect 16080 26324 16086 26376
rect 16224 26364 16252 26463
rect 17034 26460 17040 26512
rect 17092 26460 17098 26512
rect 17126 26460 17132 26512
rect 17184 26460 17190 26512
rect 17497 26503 17555 26509
rect 17497 26469 17509 26503
rect 17543 26469 17555 26503
rect 17497 26463 17555 26469
rect 16945 26367 17003 26373
rect 16945 26364 16957 26367
rect 16224 26336 16957 26364
rect 16945 26333 16957 26336
rect 16991 26333 17003 26367
rect 17052 26364 17080 26460
rect 17144 26432 17172 26460
rect 17144 26404 17264 26432
rect 17236 26373 17264 26404
rect 17129 26367 17187 26373
rect 17129 26364 17141 26367
rect 17052 26336 17141 26364
rect 16945 26327 17003 26333
rect 17129 26333 17141 26336
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17221 26367 17279 26373
rect 17221 26333 17233 26367
rect 17267 26333 17279 26367
rect 17512 26364 17540 26463
rect 18046 26460 18052 26512
rect 18104 26460 18110 26512
rect 22925 26503 22983 26509
rect 22925 26469 22937 26503
rect 22971 26500 22983 26503
rect 23014 26500 23020 26512
rect 22971 26472 23020 26500
rect 22971 26469 22983 26472
rect 22925 26463 22983 26469
rect 23014 26460 23020 26472
rect 23072 26460 23078 26512
rect 18064 26373 18092 26460
rect 22741 26435 22799 26441
rect 22741 26401 22753 26435
rect 22787 26401 22799 26435
rect 24136 26432 24164 26528
rect 24397 26435 24455 26441
rect 24397 26432 24409 26435
rect 24136 26404 24409 26432
rect 22741 26395 22799 26401
rect 24397 26401 24409 26404
rect 24443 26401 24455 26435
rect 24397 26395 24455 26401
rect 26145 26435 26203 26441
rect 26145 26401 26157 26435
rect 26191 26432 26203 26435
rect 33318 26432 33324 26444
rect 26191 26404 33324 26432
rect 26191 26401 26203 26404
rect 26145 26395 26203 26401
rect 17865 26367 17923 26373
rect 17865 26364 17877 26367
rect 17512 26336 17877 26364
rect 17221 26327 17279 26333
rect 17865 26333 17877 26336
rect 17911 26333 17923 26367
rect 17865 26327 17923 26333
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26333 18107 26367
rect 22756 26364 22784 26395
rect 33318 26392 33324 26404
rect 33376 26392 33382 26444
rect 22830 26364 22836 26376
rect 22756 26336 22836 26364
rect 18049 26327 18107 26333
rect 22830 26324 22836 26336
rect 22888 26324 22894 26376
rect 23017 26367 23075 26373
rect 23017 26333 23029 26367
rect 23063 26364 23075 26367
rect 23106 26364 23112 26376
rect 23063 26336 23112 26364
rect 23063 26333 23075 26336
rect 23017 26327 23075 26333
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 16114 26296 16120 26308
rect 15948 26268 16120 26296
rect 16114 26256 16120 26268
rect 16172 26256 16178 26308
rect 16209 26299 16267 26305
rect 16209 26265 16221 26299
rect 16255 26296 16267 26299
rect 16758 26296 16764 26308
rect 16255 26268 16764 26296
rect 16255 26265 16267 26268
rect 16209 26259 16267 26265
rect 16758 26256 16764 26268
rect 16816 26256 16822 26308
rect 17037 26299 17095 26305
rect 17037 26265 17049 26299
rect 17083 26296 17095 26299
rect 17497 26299 17555 26305
rect 17497 26296 17509 26299
rect 17083 26268 17509 26296
rect 17083 26265 17095 26268
rect 17037 26259 17095 26265
rect 17497 26265 17509 26268
rect 17543 26296 17555 26299
rect 17586 26296 17592 26308
rect 17543 26268 17592 26296
rect 17543 26265 17555 26268
rect 17497 26259 17555 26265
rect 17586 26256 17592 26268
rect 17644 26256 17650 26308
rect 17770 26256 17776 26308
rect 17828 26256 17834 26308
rect 17957 26299 18015 26305
rect 17957 26265 17969 26299
rect 18003 26296 18015 26299
rect 19242 26296 19248 26308
rect 18003 26268 19248 26296
rect 18003 26265 18015 26268
rect 17957 26259 18015 26265
rect 19242 26256 19248 26268
rect 19300 26256 19306 26308
rect 22741 26299 22799 26305
rect 22741 26265 22753 26299
rect 22787 26296 22799 26299
rect 23474 26296 23480 26308
rect 22787 26268 23480 26296
rect 22787 26265 22799 26268
rect 22741 26259 22799 26265
rect 23474 26256 23480 26268
rect 23532 26256 23538 26308
rect 24670 26256 24676 26308
rect 24728 26256 24734 26308
rect 25222 26256 25228 26308
rect 25280 26256 25286 26308
rect 17313 26231 17371 26237
rect 17313 26228 17325 26231
rect 15580 26200 17325 26228
rect 17313 26197 17325 26200
rect 17359 26228 17371 26231
rect 17788 26228 17816 26256
rect 17359 26200 17816 26228
rect 17359 26197 17371 26200
rect 17313 26191 17371 26197
rect 1104 26138 35236 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 35236 26138
rect 1104 26064 35236 26086
rect 14001 26027 14059 26033
rect 10704 25996 12434 26024
rect 4522 25916 4528 25968
rect 4580 25916 4586 25968
rect 5534 25916 5540 25968
rect 5592 25916 5598 25968
rect 10704 25900 10732 25996
rect 10965 25959 11023 25965
rect 10965 25925 10977 25959
rect 11011 25956 11023 25959
rect 11609 25959 11667 25965
rect 11609 25956 11621 25959
rect 11011 25928 11621 25956
rect 11011 25925 11023 25928
rect 10965 25919 11023 25925
rect 10686 25848 10692 25900
rect 10744 25848 10750 25900
rect 10778 25848 10784 25900
rect 10836 25848 10842 25900
rect 11164 25897 11192 25928
rect 11609 25925 11621 25928
rect 11655 25956 11667 25959
rect 11698 25956 11704 25968
rect 11655 25928 11704 25956
rect 11655 25925 11667 25928
rect 11609 25919 11667 25925
rect 11698 25916 11704 25928
rect 11756 25916 11762 25968
rect 12406 25956 12434 25996
rect 14001 25993 14013 26027
rect 14047 26024 14059 26027
rect 14182 26024 14188 26036
rect 14047 25996 14188 26024
rect 14047 25993 14059 25996
rect 14001 25987 14059 25993
rect 14182 25984 14188 25996
rect 14240 25984 14246 26036
rect 15473 26027 15531 26033
rect 15473 25993 15485 26027
rect 15519 26024 15531 26027
rect 15930 26024 15936 26036
rect 15519 25996 15936 26024
rect 15519 25993 15531 25996
rect 15473 25987 15531 25993
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 17770 25984 17776 26036
rect 17828 25984 17834 26036
rect 22186 25984 22192 26036
rect 22244 25984 22250 26036
rect 23474 25984 23480 26036
rect 23532 25984 23538 26036
rect 23661 26027 23719 26033
rect 23661 25993 23673 26027
rect 23707 26024 23719 26027
rect 24670 26024 24676 26036
rect 23707 25996 24676 26024
rect 23707 25993 23719 25996
rect 23661 25987 23719 25993
rect 24670 25984 24676 25996
rect 24728 25984 24734 26036
rect 12406 25928 14320 25956
rect 11149 25891 11207 25897
rect 11149 25857 11161 25891
rect 11195 25857 11207 25891
rect 11149 25851 11207 25857
rect 11333 25891 11391 25897
rect 11333 25857 11345 25891
rect 11379 25888 11391 25891
rect 11790 25888 11796 25900
rect 11379 25860 11796 25888
rect 11379 25857 11391 25860
rect 11333 25851 11391 25857
rect 11790 25848 11796 25860
rect 11848 25848 11854 25900
rect 11977 25891 12035 25897
rect 11977 25857 11989 25891
rect 12023 25888 12035 25891
rect 12345 25891 12403 25897
rect 12345 25888 12357 25891
rect 12023 25860 12357 25888
rect 12023 25857 12035 25860
rect 11977 25851 12035 25857
rect 12345 25857 12357 25860
rect 12391 25857 12403 25891
rect 12345 25851 12403 25857
rect 12802 25848 12808 25900
rect 12860 25888 12866 25900
rect 13832 25897 13860 25928
rect 14292 25897 14320 25928
rect 15194 25916 15200 25968
rect 15252 25956 15258 25968
rect 16209 25959 16267 25965
rect 16209 25956 16221 25959
rect 15252 25928 15700 25956
rect 15252 25916 15258 25928
rect 15672 25900 15700 25928
rect 15764 25928 16221 25956
rect 12989 25891 13047 25897
rect 12989 25888 13001 25891
rect 12860 25860 13001 25888
rect 12860 25848 12866 25860
rect 12989 25857 13001 25860
rect 13035 25857 13047 25891
rect 12989 25851 13047 25857
rect 13817 25891 13875 25897
rect 13817 25857 13829 25891
rect 13863 25857 13875 25891
rect 13817 25851 13875 25857
rect 14093 25891 14151 25897
rect 14093 25857 14105 25891
rect 14139 25857 14151 25891
rect 14093 25851 14151 25857
rect 14277 25891 14335 25897
rect 14277 25857 14289 25891
rect 14323 25857 14335 25891
rect 14277 25851 14335 25857
rect 4062 25780 4068 25832
rect 4120 25820 4126 25832
rect 4249 25823 4307 25829
rect 4249 25820 4261 25823
rect 4120 25792 4261 25820
rect 4120 25780 4126 25792
rect 4249 25789 4261 25792
rect 4295 25789 4307 25823
rect 4249 25783 4307 25789
rect 11241 25823 11299 25829
rect 11241 25789 11253 25823
rect 11287 25820 11299 25823
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 11287 25792 12173 25820
rect 11287 25789 11299 25792
rect 11241 25783 11299 25789
rect 12161 25789 12173 25792
rect 12207 25820 12219 25823
rect 12250 25820 12256 25832
rect 12207 25792 12256 25820
rect 12207 25789 12219 25792
rect 12161 25783 12219 25789
rect 12250 25780 12256 25792
rect 12308 25780 12314 25832
rect 12529 25823 12587 25829
rect 12529 25789 12541 25823
rect 12575 25820 12587 25823
rect 12897 25823 12955 25829
rect 12897 25820 12909 25823
rect 12575 25792 12909 25820
rect 12575 25789 12587 25792
rect 12529 25783 12587 25789
rect 12897 25789 12909 25792
rect 12943 25789 12955 25823
rect 13633 25823 13691 25829
rect 13633 25820 13645 25823
rect 12897 25783 12955 25789
rect 13280 25792 13645 25820
rect 5997 25755 6055 25761
rect 5997 25721 6009 25755
rect 6043 25752 6055 25755
rect 6914 25752 6920 25764
rect 6043 25724 6920 25752
rect 6043 25721 6055 25724
rect 5997 25715 6055 25721
rect 6914 25712 6920 25724
rect 6972 25712 6978 25764
rect 13280 25752 13308 25792
rect 13633 25789 13645 25792
rect 13679 25820 13691 25823
rect 14108 25820 14136 25851
rect 15102 25848 15108 25900
rect 15160 25888 15166 25900
rect 15381 25891 15439 25897
rect 15381 25888 15393 25891
rect 15160 25860 15393 25888
rect 15160 25848 15166 25860
rect 15381 25857 15393 25860
rect 15427 25857 15439 25891
rect 15381 25851 15439 25857
rect 15562 25848 15568 25900
rect 15620 25848 15626 25900
rect 15654 25848 15660 25900
rect 15712 25848 15718 25900
rect 15764 25897 15792 25928
rect 16209 25925 16221 25928
rect 16255 25925 16267 25959
rect 16209 25919 16267 25925
rect 15749 25891 15807 25897
rect 15749 25857 15761 25891
rect 15795 25857 15807 25891
rect 15749 25851 15807 25857
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25888 15991 25891
rect 16390 25888 16396 25900
rect 15979 25860 16396 25888
rect 15979 25857 15991 25860
rect 15933 25851 15991 25857
rect 13679 25792 14136 25820
rect 14185 25823 14243 25829
rect 13679 25789 13691 25792
rect 13633 25783 13691 25789
rect 14185 25789 14197 25823
rect 14231 25820 14243 25823
rect 15120 25820 15148 25848
rect 15764 25820 15792 25851
rect 16390 25848 16396 25860
rect 16448 25888 16454 25900
rect 17313 25891 17371 25897
rect 17313 25888 17325 25891
rect 16448 25860 17325 25888
rect 16448 25848 16454 25860
rect 17313 25857 17325 25860
rect 17359 25888 17371 25891
rect 17788 25888 17816 25984
rect 22094 25916 22100 25968
rect 22152 25956 22158 25968
rect 22152 25928 22508 25956
rect 22152 25916 22158 25928
rect 17359 25860 17816 25888
rect 17359 25857 17371 25860
rect 17313 25851 17371 25857
rect 18414 25848 18420 25900
rect 18472 25888 18478 25900
rect 19978 25888 19984 25900
rect 18472 25860 19984 25888
rect 18472 25848 18478 25860
rect 19978 25848 19984 25860
rect 20036 25888 20042 25900
rect 22480 25897 22508 25928
rect 22756 25928 22968 25956
rect 22756 25897 22784 25928
rect 20073 25891 20131 25897
rect 20073 25888 20085 25891
rect 20036 25860 20085 25888
rect 20036 25848 20042 25860
rect 20073 25857 20085 25860
rect 20119 25857 20131 25891
rect 20073 25851 20131 25857
rect 20257 25891 20315 25897
rect 20257 25857 20269 25891
rect 20303 25857 20315 25891
rect 20257 25851 20315 25857
rect 20441 25891 20499 25897
rect 20441 25857 20453 25891
rect 20487 25888 20499 25891
rect 20901 25891 20959 25897
rect 20901 25888 20913 25891
rect 20487 25860 20913 25888
rect 20487 25857 20499 25860
rect 20441 25851 20499 25857
rect 20901 25857 20913 25860
rect 20947 25857 20959 25891
rect 22373 25891 22431 25897
rect 22373 25888 22385 25891
rect 20901 25851 20959 25857
rect 21284 25860 22385 25888
rect 14231 25792 15148 25820
rect 15396 25792 15792 25820
rect 14231 25789 14243 25792
rect 14185 25783 14243 25789
rect 12406 25724 13308 25752
rect 13357 25755 13415 25761
rect 6086 25644 6092 25696
rect 6144 25684 6150 25696
rect 6546 25684 6552 25696
rect 6144 25656 6552 25684
rect 6144 25644 6150 25656
rect 6546 25644 6552 25656
rect 6604 25644 6610 25696
rect 6638 25644 6644 25696
rect 6696 25684 6702 25696
rect 10045 25687 10103 25693
rect 10045 25684 10057 25687
rect 6696 25656 10057 25684
rect 6696 25644 6702 25656
rect 10045 25653 10057 25656
rect 10091 25684 10103 25687
rect 10134 25684 10140 25696
rect 10091 25656 10140 25684
rect 10091 25653 10103 25656
rect 10045 25647 10103 25653
rect 10134 25644 10140 25656
rect 10192 25684 10198 25696
rect 11698 25684 11704 25696
rect 10192 25656 11704 25684
rect 10192 25644 10198 25656
rect 11698 25644 11704 25656
rect 11756 25644 11762 25696
rect 12158 25644 12164 25696
rect 12216 25684 12222 25696
rect 12406 25684 12434 25724
rect 13357 25721 13369 25755
rect 13403 25752 13415 25755
rect 13814 25752 13820 25764
rect 13403 25724 13820 25752
rect 13403 25721 13415 25724
rect 13357 25715 13415 25721
rect 13814 25712 13820 25724
rect 13872 25712 13878 25764
rect 15396 25696 15424 25792
rect 16022 25780 16028 25832
rect 16080 25780 16086 25832
rect 17126 25780 17132 25832
rect 17184 25820 17190 25832
rect 17221 25823 17279 25829
rect 17221 25820 17233 25823
rect 17184 25792 17233 25820
rect 17184 25780 17190 25792
rect 17221 25789 17233 25792
rect 17267 25789 17279 25823
rect 20272 25820 20300 25851
rect 20272 25792 20484 25820
rect 17221 25783 17279 25789
rect 15841 25755 15899 25761
rect 15841 25721 15853 25755
rect 15887 25752 15899 25755
rect 16040 25752 16068 25780
rect 15887 25724 16068 25752
rect 15887 25721 15899 25724
rect 15841 25715 15899 25721
rect 20456 25696 20484 25792
rect 20990 25780 20996 25832
rect 21048 25780 21054 25832
rect 21284 25761 21312 25860
rect 22373 25857 22385 25860
rect 22419 25857 22431 25891
rect 22373 25851 22431 25857
rect 22465 25891 22523 25897
rect 22465 25857 22477 25891
rect 22511 25857 22523 25891
rect 22465 25851 22523 25857
rect 22649 25891 22707 25897
rect 22649 25857 22661 25891
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 22741 25891 22799 25897
rect 22741 25857 22753 25891
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 21269 25755 21327 25761
rect 21269 25721 21281 25755
rect 21315 25721 21327 25755
rect 21269 25715 21327 25721
rect 12216 25656 12434 25684
rect 12216 25644 12222 25656
rect 15378 25644 15384 25696
rect 15436 25644 15442 25696
rect 17681 25687 17739 25693
rect 17681 25653 17693 25687
rect 17727 25684 17739 25687
rect 18230 25684 18236 25696
rect 17727 25656 18236 25684
rect 17727 25653 17739 25656
rect 17681 25647 17739 25653
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 20438 25644 20444 25696
rect 20496 25644 20502 25696
rect 22094 25644 22100 25696
rect 22152 25644 22158 25696
rect 22388 25684 22416 25851
rect 22664 25752 22692 25851
rect 22830 25848 22836 25900
rect 22888 25848 22894 25900
rect 22940 25829 22968 25928
rect 23492 25897 23520 25984
rect 26053 25959 26111 25965
rect 26053 25956 26065 25959
rect 25622 25928 26065 25956
rect 26053 25925 26065 25928
rect 26099 25925 26111 25959
rect 26053 25919 26111 25925
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 23937 25891 23995 25897
rect 23937 25857 23949 25891
rect 23983 25888 23995 25891
rect 24118 25888 24124 25900
rect 23983 25860 24124 25888
rect 23983 25857 23995 25860
rect 23937 25851 23995 25857
rect 24118 25848 24124 25860
rect 24176 25848 24182 25900
rect 25958 25888 25964 25900
rect 25792 25860 25964 25888
rect 22925 25823 22983 25829
rect 22925 25789 22937 25823
rect 22971 25820 22983 25823
rect 23106 25820 23112 25832
rect 22971 25792 23112 25820
rect 22971 25789 22983 25792
rect 22925 25783 22983 25789
rect 23106 25780 23112 25792
rect 23164 25780 23170 25832
rect 23293 25823 23351 25829
rect 23293 25820 23305 25823
rect 23216 25792 23305 25820
rect 23216 25761 23244 25792
rect 23293 25789 23305 25792
rect 23339 25789 23351 25823
rect 23293 25783 23351 25789
rect 24394 25780 24400 25832
rect 24452 25780 24458 25832
rect 23201 25755 23259 25761
rect 22664 25724 23060 25752
rect 23032 25696 23060 25724
rect 23201 25721 23213 25755
rect 23247 25721 23259 25755
rect 23201 25715 23259 25721
rect 22830 25684 22836 25696
rect 22388 25656 22836 25684
rect 22830 25644 22836 25656
rect 22888 25644 22894 25696
rect 23014 25644 23020 25696
rect 23072 25644 23078 25696
rect 25498 25644 25504 25696
rect 25556 25684 25562 25696
rect 25792 25684 25820 25860
rect 25958 25848 25964 25860
rect 26016 25888 26022 25900
rect 26145 25891 26203 25897
rect 26145 25888 26157 25891
rect 26016 25860 26157 25888
rect 26016 25848 26022 25860
rect 26145 25857 26157 25860
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 25869 25823 25927 25829
rect 25869 25789 25881 25823
rect 25915 25820 25927 25823
rect 33226 25820 33232 25832
rect 25915 25792 33232 25820
rect 25915 25789 25927 25792
rect 25869 25783 25927 25789
rect 33226 25780 33232 25792
rect 33284 25780 33290 25832
rect 26421 25687 26479 25693
rect 26421 25684 26433 25687
rect 25556 25656 26433 25684
rect 25556 25644 25562 25656
rect 26421 25653 26433 25656
rect 26467 25653 26479 25687
rect 26421 25647 26479 25653
rect 1104 25594 35248 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 35248 25594
rect 1104 25520 35248 25542
rect 5626 25480 5632 25492
rect 5552 25452 5632 25480
rect 4433 25347 4491 25353
rect 4433 25313 4445 25347
rect 4479 25344 4491 25347
rect 4890 25344 4896 25356
rect 4479 25316 4896 25344
rect 4479 25313 4491 25316
rect 4433 25307 4491 25313
rect 4890 25304 4896 25316
rect 4948 25304 4954 25356
rect 4062 25236 4068 25288
rect 4120 25276 4126 25288
rect 4157 25279 4215 25285
rect 4157 25276 4169 25279
rect 4120 25248 4169 25276
rect 4120 25236 4126 25248
rect 4157 25245 4169 25248
rect 4203 25245 4215 25279
rect 5552 25262 5580 25452
rect 5626 25440 5632 25452
rect 5684 25440 5690 25492
rect 8018 25440 8024 25492
rect 8076 25440 8082 25492
rect 10134 25440 10140 25492
rect 10192 25440 10198 25492
rect 10597 25483 10655 25489
rect 10597 25449 10609 25483
rect 10643 25449 10655 25483
rect 10597 25443 10655 25449
rect 7197 25415 7255 25421
rect 7197 25381 7209 25415
rect 7243 25412 7255 25415
rect 8036 25412 8064 25440
rect 7243 25384 8064 25412
rect 7243 25381 7255 25384
rect 7197 25375 7255 25381
rect 7929 25347 7987 25353
rect 7929 25344 7941 25347
rect 6932 25316 7941 25344
rect 6932 25288 6960 25316
rect 7929 25313 7941 25316
rect 7975 25313 7987 25347
rect 7929 25307 7987 25313
rect 9950 25304 9956 25356
rect 10008 25344 10014 25356
rect 10612 25344 10640 25443
rect 10686 25440 10692 25492
rect 10744 25440 10750 25492
rect 10778 25440 10784 25492
rect 10836 25480 10842 25492
rect 11057 25483 11115 25489
rect 11057 25480 11069 25483
rect 10836 25452 11069 25480
rect 10836 25440 10842 25452
rect 11057 25449 11069 25452
rect 11103 25449 11115 25483
rect 11057 25443 11115 25449
rect 11790 25440 11796 25492
rect 11848 25440 11854 25492
rect 12618 25440 12624 25492
rect 12676 25440 12682 25492
rect 12805 25483 12863 25489
rect 12805 25449 12817 25483
rect 12851 25480 12863 25483
rect 12986 25480 12992 25492
rect 12851 25452 12992 25480
rect 12851 25449 12863 25452
rect 12805 25443 12863 25449
rect 12986 25440 12992 25452
rect 13044 25440 13050 25492
rect 15838 25440 15844 25492
rect 15896 25480 15902 25492
rect 15933 25483 15991 25489
rect 15933 25480 15945 25483
rect 15896 25452 15945 25480
rect 15896 25440 15902 25452
rect 15933 25449 15945 25452
rect 15979 25449 15991 25483
rect 15933 25443 15991 25449
rect 17957 25483 18015 25489
rect 17957 25449 17969 25483
rect 18003 25480 18015 25483
rect 18003 25452 18644 25480
rect 18003 25449 18015 25452
rect 17957 25443 18015 25449
rect 10704 25412 10732 25440
rect 18616 25424 18644 25452
rect 20162 25440 20168 25492
rect 20220 25440 20226 25492
rect 20438 25480 20444 25492
rect 20272 25452 20444 25480
rect 10965 25415 11023 25421
rect 10965 25412 10977 25415
rect 10704 25384 10977 25412
rect 10965 25381 10977 25384
rect 11011 25381 11023 25415
rect 12526 25412 12532 25424
rect 10965 25375 11023 25381
rect 11256 25384 12532 25412
rect 11256 25353 11284 25384
rect 12526 25372 12532 25384
rect 12584 25372 12590 25424
rect 15654 25412 15660 25424
rect 15488 25384 15660 25412
rect 11241 25347 11299 25353
rect 11241 25344 11253 25347
rect 10008 25316 11253 25344
rect 10008 25304 10014 25316
rect 11241 25313 11253 25316
rect 11287 25313 11299 25347
rect 11241 25307 11299 25313
rect 11698 25304 11704 25356
rect 11756 25304 11762 25356
rect 12158 25344 12164 25356
rect 11808 25316 12164 25344
rect 11808 25288 11836 25316
rect 12158 25304 12164 25316
rect 12216 25304 12222 25356
rect 14737 25347 14795 25353
rect 14737 25344 14749 25347
rect 12268 25316 14749 25344
rect 4157 25239 4215 25245
rect 6914 25236 6920 25288
rect 6972 25236 6978 25288
rect 7006 25236 7012 25288
rect 7064 25276 7070 25288
rect 7101 25279 7159 25285
rect 7101 25276 7113 25279
rect 7064 25248 7113 25276
rect 7064 25236 7070 25248
rect 7101 25245 7113 25248
rect 7147 25245 7159 25279
rect 7101 25239 7159 25245
rect 7282 25236 7288 25288
rect 7340 25236 7346 25288
rect 7374 25236 7380 25288
rect 7432 25236 7438 25288
rect 7834 25236 7840 25288
rect 7892 25236 7898 25288
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25245 10655 25279
rect 10597 25239 10655 25245
rect 6178 25168 6184 25220
rect 6236 25168 6242 25220
rect 7926 25168 7932 25220
rect 7984 25208 7990 25220
rect 8113 25211 8171 25217
rect 8113 25208 8125 25211
rect 7984 25180 8125 25208
rect 7984 25168 7990 25180
rect 8113 25177 8125 25180
rect 8159 25177 8171 25211
rect 8113 25171 8171 25177
rect 10134 25168 10140 25220
rect 10192 25208 10198 25220
rect 10321 25211 10379 25217
rect 10321 25208 10333 25211
rect 10192 25180 10333 25208
rect 10192 25168 10198 25180
rect 10321 25177 10333 25180
rect 10367 25177 10379 25211
rect 10321 25171 10379 25177
rect 10612 25208 10640 25239
rect 10778 25236 10784 25288
rect 10836 25236 10842 25288
rect 11333 25279 11391 25285
rect 11333 25245 11345 25279
rect 11379 25245 11391 25279
rect 11333 25239 11391 25245
rect 11146 25208 11152 25220
rect 10612 25180 11152 25208
rect 6086 25100 6092 25152
rect 6144 25140 6150 25152
rect 6457 25143 6515 25149
rect 6457 25140 6469 25143
rect 6144 25112 6469 25140
rect 6144 25100 6150 25112
rect 6457 25109 6469 25112
rect 6503 25109 6515 25143
rect 6457 25103 6515 25109
rect 6917 25143 6975 25149
rect 6917 25109 6929 25143
rect 6963 25140 6975 25143
rect 7466 25140 7472 25152
rect 6963 25112 7472 25140
rect 6963 25109 6975 25112
rect 6917 25103 6975 25109
rect 7466 25100 7472 25112
rect 7524 25100 7530 25152
rect 7650 25100 7656 25152
rect 7708 25100 7714 25152
rect 8202 25100 8208 25152
rect 8260 25140 8266 25152
rect 9769 25143 9827 25149
rect 9769 25140 9781 25143
rect 8260 25112 9781 25140
rect 8260 25100 8266 25112
rect 9769 25109 9781 25112
rect 9815 25140 9827 25143
rect 10612 25140 10640 25180
rect 11146 25168 11152 25180
rect 11204 25208 11210 25220
rect 11348 25208 11376 25239
rect 11790 25236 11796 25288
rect 11848 25236 11854 25288
rect 12268 25285 12296 25316
rect 14737 25313 14749 25316
rect 14783 25313 14795 25347
rect 14737 25307 14795 25313
rect 11977 25279 12035 25285
rect 11977 25276 11989 25279
rect 11900 25248 11989 25276
rect 11204 25180 11376 25208
rect 11204 25168 11210 25180
rect 11606 25168 11612 25220
rect 11664 25168 11670 25220
rect 11900 25152 11928 25248
rect 11977 25245 11989 25248
rect 12023 25245 12035 25279
rect 12253 25279 12311 25285
rect 12253 25276 12265 25279
rect 11977 25239 12035 25245
rect 12084 25248 12265 25276
rect 12084 25152 12112 25248
rect 12253 25245 12265 25248
rect 12299 25245 12311 25279
rect 12253 25239 12311 25245
rect 12526 25236 12532 25288
rect 12584 25236 12590 25288
rect 14752 25276 14780 25307
rect 15289 25279 15347 25285
rect 15289 25276 15301 25279
rect 14752 25248 15301 25276
rect 15289 25245 15301 25248
rect 15335 25276 15347 25279
rect 15378 25276 15384 25288
rect 15335 25248 15384 25276
rect 15335 25245 15347 25248
rect 15289 25239 15347 25245
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 15488 25285 15516 25384
rect 15654 25372 15660 25384
rect 15712 25372 15718 25424
rect 16301 25415 16359 25421
rect 16301 25381 16313 25415
rect 16347 25412 16359 25415
rect 16390 25412 16396 25424
rect 16347 25384 16396 25412
rect 16347 25381 16359 25384
rect 16301 25375 16359 25381
rect 16390 25372 16396 25384
rect 16448 25372 16454 25424
rect 18233 25415 18291 25421
rect 18233 25381 18245 25415
rect 18279 25412 18291 25415
rect 18414 25412 18420 25424
rect 18279 25384 18420 25412
rect 18279 25381 18291 25384
rect 18233 25375 18291 25381
rect 18414 25372 18420 25384
rect 18472 25372 18478 25424
rect 18598 25372 18604 25424
rect 18656 25372 18662 25424
rect 18877 25415 18935 25421
rect 18877 25381 18889 25415
rect 18923 25412 18935 25415
rect 20272 25412 20300 25452
rect 20438 25440 20444 25452
rect 20496 25440 20502 25492
rect 20990 25440 20996 25492
rect 21048 25480 21054 25492
rect 21269 25483 21327 25489
rect 21269 25480 21281 25483
rect 21048 25452 21281 25480
rect 21048 25440 21054 25452
rect 21269 25449 21281 25452
rect 21315 25449 21327 25483
rect 21269 25443 21327 25449
rect 23293 25483 23351 25489
rect 23293 25449 23305 25483
rect 23339 25480 23351 25483
rect 24394 25480 24400 25492
rect 23339 25452 24400 25480
rect 23339 25449 23351 25452
rect 23293 25443 23351 25449
rect 24394 25440 24400 25452
rect 24452 25440 24458 25492
rect 18923 25384 20300 25412
rect 21913 25415 21971 25421
rect 18923 25381 18935 25384
rect 18877 25375 18935 25381
rect 21913 25381 21925 25415
rect 21959 25412 21971 25415
rect 21959 25384 22968 25412
rect 21959 25381 21971 25384
rect 21913 25375 21971 25381
rect 18049 25347 18107 25353
rect 15580 25316 16252 25344
rect 15580 25285 15608 25316
rect 16224 25288 16252 25316
rect 18049 25313 18061 25347
rect 18095 25344 18107 25347
rect 18509 25347 18567 25353
rect 18095 25316 18184 25344
rect 18095 25313 18107 25316
rect 18049 25307 18107 25313
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 15473 25239 15531 25245
rect 15565 25279 15623 25285
rect 15565 25245 15577 25279
rect 15611 25245 15623 25279
rect 15565 25239 15623 25245
rect 15657 25279 15715 25285
rect 15657 25245 15669 25279
rect 15703 25276 15715 25279
rect 16025 25279 16083 25285
rect 16025 25276 16037 25279
rect 15703 25248 16037 25276
rect 15703 25245 15715 25248
rect 15657 25239 15715 25245
rect 16025 25245 16037 25248
rect 16071 25245 16083 25279
rect 16025 25239 16083 25245
rect 15580 25208 15608 25239
rect 15120 25180 15608 25208
rect 15120 25152 15148 25180
rect 9815 25112 10640 25140
rect 9815 25109 9827 25112
rect 9769 25103 9827 25109
rect 11882 25100 11888 25152
rect 11940 25100 11946 25152
rect 12066 25100 12072 25152
rect 12124 25100 12130 25152
rect 13170 25100 13176 25152
rect 13228 25140 13234 25152
rect 15102 25140 15108 25152
rect 13228 25112 15108 25140
rect 13228 25100 13234 25112
rect 15102 25100 15108 25112
rect 15160 25100 15166 25152
rect 15470 25100 15476 25152
rect 15528 25140 15534 25152
rect 15672 25140 15700 25239
rect 16206 25236 16212 25288
rect 16264 25276 16270 25288
rect 16669 25279 16727 25285
rect 16669 25276 16681 25279
rect 16264 25248 16681 25276
rect 16264 25236 16270 25248
rect 16669 25245 16681 25248
rect 16715 25245 16727 25279
rect 16669 25239 16727 25245
rect 17586 25168 17592 25220
rect 17644 25208 17650 25220
rect 17865 25211 17923 25217
rect 17865 25208 17877 25211
rect 17644 25180 17877 25208
rect 17644 25168 17650 25180
rect 17865 25177 17877 25180
rect 17911 25177 17923 25211
rect 18156 25208 18184 25316
rect 18509 25313 18521 25347
rect 18555 25344 18567 25347
rect 18555 25316 19380 25344
rect 18555 25313 18567 25316
rect 18509 25307 18567 25313
rect 18230 25236 18236 25288
rect 18288 25276 18294 25288
rect 18417 25279 18475 25285
rect 18417 25276 18429 25279
rect 18288 25248 18429 25276
rect 18288 25236 18294 25248
rect 18417 25245 18429 25248
rect 18463 25245 18475 25279
rect 18417 25239 18475 25245
rect 18524 25208 18552 25307
rect 19352 25288 19380 25316
rect 20898 25304 20904 25356
rect 20956 25344 20962 25356
rect 22940 25353 22968 25384
rect 23014 25372 23020 25424
rect 23072 25412 23078 25424
rect 23477 25415 23535 25421
rect 23477 25412 23489 25415
rect 23072 25384 23489 25412
rect 23072 25372 23078 25384
rect 23477 25381 23489 25384
rect 23523 25381 23535 25415
rect 23477 25375 23535 25381
rect 21453 25347 21511 25353
rect 21453 25344 21465 25347
rect 20956 25316 21465 25344
rect 20956 25304 20962 25316
rect 21453 25313 21465 25316
rect 21499 25313 21511 25347
rect 21453 25307 21511 25313
rect 22925 25347 22983 25353
rect 22925 25313 22937 25347
rect 22971 25344 22983 25347
rect 22971 25316 23520 25344
rect 22971 25313 22983 25316
rect 22925 25307 22983 25313
rect 18693 25279 18751 25285
rect 18693 25276 18705 25279
rect 18156 25180 18552 25208
rect 18616 25248 18705 25276
rect 17865 25171 17923 25177
rect 15528 25112 15700 25140
rect 17880 25140 17908 25171
rect 18616 25140 18644 25248
rect 18693 25245 18705 25248
rect 18739 25245 18751 25279
rect 18693 25239 18751 25245
rect 19334 25236 19340 25288
rect 19392 25236 19398 25288
rect 20073 25279 20131 25285
rect 20073 25245 20085 25279
rect 20119 25276 20131 25279
rect 20346 25276 20352 25288
rect 20119 25248 20352 25276
rect 20119 25245 20131 25248
rect 20073 25239 20131 25245
rect 20346 25236 20352 25248
rect 20404 25236 20410 25288
rect 20441 25279 20499 25285
rect 20441 25245 20453 25279
rect 20487 25245 20499 25279
rect 20441 25239 20499 25245
rect 19426 25168 19432 25220
rect 19484 25208 19490 25220
rect 19705 25211 19763 25217
rect 19705 25208 19717 25211
rect 19484 25180 19717 25208
rect 19484 25168 19490 25180
rect 19705 25177 19717 25180
rect 19751 25177 19763 25211
rect 19705 25171 19763 25177
rect 19889 25211 19947 25217
rect 19889 25177 19901 25211
rect 19935 25208 19947 25211
rect 19978 25208 19984 25220
rect 19935 25180 19984 25208
rect 19935 25177 19947 25180
rect 19889 25171 19947 25177
rect 19978 25168 19984 25180
rect 20036 25168 20042 25220
rect 17880 25112 18644 25140
rect 20456 25140 20484 25239
rect 20530 25236 20536 25288
rect 20588 25276 20594 25288
rect 20625 25279 20683 25285
rect 20625 25276 20637 25279
rect 20588 25248 20637 25276
rect 20588 25236 20594 25248
rect 20625 25245 20637 25248
rect 20671 25245 20683 25279
rect 20625 25239 20683 25245
rect 20717 25279 20775 25285
rect 20717 25245 20729 25279
rect 20763 25245 20775 25279
rect 20717 25239 20775 25245
rect 20732 25208 20760 25239
rect 20806 25236 20812 25288
rect 20864 25236 20870 25288
rect 20990 25236 20996 25288
rect 21048 25276 21054 25288
rect 21085 25279 21143 25285
rect 21085 25276 21097 25279
rect 21048 25248 21097 25276
rect 21048 25236 21054 25248
rect 21085 25245 21097 25248
rect 21131 25245 21143 25279
rect 21085 25239 21143 25245
rect 21545 25279 21603 25285
rect 21545 25245 21557 25279
rect 21591 25245 21603 25279
rect 21545 25239 21603 25245
rect 23017 25279 23075 25285
rect 23017 25245 23029 25279
rect 23063 25276 23075 25279
rect 23106 25276 23112 25288
rect 23063 25248 23112 25276
rect 23063 25245 23075 25248
rect 23017 25239 23075 25245
rect 21008 25208 21036 25236
rect 20732 25180 21036 25208
rect 20806 25140 20812 25152
rect 20456 25112 20812 25140
rect 15528 25100 15534 25112
rect 20806 25100 20812 25112
rect 20864 25140 20870 25152
rect 20901 25143 20959 25149
rect 20901 25140 20913 25143
rect 20864 25112 20913 25140
rect 20864 25100 20870 25112
rect 20901 25109 20913 25112
rect 20947 25140 20959 25143
rect 21560 25140 21588 25239
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23492 25285 23520 25316
rect 23477 25279 23535 25285
rect 23477 25245 23489 25279
rect 23523 25245 23535 25279
rect 23477 25239 23535 25245
rect 23658 25236 23664 25288
rect 23716 25276 23722 25288
rect 23937 25279 23995 25285
rect 23937 25276 23949 25279
rect 23716 25248 23949 25276
rect 23716 25236 23722 25248
rect 23937 25245 23949 25248
rect 23983 25245 23995 25279
rect 23937 25239 23995 25245
rect 33134 25236 33140 25288
rect 33192 25236 33198 25288
rect 34330 25168 34336 25220
rect 34388 25168 34394 25220
rect 20947 25112 21588 25140
rect 20947 25109 20959 25112
rect 20901 25103 20959 25109
rect 1104 25050 35236 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 35236 25050
rect 1104 24976 35236 24998
rect 7006 24896 7012 24948
rect 7064 24896 7070 24948
rect 7282 24896 7288 24948
rect 7340 24936 7346 24948
rect 7926 24936 7932 24948
rect 7340 24908 7932 24936
rect 7340 24896 7346 24908
rect 7926 24896 7932 24908
rect 7984 24896 7990 24948
rect 11146 24896 11152 24948
rect 11204 24896 11210 24948
rect 11698 24896 11704 24948
rect 11756 24936 11762 24948
rect 12066 24936 12072 24948
rect 11756 24908 12072 24936
rect 11756 24896 11762 24908
rect 12066 24896 12072 24908
rect 12124 24896 12130 24948
rect 12618 24896 12624 24948
rect 12676 24936 12682 24948
rect 12713 24939 12771 24945
rect 12713 24936 12725 24939
rect 12676 24908 12725 24936
rect 12676 24896 12682 24908
rect 12713 24905 12725 24908
rect 12759 24936 12771 24939
rect 13538 24936 13544 24948
rect 12759 24908 13544 24936
rect 12759 24905 12771 24908
rect 12713 24899 12771 24905
rect 13538 24896 13544 24908
rect 13596 24896 13602 24948
rect 13909 24939 13967 24945
rect 13909 24905 13921 24939
rect 13955 24936 13967 24939
rect 13955 24908 14412 24936
rect 13955 24905 13967 24908
rect 13909 24899 13967 24905
rect 7024 24868 7052 24896
rect 9956 24880 10008 24886
rect 7834 24868 7840 24880
rect 7024 24840 7840 24868
rect 7834 24828 7840 24840
rect 7892 24868 7898 24880
rect 7892 24840 8524 24868
rect 7892 24828 7898 24840
rect 8496 24812 8524 24840
rect 11164 24868 11192 24896
rect 12437 24871 12495 24877
rect 12437 24868 12449 24871
rect 11164 24840 12449 24868
rect 12437 24837 12449 24840
rect 12483 24868 12495 24871
rect 13170 24868 13176 24880
rect 12483 24840 13176 24868
rect 12483 24837 12495 24840
rect 12437 24831 12495 24837
rect 9956 24822 10008 24828
rect 5169 24803 5227 24809
rect 5169 24769 5181 24803
rect 5215 24800 5227 24803
rect 5442 24800 5448 24812
rect 5215 24772 5448 24800
rect 5215 24769 5227 24772
rect 5169 24763 5227 24769
rect 5442 24760 5448 24772
rect 5500 24800 5506 24812
rect 5629 24803 5687 24809
rect 5629 24800 5641 24803
rect 5500 24772 5641 24800
rect 5500 24760 5506 24772
rect 5629 24769 5641 24772
rect 5675 24769 5687 24803
rect 5629 24763 5687 24769
rect 6914 24760 6920 24812
rect 6972 24760 6978 24812
rect 7466 24760 7472 24812
rect 7524 24760 7530 24812
rect 8478 24760 8484 24812
rect 8536 24760 8542 24812
rect 9214 24760 9220 24812
rect 9272 24760 9278 24812
rect 10597 24803 10655 24809
rect 10597 24800 10609 24803
rect 10520 24772 10609 24800
rect 10520 24744 10548 24772
rect 10597 24769 10609 24772
rect 10643 24800 10655 24803
rect 10778 24800 10784 24812
rect 10643 24772 10784 24800
rect 10643 24769 10655 24772
rect 10597 24763 10655 24769
rect 10778 24760 10784 24772
rect 10836 24800 10842 24812
rect 12636 24809 12664 24840
rect 13170 24828 13176 24840
rect 13228 24828 13234 24880
rect 12621 24803 12679 24809
rect 10836 24772 12572 24800
rect 10836 24760 10842 24772
rect 10502 24692 10508 24744
rect 10560 24692 10566 24744
rect 10689 24735 10747 24741
rect 10689 24701 10701 24735
rect 10735 24732 10747 24735
rect 11606 24732 11612 24744
rect 10735 24704 11612 24732
rect 10735 24701 10747 24704
rect 10689 24695 10747 24701
rect 11606 24692 11612 24704
rect 11664 24692 11670 24744
rect 12544 24732 12572 24772
rect 12621 24769 12633 24803
rect 12667 24769 12679 24803
rect 12621 24763 12679 24769
rect 12805 24803 12863 24809
rect 12805 24769 12817 24803
rect 12851 24769 12863 24803
rect 12805 24763 12863 24769
rect 12820 24732 12848 24763
rect 13354 24760 13360 24812
rect 13412 24800 13418 24812
rect 13633 24803 13691 24809
rect 13633 24800 13645 24803
rect 13412 24772 13645 24800
rect 13412 24760 13418 24772
rect 13633 24769 13645 24772
rect 13679 24769 13691 24803
rect 13633 24763 13691 24769
rect 14001 24803 14059 24809
rect 14001 24769 14013 24803
rect 14047 24769 14059 24803
rect 14384 24800 14412 24908
rect 15102 24896 15108 24948
rect 15160 24936 15166 24948
rect 15289 24939 15347 24945
rect 15289 24936 15301 24939
rect 15160 24908 15301 24936
rect 15160 24896 15166 24908
rect 15289 24905 15301 24908
rect 15335 24905 15347 24939
rect 15289 24899 15347 24905
rect 15378 24896 15384 24948
rect 15436 24936 15442 24948
rect 15436 24908 15700 24936
rect 15436 24896 15442 24908
rect 15672 24812 15700 24908
rect 19334 24896 19340 24948
rect 19392 24936 19398 24948
rect 19797 24939 19855 24945
rect 19797 24936 19809 24939
rect 19392 24908 19809 24936
rect 19392 24896 19398 24908
rect 19797 24905 19809 24908
rect 19843 24905 19855 24939
rect 19797 24899 19855 24905
rect 20990 24896 20996 24948
rect 21048 24896 21054 24948
rect 19426 24868 19432 24880
rect 16132 24840 16344 24868
rect 14550 24800 14556 24812
rect 14384 24772 14556 24800
rect 14001 24763 14059 24769
rect 12544 24704 12848 24732
rect 13814 24692 13820 24744
rect 13872 24732 13878 24744
rect 13909 24735 13967 24741
rect 13909 24732 13921 24735
rect 13872 24704 13921 24732
rect 13872 24692 13878 24704
rect 13909 24701 13921 24704
rect 13955 24732 13967 24735
rect 14016 24732 14044 24763
rect 14550 24760 14556 24772
rect 14608 24760 14614 24812
rect 14645 24803 14703 24809
rect 14645 24769 14657 24803
rect 14691 24769 14703 24803
rect 14645 24763 14703 24769
rect 13955 24704 14044 24732
rect 13955 24701 13967 24704
rect 13909 24695 13967 24701
rect 14090 24692 14096 24744
rect 14148 24692 14154 24744
rect 8297 24667 8355 24673
rect 8297 24633 8309 24667
rect 8343 24664 8355 24667
rect 11330 24664 11336 24676
rect 8343 24636 11336 24664
rect 8343 24633 8355 24636
rect 8297 24627 8355 24633
rect 11330 24624 11336 24636
rect 11388 24624 11394 24676
rect 13354 24624 13360 24676
rect 13412 24624 13418 24676
rect 13722 24624 13728 24676
rect 13780 24664 13786 24676
rect 14369 24667 14427 24673
rect 13780 24636 14228 24664
rect 13780 24624 13786 24636
rect 5166 24556 5172 24608
rect 5224 24596 5230 24608
rect 5261 24599 5319 24605
rect 5261 24596 5273 24599
rect 5224 24568 5273 24596
rect 5224 24556 5230 24568
rect 5261 24565 5273 24568
rect 5307 24565 5319 24599
rect 5261 24559 5319 24565
rect 6086 24556 6092 24608
rect 6144 24556 6150 24608
rect 13372 24596 13400 24624
rect 14090 24596 14096 24608
rect 13372 24568 14096 24596
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14200 24605 14228 24636
rect 14369 24633 14381 24667
rect 14415 24664 14427 24667
rect 14660 24664 14688 24763
rect 15010 24760 15016 24812
rect 15068 24800 15074 24812
rect 15470 24800 15476 24812
rect 15068 24772 15476 24800
rect 15068 24760 15074 24772
rect 15470 24760 15476 24772
rect 15528 24760 15534 24812
rect 15654 24809 15660 24812
rect 15627 24803 15660 24809
rect 15627 24769 15639 24803
rect 15627 24763 15660 24769
rect 15654 24760 15660 24763
rect 15712 24760 15718 24812
rect 16132 24800 16160 24840
rect 15764 24772 16160 24800
rect 14829 24735 14887 24741
rect 14829 24701 14841 24735
rect 14875 24732 14887 24735
rect 15764 24732 15792 24772
rect 16206 24760 16212 24812
rect 16264 24760 16270 24812
rect 16316 24800 16344 24840
rect 19168 24840 19432 24868
rect 19168 24800 19196 24840
rect 19426 24828 19432 24840
rect 19484 24828 19490 24880
rect 19628 24840 19840 24868
rect 16316 24772 19196 24800
rect 19245 24803 19303 24809
rect 19245 24769 19257 24803
rect 19291 24800 19303 24803
rect 19334 24800 19340 24812
rect 19291 24772 19340 24800
rect 19291 24769 19303 24772
rect 19245 24763 19303 24769
rect 19334 24760 19340 24772
rect 19392 24800 19398 24812
rect 19628 24800 19656 24840
rect 19392 24772 19656 24800
rect 19705 24803 19763 24809
rect 19392 24760 19398 24772
rect 19705 24769 19717 24803
rect 19751 24769 19763 24803
rect 19812 24800 19840 24840
rect 20456 24840 21128 24868
rect 19889 24803 19947 24809
rect 19889 24800 19901 24803
rect 19812 24772 19901 24800
rect 19705 24763 19763 24769
rect 19889 24769 19901 24772
rect 19935 24769 19947 24803
rect 19889 24763 19947 24769
rect 14875 24704 15792 24732
rect 15841 24735 15899 24741
rect 14875 24701 14887 24704
rect 14829 24695 14887 24701
rect 15841 24701 15853 24735
rect 15887 24732 15899 24735
rect 15933 24735 15991 24741
rect 15933 24732 15945 24735
rect 15887 24704 15945 24732
rect 15887 24701 15899 24704
rect 15841 24695 15899 24701
rect 15933 24701 15945 24704
rect 15979 24701 15991 24735
rect 15933 24695 15991 24701
rect 16114 24692 16120 24744
rect 16172 24692 16178 24744
rect 19153 24735 19211 24741
rect 19153 24732 19165 24735
rect 18524 24704 19165 24732
rect 14415 24636 14688 24664
rect 16025 24667 16083 24673
rect 14415 24633 14427 24636
rect 14369 24627 14427 24633
rect 16025 24633 16037 24667
rect 16071 24664 16083 24667
rect 16132 24664 16160 24692
rect 16071 24636 16160 24664
rect 16071 24633 16083 24636
rect 16025 24627 16083 24633
rect 18524 24608 18552 24704
rect 19153 24701 19165 24704
rect 19199 24732 19211 24735
rect 19720 24732 19748 24763
rect 19199 24704 19748 24732
rect 19199 24701 19211 24704
rect 19153 24695 19211 24701
rect 19794 24692 19800 24744
rect 19852 24732 19858 24744
rect 20456 24741 20484 24840
rect 20533 24803 20591 24809
rect 20533 24769 20545 24803
rect 20579 24800 20591 24803
rect 21100 24800 21128 24840
rect 21177 24803 21235 24809
rect 21177 24800 21189 24803
rect 20579 24772 21036 24800
rect 21100 24772 21189 24800
rect 20579 24769 20591 24772
rect 20533 24763 20591 24769
rect 20441 24735 20499 24741
rect 20441 24732 20453 24735
rect 19852 24704 20453 24732
rect 19852 24692 19858 24704
rect 20441 24701 20453 24704
rect 20487 24701 20499 24735
rect 20441 24695 20499 24701
rect 19613 24667 19671 24673
rect 19613 24633 19625 24667
rect 19659 24664 19671 24667
rect 19978 24664 19984 24676
rect 19659 24636 19984 24664
rect 19659 24633 19671 24636
rect 19613 24627 19671 24633
rect 19978 24624 19984 24636
rect 20036 24664 20042 24676
rect 20548 24664 20576 24763
rect 20898 24692 20904 24744
rect 20956 24692 20962 24744
rect 21008 24732 21036 24772
rect 21177 24769 21189 24772
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 21361 24735 21419 24741
rect 21361 24732 21373 24735
rect 21008 24704 21373 24732
rect 21361 24701 21373 24704
rect 21407 24701 21419 24735
rect 21361 24695 21419 24701
rect 20036 24636 20576 24664
rect 20036 24624 20042 24636
rect 14185 24599 14243 24605
rect 14185 24565 14197 24599
rect 14231 24565 14243 24599
rect 14185 24559 14243 24565
rect 16114 24556 16120 24608
rect 16172 24556 16178 24608
rect 18506 24556 18512 24608
rect 18564 24556 18570 24608
rect 1104 24506 35248 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 35248 24506
rect 1104 24432 35248 24454
rect 6196 24364 8064 24392
rect 6196 24265 6224 24364
rect 8036 24336 8064 24364
rect 8846 24352 8852 24404
rect 8904 24392 8910 24404
rect 11149 24395 11207 24401
rect 11149 24392 11161 24395
rect 8904 24364 11161 24392
rect 8904 24352 8910 24364
rect 11149 24361 11161 24364
rect 11195 24361 11207 24395
rect 11149 24355 11207 24361
rect 11609 24395 11667 24401
rect 11609 24361 11621 24395
rect 11655 24392 11667 24395
rect 11790 24392 11796 24404
rect 11655 24364 11796 24392
rect 11655 24361 11667 24364
rect 11609 24355 11667 24361
rect 6641 24327 6699 24333
rect 6641 24293 6653 24327
rect 6687 24324 6699 24327
rect 6687 24296 7052 24324
rect 6687 24293 6699 24296
rect 6641 24287 6699 24293
rect 6181 24259 6239 24265
rect 6181 24225 6193 24259
rect 6227 24225 6239 24259
rect 6181 24219 6239 24225
rect 934 24148 940 24200
rect 992 24188 998 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 992 24160 1409 24188
rect 992 24148 998 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 3602 24148 3608 24200
rect 3660 24188 3666 24200
rect 4062 24188 4068 24200
rect 3660 24160 4068 24188
rect 3660 24148 3666 24160
rect 4062 24148 4068 24160
rect 4120 24188 4126 24200
rect 4157 24191 4215 24197
rect 4157 24188 4169 24191
rect 4120 24160 4169 24188
rect 4120 24148 4126 24160
rect 4157 24157 4169 24160
rect 4203 24157 4215 24191
rect 4157 24151 4215 24157
rect 6549 24191 6607 24197
rect 6549 24157 6561 24191
rect 6595 24157 6607 24191
rect 6549 24151 6607 24157
rect 6733 24191 6791 24197
rect 6733 24157 6745 24191
rect 6779 24157 6791 24191
rect 7024 24188 7052 24296
rect 8018 24284 8024 24336
rect 8076 24284 8082 24336
rect 11164 24324 11192 24355
rect 11790 24352 11796 24364
rect 11848 24352 11854 24404
rect 11882 24352 11888 24404
rect 11940 24352 11946 24404
rect 11974 24352 11980 24404
rect 12032 24392 12038 24404
rect 12161 24395 12219 24401
rect 12161 24392 12173 24395
rect 12032 24364 12173 24392
rect 12032 24352 12038 24364
rect 12161 24361 12173 24364
rect 12207 24361 12219 24395
rect 12161 24355 12219 24361
rect 12434 24352 12440 24404
rect 12492 24392 12498 24404
rect 12529 24395 12587 24401
rect 12529 24392 12541 24395
rect 12492 24364 12541 24392
rect 12492 24352 12498 24364
rect 12529 24361 12541 24364
rect 12575 24392 12587 24395
rect 12710 24392 12716 24404
rect 12575 24364 12716 24392
rect 12575 24361 12587 24364
rect 12529 24355 12587 24361
rect 12710 24352 12716 24364
rect 12768 24352 12774 24404
rect 12802 24352 12808 24404
rect 12860 24352 12866 24404
rect 13633 24395 13691 24401
rect 13633 24361 13645 24395
rect 13679 24392 13691 24395
rect 13722 24392 13728 24404
rect 13679 24364 13728 24392
rect 13679 24361 13691 24364
rect 13633 24355 13691 24361
rect 13722 24352 13728 24364
rect 13780 24352 13786 24404
rect 14277 24395 14335 24401
rect 14277 24392 14289 24395
rect 13832 24364 14289 24392
rect 12250 24324 12256 24336
rect 11164 24296 12256 24324
rect 9214 24216 9220 24268
rect 9272 24216 9278 24268
rect 7469 24191 7527 24197
rect 7469 24188 7481 24191
rect 7024 24160 7481 24188
rect 6733 24151 6791 24157
rect 7469 24157 7481 24160
rect 7515 24157 7527 24191
rect 7469 24151 7527 24157
rect 4433 24123 4491 24129
rect 4433 24120 4445 24123
rect 1596 24092 4445 24120
rect 1596 24061 1624 24092
rect 4433 24089 4445 24092
rect 4479 24089 4491 24123
rect 4433 24083 4491 24089
rect 5166 24080 5172 24132
rect 5224 24080 5230 24132
rect 1581 24055 1639 24061
rect 1581 24021 1593 24055
rect 1627 24021 1639 24055
rect 6564 24052 6592 24151
rect 6748 24120 6776 24151
rect 8018 24148 8024 24200
rect 8076 24148 8082 24200
rect 8478 24148 8484 24200
rect 8536 24188 8542 24200
rect 9125 24191 9183 24197
rect 9125 24188 9137 24191
rect 8536 24160 9137 24188
rect 8536 24148 8542 24160
rect 9125 24157 9137 24160
rect 9171 24157 9183 24191
rect 9125 24151 9183 24157
rect 11330 24148 11336 24200
rect 11388 24148 11394 24200
rect 11422 24148 11428 24200
rect 11480 24148 11486 24200
rect 11716 24197 11744 24296
rect 12250 24284 12256 24296
rect 12308 24324 12314 24336
rect 12820 24324 12848 24352
rect 13832 24333 13860 24364
rect 14277 24361 14289 24364
rect 14323 24361 14335 24395
rect 14277 24355 14335 24361
rect 15102 24352 15108 24404
rect 15160 24392 15166 24404
rect 15289 24395 15347 24401
rect 15289 24392 15301 24395
rect 15160 24364 15301 24392
rect 15160 24352 15166 24364
rect 15289 24361 15301 24364
rect 15335 24392 15347 24395
rect 16114 24392 16120 24404
rect 15335 24364 16120 24392
rect 15335 24361 15347 24364
rect 15289 24355 15347 24361
rect 16114 24352 16120 24364
rect 16172 24352 16178 24404
rect 17586 24352 17592 24404
rect 17644 24352 17650 24404
rect 18506 24352 18512 24404
rect 18564 24352 18570 24404
rect 18598 24352 18604 24404
rect 18656 24352 18662 24404
rect 24118 24352 24124 24404
rect 24176 24352 24182 24404
rect 13817 24327 13875 24333
rect 13817 24324 13829 24327
rect 12308 24296 12480 24324
rect 12820 24296 13829 24324
rect 12308 24284 12314 24296
rect 11793 24259 11851 24265
rect 11793 24225 11805 24259
rect 11839 24225 11851 24259
rect 11793 24219 11851 24225
rect 11885 24259 11943 24265
rect 11885 24225 11897 24259
rect 11931 24256 11943 24259
rect 12069 24259 12127 24265
rect 11931 24228 12020 24256
rect 11931 24225 11943 24228
rect 11885 24219 11943 24225
rect 11701 24191 11759 24197
rect 11701 24157 11713 24191
rect 11747 24157 11759 24191
rect 11701 24151 11759 24157
rect 7282 24120 7288 24132
rect 6748 24092 7288 24120
rect 7282 24080 7288 24092
rect 7340 24080 7346 24132
rect 9674 24120 9680 24132
rect 8418 24092 9680 24120
rect 9674 24080 9680 24092
rect 9732 24120 9738 24132
rect 10502 24120 10508 24132
rect 9732 24092 10508 24120
rect 9732 24080 9738 24092
rect 10502 24080 10508 24092
rect 10560 24080 10566 24132
rect 11149 24123 11207 24129
rect 11149 24089 11161 24123
rect 11195 24089 11207 24123
rect 11348 24120 11376 24148
rect 11808 24120 11836 24219
rect 11992 24200 12020 24228
rect 12069 24225 12081 24259
rect 12115 24256 12127 24259
rect 12342 24256 12348 24268
rect 12115 24228 12348 24256
rect 12115 24225 12127 24228
rect 12069 24219 12127 24225
rect 11974 24148 11980 24200
rect 12032 24148 12038 24200
rect 11882 24120 11888 24132
rect 11348 24092 11888 24120
rect 11149 24083 11207 24089
rect 7098 24052 7104 24064
rect 6564 24024 7104 24052
rect 1581 24015 1639 24021
rect 7098 24012 7104 24024
rect 7156 24052 7162 24064
rect 7374 24052 7380 24064
rect 7156 24024 7380 24052
rect 7156 24012 7162 24024
rect 7374 24012 7380 24024
rect 7432 24012 7438 24064
rect 9490 24012 9496 24064
rect 9548 24012 9554 24064
rect 11164 24052 11192 24083
rect 11882 24080 11888 24092
rect 11940 24080 11946 24132
rect 12084 24052 12112 24219
rect 12342 24216 12348 24228
rect 12400 24216 12406 24268
rect 12452 24265 12480 24296
rect 13817 24293 13829 24296
rect 13863 24293 13875 24327
rect 13817 24287 13875 24293
rect 15654 24284 15660 24336
rect 15712 24284 15718 24336
rect 18693 24327 18751 24333
rect 18693 24324 18705 24327
rect 18156 24296 18705 24324
rect 12437 24259 12495 24265
rect 12437 24225 12449 24259
rect 12483 24256 12495 24259
rect 12483 24228 12848 24256
rect 12483 24225 12495 24228
rect 12437 24219 12495 24225
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 11164 24024 12112 24052
rect 12544 24052 12572 24151
rect 12618 24148 12624 24200
rect 12676 24148 12682 24200
rect 12820 24197 12848 24228
rect 16758 24216 16764 24268
rect 16816 24256 16822 24268
rect 17037 24259 17095 24265
rect 17037 24256 17049 24259
rect 16816 24228 17049 24256
rect 16816 24216 16822 24228
rect 17037 24225 17049 24228
rect 17083 24225 17095 24259
rect 17037 24219 17095 24225
rect 17313 24259 17371 24265
rect 17313 24225 17325 24259
rect 17359 24256 17371 24259
rect 18156 24256 18184 24296
rect 18693 24293 18705 24296
rect 18739 24293 18751 24327
rect 18693 24287 18751 24293
rect 17359 24228 18184 24256
rect 17359 24225 17371 24228
rect 17313 24219 17371 24225
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24157 12863 24191
rect 12805 24151 12863 24157
rect 12989 24191 13047 24197
rect 12989 24157 13001 24191
rect 13035 24188 13047 24191
rect 13078 24188 13084 24200
rect 13035 24160 13084 24188
rect 13035 24157 13047 24160
rect 12989 24151 13047 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13173 24191 13231 24197
rect 13173 24157 13185 24191
rect 13219 24157 13231 24191
rect 13173 24151 13231 24157
rect 12710 24080 12716 24132
rect 12768 24120 12774 24132
rect 13188 24120 13216 24151
rect 13262 24148 13268 24200
rect 13320 24148 13326 24200
rect 13357 24191 13415 24197
rect 13357 24157 13369 24191
rect 13403 24190 13415 24191
rect 13403 24162 13492 24190
rect 13403 24157 13415 24162
rect 13357 24151 13415 24157
rect 12768 24092 13216 24120
rect 12768 24080 12774 24092
rect 12802 24052 12808 24064
rect 12544 24024 12808 24052
rect 12802 24012 12808 24024
rect 12860 24052 12866 24064
rect 13464 24052 13492 24162
rect 13538 24148 13544 24200
rect 13596 24188 13602 24200
rect 13725 24191 13783 24197
rect 13725 24188 13737 24191
rect 13596 24160 13737 24188
rect 13596 24148 13602 24160
rect 13725 24157 13737 24160
rect 13771 24157 13783 24191
rect 13909 24191 13967 24197
rect 13909 24188 13921 24191
rect 13725 24151 13783 24157
rect 13832 24160 13921 24188
rect 13832 24052 13860 24160
rect 13909 24157 13921 24160
rect 13955 24157 13967 24191
rect 13909 24151 13967 24157
rect 14918 24148 14924 24200
rect 14976 24188 14982 24200
rect 15194 24188 15200 24200
rect 14976 24160 15200 24188
rect 14976 24148 14982 24160
rect 15194 24148 15200 24160
rect 15252 24148 15258 24200
rect 14090 24080 14096 24132
rect 14148 24080 14154 24132
rect 16776 24120 16804 24216
rect 16850 24148 16856 24200
rect 16908 24188 16914 24200
rect 18156 24197 18184 24228
rect 18233 24259 18291 24265
rect 18233 24225 18245 24259
rect 18279 24225 18291 24259
rect 24136 24256 24164 24352
rect 24397 24259 24455 24265
rect 24397 24256 24409 24259
rect 24136 24228 24409 24256
rect 18233 24219 18291 24225
rect 24397 24225 24409 24228
rect 24443 24225 24455 24259
rect 24397 24219 24455 24225
rect 16945 24191 17003 24197
rect 16945 24188 16957 24191
rect 16908 24160 16957 24188
rect 16908 24148 16914 24160
rect 16945 24157 16957 24160
rect 16991 24188 17003 24191
rect 17405 24191 17463 24197
rect 17405 24188 17417 24191
rect 16991 24160 17417 24188
rect 16991 24157 17003 24160
rect 16945 24151 17003 24157
rect 17405 24157 17417 24160
rect 17451 24157 17463 24191
rect 17405 24151 17463 24157
rect 17589 24191 17647 24197
rect 17589 24157 17601 24191
rect 17635 24157 17647 24191
rect 17589 24151 17647 24157
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24157 18199 24191
rect 18141 24151 18199 24157
rect 17604 24120 17632 24151
rect 18248 24120 18276 24219
rect 19061 24123 19119 24129
rect 19061 24120 19073 24123
rect 16776 24092 17632 24120
rect 18156 24092 19073 24120
rect 18156 24064 18184 24092
rect 19061 24089 19073 24092
rect 19107 24089 19119 24123
rect 19061 24083 19119 24089
rect 24670 24080 24676 24132
rect 24728 24080 24734 24132
rect 24946 24080 24952 24132
rect 25004 24120 25010 24132
rect 25004 24092 25162 24120
rect 25004 24080 25010 24092
rect 12860 24024 13860 24052
rect 12860 24012 12866 24024
rect 13998 24012 14004 24064
rect 14056 24052 14062 24064
rect 14293 24055 14351 24061
rect 14293 24052 14305 24055
rect 14056 24024 14305 24052
rect 14056 24012 14062 24024
rect 14293 24021 14305 24024
rect 14339 24021 14351 24055
rect 14293 24015 14351 24021
rect 14458 24012 14464 24064
rect 14516 24012 14522 24064
rect 18138 24012 18144 24064
rect 18196 24012 18202 24064
rect 26145 24055 26203 24061
rect 26145 24021 26157 24055
rect 26191 24052 26203 24055
rect 33134 24052 33140 24064
rect 26191 24024 33140 24052
rect 26191 24021 26203 24024
rect 26145 24015 26203 24021
rect 33134 24012 33140 24024
rect 33192 24012 33198 24064
rect 1104 23962 35236 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 35236 23962
rect 1104 23888 35236 23910
rect 9214 23808 9220 23860
rect 9272 23808 9278 23860
rect 12710 23808 12716 23860
rect 12768 23848 12774 23860
rect 12768 23820 13216 23848
rect 12768 23808 12774 23820
rect 4982 23740 4988 23792
rect 5040 23740 5046 23792
rect 6914 23780 6920 23792
rect 6656 23752 6920 23780
rect 6178 23672 6184 23724
rect 6236 23712 6242 23724
rect 6656 23721 6684 23752
rect 6914 23740 6920 23752
rect 6972 23740 6978 23792
rect 7282 23740 7288 23792
rect 7340 23780 7346 23792
rect 9125 23783 9183 23789
rect 7340 23752 8432 23780
rect 7340 23740 7346 23752
rect 6641 23715 6699 23721
rect 6641 23712 6653 23715
rect 6236 23684 6653 23712
rect 6236 23672 6242 23684
rect 6641 23681 6653 23684
rect 6687 23681 6699 23715
rect 6641 23675 6699 23681
rect 6822 23672 6828 23724
rect 6880 23712 6886 23724
rect 7377 23715 7435 23721
rect 7377 23712 7389 23715
rect 6880 23684 7389 23712
rect 6880 23672 6886 23684
rect 7377 23681 7389 23684
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 7650 23672 7656 23724
rect 7708 23672 7714 23724
rect 8018 23672 8024 23724
rect 8076 23672 8082 23724
rect 8404 23721 8432 23752
rect 9125 23749 9137 23783
rect 9171 23780 9183 23783
rect 9232 23780 9260 23808
rect 9171 23752 9260 23780
rect 12345 23783 12403 23789
rect 9171 23749 9183 23752
rect 9125 23743 9183 23749
rect 12345 23749 12357 23783
rect 12391 23780 12403 23783
rect 12391 23752 12848 23780
rect 12391 23749 12403 23752
rect 12345 23743 12403 23749
rect 12820 23724 12848 23752
rect 8389 23715 8447 23721
rect 8389 23681 8401 23715
rect 8435 23681 8447 23715
rect 8389 23675 8447 23681
rect 8941 23715 8999 23721
rect 8941 23681 8953 23715
rect 8987 23712 8999 23715
rect 9766 23712 9772 23724
rect 8987 23684 9772 23712
rect 8987 23681 8999 23684
rect 8941 23675 8999 23681
rect 3602 23604 3608 23656
rect 3660 23644 3666 23656
rect 3973 23647 4031 23653
rect 3973 23644 3985 23647
rect 3660 23616 3985 23644
rect 3660 23604 3666 23616
rect 3973 23613 3985 23616
rect 4019 23613 4031 23647
rect 3973 23607 4031 23613
rect 4249 23647 4307 23653
rect 4249 23613 4261 23647
rect 4295 23644 4307 23647
rect 4614 23644 4620 23656
rect 4295 23616 4620 23644
rect 4295 23613 4307 23616
rect 4249 23607 4307 23613
rect 4614 23604 4620 23616
rect 4672 23604 4678 23656
rect 5994 23604 6000 23656
rect 6052 23604 6058 23656
rect 8202 23604 8208 23656
rect 8260 23644 8266 23656
rect 8956 23644 8984 23675
rect 9766 23672 9772 23684
rect 9824 23712 9830 23724
rect 9861 23715 9919 23721
rect 9861 23712 9873 23715
rect 9824 23684 9873 23712
rect 9824 23672 9830 23684
rect 9861 23681 9873 23684
rect 9907 23681 9919 23715
rect 9861 23675 9919 23681
rect 10410 23672 10416 23724
rect 10468 23712 10474 23724
rect 10505 23715 10563 23721
rect 10505 23712 10517 23715
rect 10468 23684 10517 23712
rect 10468 23672 10474 23684
rect 10505 23681 10517 23684
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 11422 23672 11428 23724
rect 11480 23712 11486 23724
rect 12066 23712 12072 23724
rect 11480 23684 12072 23712
rect 11480 23672 11486 23684
rect 12066 23672 12072 23684
rect 12124 23712 12130 23724
rect 12253 23715 12311 23721
rect 12253 23712 12265 23715
rect 12124 23684 12265 23712
rect 12124 23672 12130 23684
rect 12253 23681 12265 23684
rect 12299 23681 12311 23715
rect 12253 23675 12311 23681
rect 12437 23715 12495 23721
rect 12437 23681 12449 23715
rect 12483 23681 12495 23715
rect 12437 23675 12495 23681
rect 12452 23644 12480 23675
rect 12802 23672 12808 23724
rect 12860 23672 12866 23724
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 8260 23616 8984 23644
rect 11992 23616 12480 23644
rect 8260 23604 8266 23616
rect 11992 23588 12020 23616
rect 7101 23579 7159 23585
rect 7101 23545 7113 23579
rect 7147 23576 7159 23579
rect 10502 23576 10508 23588
rect 7147 23548 10508 23576
rect 7147 23545 7159 23548
rect 7101 23539 7159 23545
rect 10502 23536 10508 23548
rect 10560 23536 10566 23588
rect 11974 23536 11980 23588
rect 12032 23536 12038 23588
rect 12912 23576 12940 23675
rect 13078 23672 13084 23724
rect 13136 23672 13142 23724
rect 13188 23721 13216 23820
rect 13722 23808 13728 23860
rect 13780 23808 13786 23860
rect 13817 23851 13875 23857
rect 13817 23817 13829 23851
rect 13863 23848 13875 23851
rect 13998 23848 14004 23860
rect 13863 23820 14004 23848
rect 13863 23817 13875 23820
rect 13817 23811 13875 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 14458 23808 14464 23860
rect 14516 23808 14522 23860
rect 20806 23808 20812 23860
rect 20864 23848 20870 23860
rect 20901 23851 20959 23857
rect 20901 23848 20913 23851
rect 20864 23820 20913 23848
rect 20864 23808 20870 23820
rect 20901 23817 20913 23820
rect 20947 23817 20959 23851
rect 23658 23848 23664 23860
rect 20901 23811 20959 23817
rect 23032 23820 23664 23848
rect 13740 23721 13768 23808
rect 13173 23715 13231 23721
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13725 23715 13783 23721
rect 13725 23681 13737 23715
rect 13771 23681 13783 23715
rect 14476 23712 14504 23808
rect 23032 23724 23060 23820
rect 23658 23808 23664 23820
rect 23716 23808 23722 23860
rect 24670 23808 24676 23860
rect 24728 23808 24734 23860
rect 24946 23808 24952 23860
rect 25004 23808 25010 23860
rect 23106 23740 23112 23792
rect 23164 23740 23170 23792
rect 20622 23712 20628 23724
rect 14476 23684 20628 23712
rect 13725 23675 13783 23681
rect 20622 23672 20628 23684
rect 20680 23672 20686 23724
rect 21082 23672 21088 23724
rect 21140 23672 21146 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21468 23684 22017 23712
rect 21468 23656 21496 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22833 23715 22891 23721
rect 22833 23712 22845 23715
rect 22005 23675 22063 23681
rect 22388 23684 22845 23712
rect 13357 23647 13415 23653
rect 13357 23613 13369 23647
rect 13403 23644 13415 23647
rect 14090 23644 14096 23656
rect 13403 23616 14096 23644
rect 13403 23613 13415 23616
rect 13357 23607 13415 23613
rect 14090 23604 14096 23616
rect 14148 23604 14154 23656
rect 20438 23604 20444 23656
rect 20496 23604 20502 23656
rect 21361 23647 21419 23653
rect 21361 23613 21373 23647
rect 21407 23644 21419 23647
rect 21450 23644 21456 23656
rect 21407 23616 21456 23644
rect 21407 23613 21419 23616
rect 21361 23607 21419 23613
rect 21450 23604 21456 23616
rect 21508 23604 21514 23656
rect 21910 23604 21916 23656
rect 21968 23604 21974 23656
rect 13262 23576 13268 23588
rect 12912 23548 13268 23576
rect 13262 23536 13268 23548
rect 13320 23576 13326 23588
rect 13538 23576 13544 23588
rect 13320 23548 13544 23576
rect 13320 23536 13326 23548
rect 13538 23536 13544 23548
rect 13596 23536 13602 23588
rect 20809 23579 20867 23585
rect 20809 23545 20821 23579
rect 20855 23576 20867 23579
rect 21174 23576 21180 23588
rect 20855 23548 21180 23576
rect 20855 23545 20867 23548
rect 20809 23539 20867 23545
rect 21174 23536 21180 23548
rect 21232 23576 21238 23588
rect 22388 23585 22416 23684
rect 22833 23681 22845 23684
rect 22879 23681 22891 23715
rect 22833 23675 22891 23681
rect 22848 23644 22876 23675
rect 23014 23672 23020 23724
rect 23072 23672 23078 23724
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23712 23259 23715
rect 23382 23712 23388 23724
rect 23247 23684 23388 23712
rect 23247 23681 23259 23684
rect 23201 23675 23259 23681
rect 23382 23672 23388 23684
rect 23440 23712 23446 23724
rect 23477 23715 23535 23721
rect 23477 23712 23489 23715
rect 23440 23684 23489 23712
rect 23440 23672 23446 23684
rect 23477 23681 23489 23684
rect 23523 23681 23535 23715
rect 23477 23675 23535 23681
rect 23569 23647 23627 23653
rect 23569 23644 23581 23647
rect 22848 23616 23581 23644
rect 23569 23613 23581 23616
rect 23615 23613 23627 23647
rect 23569 23607 23627 23613
rect 23845 23647 23903 23653
rect 23845 23613 23857 23647
rect 23891 23644 23903 23647
rect 24688 23644 24716 23808
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23712 24915 23715
rect 24903 23684 25452 23712
rect 24903 23681 24915 23684
rect 24857 23675 24915 23681
rect 23891 23616 24716 23644
rect 23891 23613 23903 23616
rect 23845 23607 23903 23613
rect 21269 23579 21327 23585
rect 21269 23576 21281 23579
rect 21232 23548 21281 23576
rect 21232 23536 21238 23548
rect 21269 23545 21281 23548
rect 21315 23545 21327 23579
rect 21269 23539 21327 23545
rect 22373 23579 22431 23585
rect 22373 23545 22385 23579
rect 22419 23545 22431 23579
rect 22373 23539 22431 23545
rect 11333 23511 11391 23517
rect 11333 23477 11345 23511
rect 11379 23508 11391 23511
rect 11882 23508 11888 23520
rect 11379 23480 11888 23508
rect 11379 23477 11391 23480
rect 11333 23471 11391 23477
rect 11882 23468 11888 23480
rect 11940 23508 11946 23520
rect 23014 23508 23020 23520
rect 11940 23480 23020 23508
rect 11940 23468 11946 23480
rect 23014 23468 23020 23480
rect 23072 23468 23078 23520
rect 25424 23517 25452 23684
rect 25409 23511 25467 23517
rect 25409 23477 25421 23511
rect 25455 23508 25467 23511
rect 25498 23508 25504 23520
rect 25455 23480 25504 23508
rect 25455 23477 25467 23480
rect 25409 23471 25467 23477
rect 25498 23468 25504 23480
rect 25556 23468 25562 23520
rect 1104 23418 35248 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 35248 23418
rect 1104 23344 35248 23366
rect 4982 23264 4988 23316
rect 5040 23304 5046 23316
rect 5077 23307 5135 23313
rect 5077 23304 5089 23307
rect 5040 23276 5089 23304
rect 5040 23264 5046 23276
rect 5077 23273 5089 23276
rect 5123 23273 5135 23307
rect 5077 23267 5135 23273
rect 5442 23264 5448 23316
rect 5500 23264 5506 23316
rect 7098 23264 7104 23316
rect 7156 23304 7162 23316
rect 8202 23304 8208 23316
rect 7156 23276 8208 23304
rect 7156 23264 7162 23276
rect 8202 23264 8208 23276
rect 8260 23264 8266 23316
rect 13078 23264 13084 23316
rect 13136 23304 13142 23316
rect 15838 23304 15844 23316
rect 13136 23276 15844 23304
rect 13136 23264 13142 23276
rect 15838 23264 15844 23276
rect 15896 23264 15902 23316
rect 16209 23307 16267 23313
rect 16209 23273 16221 23307
rect 16255 23304 16267 23307
rect 16850 23304 16856 23316
rect 16255 23276 16856 23304
rect 16255 23273 16267 23276
rect 16209 23267 16267 23273
rect 16850 23264 16856 23276
rect 16908 23264 16914 23316
rect 20073 23307 20131 23313
rect 20073 23273 20085 23307
rect 20119 23304 20131 23307
rect 20438 23304 20444 23316
rect 20119 23276 20444 23304
rect 20119 23273 20131 23276
rect 20073 23267 20131 23273
rect 20438 23264 20444 23276
rect 20496 23264 20502 23316
rect 21637 23307 21695 23313
rect 21637 23273 21649 23307
rect 21683 23304 21695 23307
rect 21910 23304 21916 23316
rect 21683 23276 21916 23304
rect 21683 23273 21695 23276
rect 21637 23267 21695 23273
rect 21910 23264 21916 23276
rect 21968 23264 21974 23316
rect 22557 23307 22615 23313
rect 22557 23273 22569 23307
rect 22603 23304 22615 23307
rect 23014 23304 23020 23316
rect 22603 23276 23020 23304
rect 22603 23273 22615 23276
rect 22557 23267 22615 23273
rect 23014 23264 23020 23276
rect 23072 23264 23078 23316
rect 4893 23239 4951 23245
rect 4893 23205 4905 23239
rect 4939 23236 4951 23239
rect 5460 23236 5488 23264
rect 4939 23208 5488 23236
rect 12161 23239 12219 23245
rect 4939 23205 4951 23208
rect 4893 23199 4951 23205
rect 5000 23109 5028 23208
rect 12161 23205 12173 23239
rect 12207 23236 12219 23239
rect 12618 23236 12624 23248
rect 12207 23208 12624 23236
rect 12207 23205 12219 23208
rect 12161 23199 12219 23205
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 20993 23239 21051 23245
rect 14936 23208 20944 23236
rect 6822 23128 6828 23180
rect 6880 23128 6886 23180
rect 8021 23171 8079 23177
rect 8021 23137 8033 23171
rect 8067 23168 8079 23171
rect 12802 23168 12808 23180
rect 8067 23140 8616 23168
rect 8067 23137 8079 23140
rect 8021 23131 8079 23137
rect 4985 23103 5043 23109
rect 4985 23069 4997 23103
rect 5031 23069 5043 23103
rect 4985 23063 5043 23069
rect 6914 23060 6920 23112
rect 6972 23060 6978 23112
rect 7926 23060 7932 23112
rect 7984 23060 7990 23112
rect 8588 22976 8616 23140
rect 12360 23140 12808 23168
rect 9766 23060 9772 23112
rect 9824 23060 9830 23112
rect 10410 23060 10416 23112
rect 10468 23060 10474 23112
rect 12066 23060 12072 23112
rect 12124 23060 12130 23112
rect 12250 23060 12256 23112
rect 12308 23060 12314 23112
rect 12360 23109 12388 23140
rect 12802 23128 12808 23140
rect 12860 23128 12866 23180
rect 12345 23103 12403 23109
rect 12345 23069 12357 23103
rect 12391 23069 12403 23103
rect 12454 23103 12512 23109
rect 12454 23100 12466 23103
rect 12345 23063 12403 23069
rect 12452 23069 12466 23100
rect 12500 23069 12512 23103
rect 12452 23063 12512 23069
rect 12621 23103 12679 23109
rect 12621 23069 12633 23103
rect 12667 23100 12679 23103
rect 13173 23103 13231 23109
rect 13173 23100 13185 23103
rect 12667 23072 13185 23100
rect 12667 23069 12679 23072
rect 12621 23063 12679 23069
rect 13173 23069 13185 23072
rect 13219 23069 13231 23103
rect 13173 23063 13231 23069
rect 12268 23032 12296 23060
rect 12452 23032 12480 23063
rect 13354 23060 13360 23112
rect 13412 23060 13418 23112
rect 11086 23004 12204 23032
rect 12268 23004 12480 23032
rect 5626 22924 5632 22976
rect 5684 22964 5690 22976
rect 6086 22964 6092 22976
rect 5684 22936 6092 22964
rect 5684 22924 5690 22936
rect 6086 22924 6092 22936
rect 6144 22924 6150 22976
rect 8294 22924 8300 22976
rect 8352 22924 8358 22976
rect 8570 22924 8576 22976
rect 8628 22924 8634 22976
rect 12176 22964 12204 23004
rect 12710 22992 12716 23044
rect 12768 22992 12774 23044
rect 12802 22992 12808 23044
rect 12860 23032 12866 23044
rect 12897 23035 12955 23041
rect 12897 23032 12909 23035
rect 12860 23004 12909 23032
rect 12860 22992 12866 23004
rect 12897 23001 12909 23004
rect 12943 23001 12955 23035
rect 14936 23032 14964 23208
rect 15286 23128 15292 23180
rect 15344 23128 15350 23180
rect 16666 23128 16672 23180
rect 16724 23128 16730 23180
rect 19426 23128 19432 23180
rect 19484 23168 19490 23180
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 19484 23140 19717 23168
rect 19484 23128 19490 23140
rect 19705 23137 19717 23140
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 15381 23103 15439 23109
rect 15381 23069 15393 23103
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 12897 22995 12955 23001
rect 13004 23004 14964 23032
rect 13004 22964 13032 23004
rect 12176 22936 13032 22964
rect 13262 22924 13268 22976
rect 13320 22924 13326 22976
rect 14826 22924 14832 22976
rect 14884 22964 14890 22976
rect 15396 22964 15424 23063
rect 16022 23060 16028 23112
rect 16080 23060 16086 23112
rect 16485 23103 16543 23109
rect 16485 23069 16497 23103
rect 16531 23100 16543 23103
rect 16684 23100 16712 23128
rect 16531 23072 16712 23100
rect 16761 23103 16819 23109
rect 16531 23069 16543 23072
rect 16485 23063 16543 23069
rect 16761 23069 16773 23103
rect 16807 23069 16819 23103
rect 16761 23063 16819 23069
rect 19797 23103 19855 23109
rect 19797 23069 19809 23103
rect 19843 23100 19855 23103
rect 19978 23100 19984 23112
rect 19843 23072 19984 23100
rect 19843 23069 19855 23072
rect 19797 23063 19855 23069
rect 16393 23035 16451 23041
rect 16393 23032 16405 23035
rect 15764 23004 16405 23032
rect 15764 22973 15792 23004
rect 16393 23001 16405 23004
rect 16439 23032 16451 23035
rect 16776 23032 16804 23063
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20438 23060 20444 23112
rect 20496 23100 20502 23112
rect 20809 23103 20867 23109
rect 20809 23100 20821 23103
rect 20496 23072 20821 23100
rect 20496 23060 20502 23072
rect 20809 23069 20821 23072
rect 20855 23069 20867 23103
rect 20916 23100 20944 23208
rect 20993 23205 21005 23239
rect 21039 23236 21051 23239
rect 21082 23236 21088 23248
rect 21039 23208 21088 23236
rect 21039 23205 21051 23208
rect 20993 23199 21051 23205
rect 21082 23196 21088 23208
rect 21140 23236 21146 23248
rect 21453 23239 21511 23245
rect 21453 23236 21465 23239
rect 21140 23208 21465 23236
rect 21140 23196 21146 23208
rect 21453 23205 21465 23208
rect 21499 23205 21511 23239
rect 21453 23199 21511 23205
rect 21174 23128 21180 23180
rect 21232 23128 21238 23180
rect 22094 23100 22100 23112
rect 20916 23072 22100 23100
rect 20809 23063 20867 23069
rect 22094 23060 22100 23072
rect 22152 23100 22158 23112
rect 22646 23100 22652 23112
rect 22152 23072 22652 23100
rect 22152 23060 22158 23072
rect 22646 23060 22652 23072
rect 22704 23060 22710 23112
rect 33134 23060 33140 23112
rect 33192 23060 33198 23112
rect 16439 23004 16804 23032
rect 16868 23004 17264 23032
rect 16439 23001 16451 23004
rect 16393 22995 16451 23001
rect 14884 22936 15424 22964
rect 15749 22967 15807 22973
rect 14884 22924 14890 22936
rect 15749 22933 15761 22967
rect 15795 22933 15807 22967
rect 15749 22927 15807 22933
rect 15838 22924 15844 22976
rect 15896 22964 15902 22976
rect 16868 22964 16896 23004
rect 15896 22936 16896 22964
rect 15896 22924 15902 22936
rect 17126 22924 17132 22976
rect 17184 22924 17190 22976
rect 17236 22964 17264 23004
rect 20622 22992 20628 23044
rect 20680 22992 20686 23044
rect 34333 23035 34391 23041
rect 34333 23001 34345 23035
rect 34379 23032 34391 23035
rect 34882 23032 34888 23044
rect 34379 23004 34888 23032
rect 34379 23001 34391 23004
rect 34333 22995 34391 23001
rect 34882 22992 34888 23004
rect 34940 22992 34946 23044
rect 20714 22964 20720 22976
rect 17236 22936 20720 22964
rect 20714 22924 20720 22936
rect 20772 22924 20778 22976
rect 1104 22874 35236 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 35236 22874
rect 1104 22800 35236 22822
rect 5442 22720 5448 22772
rect 5500 22760 5506 22772
rect 5997 22763 6055 22769
rect 5997 22760 6009 22763
rect 5500 22732 6009 22760
rect 5500 22720 5506 22732
rect 3878 22652 3884 22704
rect 3936 22652 3942 22704
rect 5629 22695 5687 22701
rect 5629 22692 5641 22695
rect 5106 22664 5641 22692
rect 5629 22661 5641 22664
rect 5675 22661 5687 22695
rect 5629 22655 5687 22661
rect 5736 22633 5764 22732
rect 5997 22729 6009 22732
rect 6043 22729 6055 22763
rect 5997 22723 6055 22729
rect 9490 22720 9496 22772
rect 9548 22760 9554 22772
rect 10229 22763 10287 22769
rect 10229 22760 10241 22763
rect 9548 22732 10241 22760
rect 9548 22720 9554 22732
rect 10229 22729 10241 22732
rect 10275 22729 10287 22763
rect 12710 22760 12716 22772
rect 10229 22723 10287 22729
rect 12406 22732 12716 22760
rect 8846 22652 8852 22704
rect 8904 22652 8910 22704
rect 9769 22695 9827 22701
rect 9769 22661 9781 22695
rect 9815 22692 9827 22695
rect 12066 22692 12072 22704
rect 9815 22664 12072 22692
rect 9815 22661 9827 22664
rect 9769 22655 9827 22661
rect 5721 22627 5779 22633
rect 5721 22593 5733 22627
rect 5767 22593 5779 22627
rect 5721 22587 5779 22593
rect 6549 22627 6607 22633
rect 6549 22593 6561 22627
rect 6595 22624 6607 22627
rect 6822 22624 6828 22636
rect 6595 22596 6828 22624
rect 6595 22593 6607 22596
rect 6549 22587 6607 22593
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 6914 22584 6920 22636
rect 6972 22624 6978 22636
rect 7009 22627 7067 22633
rect 7009 22624 7021 22627
rect 6972 22596 7021 22624
rect 6972 22584 6978 22596
rect 7009 22593 7021 22596
rect 7055 22593 7067 22627
rect 7009 22587 7067 22593
rect 7926 22584 7932 22636
rect 7984 22584 7990 22636
rect 8570 22584 8576 22636
rect 8628 22584 8634 22636
rect 8754 22584 8760 22636
rect 8812 22624 8818 22636
rect 9784 22624 9812 22655
rect 12066 22652 12072 22664
rect 12124 22692 12130 22704
rect 12406 22692 12434 22732
rect 12710 22720 12716 22732
rect 12768 22720 12774 22772
rect 14829 22763 14887 22769
rect 14829 22729 14841 22763
rect 14875 22729 14887 22763
rect 14829 22723 14887 22729
rect 12124 22664 12434 22692
rect 14844 22692 14872 22723
rect 15010 22720 15016 22772
rect 15068 22760 15074 22772
rect 15657 22763 15715 22769
rect 15068 22732 15608 22760
rect 15068 22720 15074 22732
rect 15580 22692 15608 22732
rect 15657 22729 15669 22763
rect 15703 22760 15715 22763
rect 16022 22760 16028 22772
rect 15703 22732 16028 22760
rect 15703 22729 15715 22732
rect 15657 22723 15715 22729
rect 16022 22720 16028 22732
rect 16080 22720 16086 22772
rect 17126 22720 17132 22772
rect 17184 22720 17190 22772
rect 19334 22720 19340 22772
rect 19392 22720 19398 22772
rect 19426 22720 19432 22772
rect 19484 22720 19490 22772
rect 22649 22763 22707 22769
rect 22649 22729 22661 22763
rect 22695 22760 22707 22763
rect 23014 22760 23020 22772
rect 22695 22732 23020 22760
rect 22695 22729 22707 22732
rect 22649 22723 22707 22729
rect 14844 22664 15424 22692
rect 15580 22664 15976 22692
rect 12124 22652 12130 22664
rect 15396 22636 15424 22664
rect 8812 22596 9812 22624
rect 10505 22627 10563 22633
rect 8812 22584 8818 22596
rect 10505 22593 10517 22627
rect 10551 22624 10563 22627
rect 13354 22624 13360 22636
rect 10551 22596 13360 22624
rect 10551 22593 10563 22596
rect 10505 22587 10563 22593
rect 13354 22584 13360 22596
rect 13412 22584 13418 22636
rect 14369 22627 14427 22633
rect 14369 22593 14381 22627
rect 14415 22624 14427 22627
rect 14550 22624 14556 22636
rect 14415 22596 14556 22624
rect 14415 22593 14427 22596
rect 14369 22587 14427 22593
rect 14550 22584 14556 22596
rect 14608 22584 14614 22636
rect 14642 22584 14648 22636
rect 14700 22584 14706 22636
rect 14921 22627 14979 22633
rect 14921 22624 14933 22627
rect 14752 22596 14933 22624
rect 3602 22516 3608 22568
rect 3660 22516 3666 22568
rect 5353 22559 5411 22565
rect 5353 22525 5365 22559
rect 5399 22556 5411 22559
rect 6270 22556 6276 22568
rect 5399 22528 6276 22556
rect 5399 22525 5411 22528
rect 5353 22519 5411 22525
rect 6270 22516 6276 22528
rect 6328 22556 6334 22568
rect 6457 22559 6515 22565
rect 6457 22556 6469 22559
rect 6328 22528 6469 22556
rect 6328 22516 6334 22528
rect 6457 22525 6469 22528
rect 6503 22525 6515 22559
rect 9582 22556 9588 22568
rect 6457 22519 6515 22525
rect 9416 22528 9588 22556
rect 8294 22448 8300 22500
rect 8352 22488 8358 22500
rect 9416 22488 9444 22528
rect 9582 22516 9588 22528
rect 9640 22556 9646 22568
rect 10321 22559 10379 22565
rect 10321 22556 10333 22559
rect 9640 22528 10333 22556
rect 9640 22516 9646 22528
rect 10321 22525 10333 22528
rect 10367 22525 10379 22559
rect 10321 22519 10379 22525
rect 11974 22516 11980 22568
rect 12032 22556 12038 22568
rect 14458 22556 14464 22568
rect 12032 22528 14464 22556
rect 12032 22516 12038 22528
rect 14458 22516 14464 22528
rect 14516 22516 14522 22568
rect 8352 22460 9444 22488
rect 8352 22448 8358 22460
rect 9674 22448 9680 22500
rect 9732 22488 9738 22500
rect 9769 22491 9827 22497
rect 9769 22488 9781 22491
rect 9732 22460 9781 22488
rect 9732 22448 9738 22460
rect 9769 22457 9781 22460
rect 9815 22488 9827 22491
rect 10226 22488 10232 22500
rect 9815 22460 10232 22488
rect 9815 22457 9827 22460
rect 9769 22451 9827 22457
rect 10226 22448 10232 22460
rect 10284 22488 10290 22500
rect 12710 22488 12716 22500
rect 10284 22460 12716 22488
rect 10284 22448 10290 22460
rect 12710 22448 12716 22460
rect 12768 22448 12774 22500
rect 14752 22488 14780 22596
rect 14921 22593 14933 22596
rect 14967 22593 14979 22627
rect 15289 22627 15347 22633
rect 15289 22624 15301 22627
rect 14921 22587 14979 22593
rect 15028 22596 15301 22624
rect 14826 22516 14832 22568
rect 14884 22556 14890 22568
rect 15028 22556 15056 22596
rect 15289 22593 15301 22596
rect 15335 22593 15347 22627
rect 15289 22587 15347 22593
rect 15378 22584 15384 22636
rect 15436 22584 15442 22636
rect 15470 22584 15476 22636
rect 15528 22624 15534 22636
rect 15948 22633 15976 22664
rect 15749 22627 15807 22633
rect 15749 22624 15761 22627
rect 15528 22596 15761 22624
rect 15528 22584 15534 22596
rect 15749 22593 15761 22596
rect 15795 22593 15807 22627
rect 15749 22587 15807 22593
rect 15933 22627 15991 22633
rect 15933 22593 15945 22627
rect 15979 22593 15991 22627
rect 17144 22624 17172 22720
rect 17788 22664 18460 22692
rect 17788 22633 17816 22664
rect 18432 22633 18460 22664
rect 17773 22627 17831 22633
rect 17773 22624 17785 22627
rect 17144 22596 17785 22624
rect 15933 22587 15991 22593
rect 17773 22593 17785 22596
rect 17819 22593 17831 22627
rect 18233 22627 18291 22633
rect 18233 22624 18245 22627
rect 17773 22587 17831 22593
rect 17880 22596 18245 22624
rect 14884 22528 15056 22556
rect 14884 22516 14890 22528
rect 15102 22516 15108 22568
rect 15160 22516 15166 22568
rect 15197 22559 15255 22565
rect 15197 22525 15209 22559
rect 15243 22556 15255 22559
rect 15838 22556 15844 22568
rect 15243 22528 15844 22556
rect 15243 22525 15255 22528
rect 15197 22519 15255 22525
rect 15838 22516 15844 22528
rect 15896 22516 15902 22568
rect 17218 22516 17224 22568
rect 17276 22556 17282 22568
rect 17681 22559 17739 22565
rect 17681 22556 17693 22559
rect 17276 22528 17693 22556
rect 17276 22516 17282 22528
rect 17681 22525 17693 22528
rect 17727 22556 17739 22559
rect 17880 22556 17908 22596
rect 18233 22593 18245 22596
rect 18279 22593 18291 22627
rect 18233 22587 18291 22593
rect 18417 22627 18475 22633
rect 18417 22593 18429 22627
rect 18463 22593 18475 22627
rect 18417 22587 18475 22593
rect 18693 22627 18751 22633
rect 18693 22593 18705 22627
rect 18739 22593 18751 22627
rect 19444 22624 19472 22720
rect 19551 22627 19609 22633
rect 19551 22624 19563 22627
rect 18693 22587 18751 22593
rect 19076 22596 19563 22624
rect 17727 22528 17908 22556
rect 18141 22559 18199 22565
rect 17727 22525 17739 22528
rect 17681 22519 17739 22525
rect 18141 22525 18153 22559
rect 18187 22556 18199 22559
rect 18322 22556 18328 22568
rect 18187 22528 18328 22556
rect 18187 22525 18199 22528
rect 18141 22519 18199 22525
rect 18322 22516 18328 22528
rect 18380 22556 18386 22568
rect 18708 22556 18736 22587
rect 18380 22528 18736 22556
rect 18380 22516 18386 22528
rect 18782 22516 18788 22568
rect 18840 22516 18846 22568
rect 19076 22565 19104 22596
rect 19551 22593 19563 22596
rect 19597 22593 19609 22627
rect 19551 22587 19609 22593
rect 19705 22627 19763 22633
rect 19705 22593 19717 22627
rect 19751 22624 19763 22627
rect 19978 22624 19984 22636
rect 19751 22596 19984 22624
rect 19751 22593 19763 22596
rect 19705 22587 19763 22593
rect 19978 22584 19984 22596
rect 20036 22584 20042 22636
rect 22554 22584 22560 22636
rect 22612 22624 22618 22636
rect 22756 22633 22784 22732
rect 23014 22720 23020 22732
rect 23072 22720 23078 22772
rect 23382 22720 23388 22772
rect 23440 22720 23446 22772
rect 23845 22763 23903 22769
rect 23845 22729 23857 22763
rect 23891 22760 23903 22763
rect 24118 22760 24124 22772
rect 23891 22732 24124 22760
rect 23891 22729 23903 22732
rect 23845 22723 23903 22729
rect 22741 22627 22799 22633
rect 22741 22624 22753 22627
rect 22612 22596 22753 22624
rect 22612 22584 22618 22596
rect 22741 22593 22753 22596
rect 22787 22593 22799 22627
rect 22741 22587 22799 22593
rect 22922 22584 22928 22636
rect 22980 22584 22986 22636
rect 23198 22584 23204 22636
rect 23256 22584 23262 22636
rect 23952 22633 23980 22732
rect 24118 22720 24124 22732
rect 24176 22720 24182 22772
rect 33134 22720 33140 22772
rect 33192 22720 33198 22772
rect 25869 22695 25927 22701
rect 25869 22692 25881 22695
rect 25438 22664 25881 22692
rect 25869 22661 25881 22664
rect 25915 22661 25927 22695
rect 25869 22655 25927 22661
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22593 23995 22627
rect 23937 22587 23995 22593
rect 25498 22584 25504 22636
rect 25556 22624 25562 22636
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 25556 22596 25973 22624
rect 25556 22584 25562 22596
rect 25961 22593 25973 22596
rect 26007 22624 26019 22627
rect 26237 22627 26295 22633
rect 26237 22624 26249 22627
rect 26007 22596 26249 22624
rect 26007 22593 26019 22596
rect 25961 22587 26019 22593
rect 26237 22593 26249 22596
rect 26283 22593 26295 22627
rect 26237 22587 26295 22593
rect 19061 22559 19119 22565
rect 19061 22525 19073 22559
rect 19107 22525 19119 22559
rect 19061 22519 19119 22525
rect 24210 22516 24216 22568
rect 24268 22516 24274 22568
rect 25685 22559 25743 22565
rect 25685 22525 25697 22559
rect 25731 22556 25743 22559
rect 33152 22556 33180 22720
rect 25731 22528 33180 22556
rect 25731 22525 25743 22528
rect 25685 22519 25743 22525
rect 14384 22460 15240 22488
rect 10318 22380 10324 22432
rect 10376 22420 10382 22432
rect 14384 22429 14412 22460
rect 15212 22432 15240 22460
rect 14369 22423 14427 22429
rect 14369 22420 14381 22423
rect 10376 22392 14381 22420
rect 10376 22380 10382 22392
rect 14369 22389 14381 22392
rect 14415 22389 14427 22423
rect 14369 22383 14427 22389
rect 14550 22380 14556 22432
rect 14608 22420 14614 22432
rect 15102 22420 15108 22432
rect 14608 22392 15108 22420
rect 14608 22380 14614 22392
rect 15102 22380 15108 22392
rect 15160 22380 15166 22432
rect 15194 22380 15200 22432
rect 15252 22380 15258 22432
rect 18230 22380 18236 22432
rect 18288 22380 18294 22432
rect 1104 22330 35248 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 35248 22330
rect 1104 22256 35248 22278
rect 5810 22176 5816 22228
rect 5868 22176 5874 22228
rect 5994 22176 6000 22228
rect 6052 22176 6058 22228
rect 6914 22176 6920 22228
rect 6972 22216 6978 22228
rect 8110 22216 8116 22228
rect 6972 22188 8116 22216
rect 6972 22176 6978 22188
rect 8110 22176 8116 22188
rect 8168 22176 8174 22228
rect 9398 22176 9404 22228
rect 9456 22216 9462 22228
rect 10318 22216 10324 22228
rect 9456 22188 10324 22216
rect 9456 22176 9462 22188
rect 10318 22176 10324 22188
rect 10376 22176 10382 22228
rect 10410 22176 10416 22228
rect 10468 22176 10474 22228
rect 11517 22219 11575 22225
rect 10520 22188 11001 22216
rect 6012 22148 6040 22176
rect 6638 22148 6644 22160
rect 5552 22120 6644 22148
rect 934 21972 940 22024
rect 992 22012 998 22024
rect 5552 22021 5580 22120
rect 6638 22108 6644 22120
rect 6696 22148 6702 22160
rect 7742 22148 7748 22160
rect 6696 22120 7748 22148
rect 6696 22108 6702 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 7837 22151 7895 22157
rect 7837 22117 7849 22151
rect 7883 22148 7895 22151
rect 8202 22148 8208 22160
rect 7883 22120 8208 22148
rect 7883 22117 7895 22120
rect 7837 22111 7895 22117
rect 8202 22108 8208 22120
rect 8260 22108 8266 22160
rect 8570 22108 8576 22160
rect 8628 22148 8634 22160
rect 9125 22151 9183 22157
rect 9125 22148 9137 22151
rect 8628 22120 9137 22148
rect 8628 22108 8634 22120
rect 9125 22117 9137 22120
rect 9171 22117 9183 22151
rect 10428 22148 10456 22176
rect 9125 22111 9183 22117
rect 9232 22120 10456 22148
rect 9232 22080 9260 22120
rect 7760 22052 8064 22080
rect 1397 22015 1455 22021
rect 1397 22012 1409 22015
rect 992 21984 1409 22012
rect 992 21972 998 21984
rect 1397 21981 1409 21984
rect 1443 21981 1455 22015
rect 1397 21975 1455 21981
rect 5537 22015 5595 22021
rect 5537 21981 5549 22015
rect 5583 21981 5595 22015
rect 5537 21975 5595 21981
rect 5629 22015 5687 22021
rect 5629 21981 5641 22015
rect 5675 22012 5687 22015
rect 5902 22012 5908 22024
rect 5675 21984 5908 22012
rect 5675 21981 5687 21984
rect 5629 21975 5687 21981
rect 5902 21972 5908 21984
rect 5960 21972 5966 22024
rect 5994 21972 6000 22024
rect 6052 21972 6058 22024
rect 6178 21972 6184 22024
rect 6236 22012 6242 22024
rect 6365 22015 6423 22021
rect 6365 22012 6377 22015
rect 6236 21984 6377 22012
rect 6236 21972 6242 21984
rect 6365 21981 6377 21984
rect 6411 21981 6423 22015
rect 6365 21975 6423 21981
rect 5813 21947 5871 21953
rect 5813 21913 5825 21947
rect 5859 21944 5871 21947
rect 7760 21944 7788 22052
rect 7929 22015 7987 22021
rect 7929 21981 7941 22015
rect 7975 21981 7987 22015
rect 7929 21975 7987 21981
rect 5859 21916 7788 21944
rect 5859 21913 5871 21916
rect 5813 21907 5871 21913
rect 7944 21888 7972 21975
rect 8036 21944 8064 22052
rect 8128 22052 9260 22080
rect 8128 22024 8156 22052
rect 8110 21972 8116 22024
rect 8168 21972 8174 22024
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 22012 8355 22015
rect 8386 22012 8392 22024
rect 8343 21984 8392 22012
rect 8343 21981 8355 21984
rect 8297 21975 8355 21981
rect 8386 21972 8392 21984
rect 8444 21972 8450 22024
rect 9140 22021 9168 22052
rect 10226 22040 10232 22092
rect 10284 22040 10290 22092
rect 10520 22080 10548 22188
rect 10870 22108 10876 22160
rect 10928 22108 10934 22160
rect 10973 22148 11001 22188
rect 11517 22185 11529 22219
rect 11563 22216 11575 22219
rect 14826 22216 14832 22228
rect 11563 22188 14832 22216
rect 11563 22185 11575 22188
rect 11517 22179 11575 22185
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 15286 22176 15292 22228
rect 15344 22216 15350 22228
rect 15381 22219 15439 22225
rect 15381 22216 15393 22219
rect 15344 22188 15393 22216
rect 15344 22176 15350 22188
rect 15381 22185 15393 22188
rect 15427 22185 15439 22219
rect 15381 22179 15439 22185
rect 18138 22176 18144 22228
rect 18196 22216 18202 22228
rect 18233 22219 18291 22225
rect 18233 22216 18245 22219
rect 18196 22188 18245 22216
rect 18196 22176 18202 22188
rect 18233 22185 18245 22188
rect 18279 22185 18291 22219
rect 18233 22179 18291 22185
rect 19978 22176 19984 22228
rect 20036 22216 20042 22228
rect 20625 22219 20683 22225
rect 20625 22216 20637 22219
rect 20036 22188 20637 22216
rect 20036 22176 20042 22188
rect 20625 22185 20637 22188
rect 20671 22185 20683 22219
rect 20625 22179 20683 22185
rect 21450 22176 21456 22228
rect 21508 22176 21514 22228
rect 23293 22219 23351 22225
rect 23293 22185 23305 22219
rect 23339 22216 23351 22219
rect 24210 22216 24216 22228
rect 23339 22188 24216 22216
rect 23339 22185 23351 22188
rect 23293 22179 23351 22185
rect 24210 22176 24216 22188
rect 24268 22176 24274 22228
rect 12618 22148 12624 22160
rect 10973 22120 12624 22148
rect 12618 22108 12624 22120
rect 12676 22108 12682 22160
rect 12989 22151 13047 22157
rect 12989 22117 13001 22151
rect 13035 22148 13047 22151
rect 13035 22120 13124 22148
rect 13035 22117 13047 22120
rect 12989 22111 13047 22117
rect 13096 22092 13124 22120
rect 13262 22108 13268 22160
rect 13320 22148 13326 22160
rect 20162 22148 20168 22160
rect 13320 22120 20168 22148
rect 13320 22108 13326 22120
rect 20162 22108 20168 22120
rect 20220 22108 20226 22160
rect 20809 22151 20867 22157
rect 20809 22117 20821 22151
rect 20855 22148 20867 22151
rect 21082 22148 21088 22160
rect 20855 22120 21088 22148
rect 20855 22117 20867 22120
rect 20809 22111 20867 22117
rect 21082 22108 21088 22120
rect 21140 22108 21146 22160
rect 22189 22151 22247 22157
rect 22189 22117 22201 22151
rect 22235 22148 22247 22151
rect 22922 22148 22928 22160
rect 22235 22120 22928 22148
rect 22235 22117 22247 22120
rect 22189 22111 22247 22117
rect 22922 22108 22928 22120
rect 22980 22108 22986 22160
rect 11149 22083 11207 22089
rect 11149 22080 11161 22083
rect 10336 22052 10548 22080
rect 10704 22052 11161 22080
rect 9125 22015 9183 22021
rect 9125 21981 9137 22015
rect 9171 22012 9183 22015
rect 9493 22015 9551 22021
rect 9171 21984 9205 22012
rect 9171 21981 9183 21984
rect 9125 21975 9183 21981
rect 9493 21981 9505 22015
rect 9539 21981 9551 22015
rect 9493 21975 9551 21981
rect 8404 21944 8432 21972
rect 9508 21944 9536 21975
rect 9858 21972 9864 22024
rect 9916 21972 9922 22024
rect 10137 22015 10195 22021
rect 10137 21981 10149 22015
rect 10183 22012 10195 22015
rect 10336 22012 10364 22052
rect 10183 21984 10364 22012
rect 10413 22015 10471 22021
rect 10183 21981 10195 21984
rect 10137 21975 10195 21981
rect 10413 21981 10425 22015
rect 10459 22012 10471 22015
rect 10594 22012 10600 22024
rect 10459 21984 10600 22012
rect 10459 21981 10471 21984
rect 10413 21975 10471 21981
rect 10594 21972 10600 21984
rect 10652 21972 10658 22024
rect 8036 21916 9536 21944
rect 1578 21836 1584 21888
rect 1636 21836 1642 21888
rect 5350 21836 5356 21888
rect 5408 21836 5414 21888
rect 7926 21836 7932 21888
rect 7984 21836 7990 21888
rect 10042 21836 10048 21888
rect 10100 21876 10106 21888
rect 10597 21879 10655 21885
rect 10597 21876 10609 21879
rect 10100 21848 10609 21876
rect 10100 21836 10106 21848
rect 10597 21845 10609 21848
rect 10643 21876 10655 21879
rect 10704 21876 10732 22052
rect 10781 22015 10839 22021
rect 10781 21981 10793 22015
rect 10827 21981 10839 22015
rect 10781 21975 10839 21981
rect 10888 22006 10916 22052
rect 11149 22049 11161 22052
rect 11195 22049 11207 22083
rect 11149 22043 11207 22049
rect 12452 22052 13032 22080
rect 10965 22015 11023 22021
rect 10965 22006 10977 22015
rect 10888 21981 10977 22006
rect 11011 21981 11023 22015
rect 10888 21978 11023 21981
rect 10965 21975 11023 21978
rect 11057 22015 11115 22021
rect 11057 21981 11069 22015
rect 11103 22012 11115 22015
rect 11238 22012 11244 22024
rect 11103 21984 11244 22012
rect 11103 21981 11115 21984
rect 11057 21975 11115 21981
rect 10796 21944 10824 21975
rect 10796 21916 10916 21944
rect 10778 21876 10784 21888
rect 10643 21848 10784 21876
rect 10643 21845 10655 21848
rect 10597 21839 10655 21845
rect 10778 21836 10784 21848
rect 10836 21836 10842 21888
rect 10888 21876 10916 21916
rect 11072 21876 11100 21975
rect 11238 21972 11244 21984
rect 11296 21972 11302 22024
rect 11333 22015 11391 22021
rect 11333 21981 11345 22015
rect 11379 22012 11391 22015
rect 12452 22012 12480 22052
rect 11379 21984 12480 22012
rect 11379 21981 11391 21984
rect 11333 21975 11391 21981
rect 12526 21972 12532 22024
rect 12584 22012 12590 22024
rect 12713 22015 12771 22021
rect 12713 22012 12725 22015
rect 12584 21984 12725 22012
rect 12584 21972 12590 21984
rect 12713 21981 12725 21984
rect 12759 22012 12771 22015
rect 13004 22012 13032 22052
rect 13078 22040 13084 22092
rect 13136 22080 13142 22092
rect 20349 22083 20407 22089
rect 13136 22052 13768 22080
rect 13136 22040 13142 22052
rect 12759 21984 12940 22012
rect 13004 21984 13492 22012
rect 12759 21981 12771 21984
rect 12713 21975 12771 21981
rect 12912 21888 12940 21984
rect 12999 21947 13057 21953
rect 12999 21913 13011 21947
rect 13045 21944 13057 21947
rect 13464 21944 13492 21984
rect 13538 21972 13544 22024
rect 13596 21972 13602 22024
rect 13740 22021 13768 22052
rect 14476 22052 15056 22080
rect 14476 22024 14504 22052
rect 15028 22024 15056 22052
rect 20349 22049 20361 22083
rect 20395 22080 20407 22083
rect 20395 22052 21312 22080
rect 20395 22049 20407 22052
rect 20349 22043 20407 22049
rect 21284 22024 21312 22052
rect 21726 22040 21732 22092
rect 21784 22040 21790 22092
rect 22940 22080 22968 22108
rect 23109 22083 23167 22089
rect 23109 22080 23121 22083
rect 22940 22052 23121 22080
rect 23109 22049 23121 22052
rect 23155 22049 23167 22083
rect 23109 22043 23167 22049
rect 13725 22015 13783 22021
rect 13725 21981 13737 22015
rect 13771 21981 13783 22015
rect 13725 21975 13783 21981
rect 14458 21972 14464 22024
rect 14516 21972 14522 22024
rect 14734 21972 14740 22024
rect 14792 21972 14798 22024
rect 14918 21972 14924 22024
rect 14976 21972 14982 22024
rect 15010 21972 15016 22024
rect 15068 21972 15074 22024
rect 15102 21972 15108 22024
rect 15160 22012 15166 22024
rect 15470 22012 15476 22024
rect 15160 21984 15476 22012
rect 15160 21972 15166 21984
rect 15470 21972 15476 21984
rect 15528 21972 15534 22024
rect 16390 21972 16396 22024
rect 16448 21972 16454 22024
rect 18230 21972 18236 22024
rect 18288 21972 18294 22024
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 18417 22015 18475 22021
rect 18417 22012 18429 22015
rect 18380 21984 18429 22012
rect 18380 21972 18386 21984
rect 18417 21981 18429 21984
rect 18463 21981 18475 22015
rect 18417 21975 18475 21981
rect 18509 22015 18567 22021
rect 18509 21981 18521 22015
rect 18555 22012 18567 22015
rect 18874 22012 18880 22024
rect 18555 21984 18880 22012
rect 18555 21981 18567 21984
rect 18509 21975 18567 21981
rect 18874 21972 18880 21984
rect 18932 21972 18938 22024
rect 19889 22015 19947 22021
rect 19889 21981 19901 22015
rect 19935 22012 19947 22015
rect 19935 21984 20116 22012
rect 19935 21981 19947 21984
rect 19889 21975 19947 21981
rect 14550 21944 14556 21956
rect 13045 21916 13308 21944
rect 13464 21916 14556 21944
rect 13045 21913 13057 21916
rect 12999 21907 13057 21913
rect 13280 21888 13308 21916
rect 14550 21904 14556 21916
rect 14608 21904 14614 21956
rect 14642 21904 14648 21956
rect 14700 21944 14706 21956
rect 15120 21944 15148 21972
rect 16117 21947 16175 21953
rect 16117 21944 16129 21947
rect 14700 21916 15148 21944
rect 15948 21916 16129 21944
rect 14700 21904 14706 21916
rect 15948 21888 15976 21916
rect 16117 21913 16129 21916
rect 16163 21913 16175 21947
rect 16301 21947 16359 21953
rect 16301 21944 16313 21947
rect 16117 21907 16175 21913
rect 16224 21916 16313 21944
rect 16224 21888 16252 21916
rect 16301 21913 16313 21916
rect 16347 21913 16359 21947
rect 16301 21907 16359 21913
rect 10888 21848 11100 21876
rect 11330 21836 11336 21888
rect 11388 21876 11394 21888
rect 12802 21876 12808 21888
rect 11388 21848 12808 21876
rect 11388 21836 11394 21848
rect 12802 21836 12808 21848
rect 12860 21836 12866 21888
rect 12894 21836 12900 21888
rect 12952 21836 12958 21888
rect 13262 21836 13268 21888
rect 13320 21836 13326 21888
rect 13633 21879 13691 21885
rect 13633 21845 13645 21879
rect 13679 21876 13691 21879
rect 13814 21876 13820 21888
rect 13679 21848 13820 21876
rect 13679 21845 13691 21848
rect 13633 21839 13691 21845
rect 13814 21836 13820 21848
rect 13872 21836 13878 21888
rect 15930 21836 15936 21888
rect 15988 21836 15994 21888
rect 16206 21836 16212 21888
rect 16264 21836 16270 21888
rect 16393 21879 16451 21885
rect 16393 21845 16405 21879
rect 16439 21876 16451 21879
rect 17402 21876 17408 21888
rect 16439 21848 17408 21876
rect 16439 21845 16451 21848
rect 16393 21839 16451 21845
rect 17402 21836 17408 21848
rect 17460 21836 17466 21888
rect 19978 21836 19984 21888
rect 20036 21836 20042 21888
rect 20088 21876 20116 21984
rect 20162 21972 20168 22024
rect 20220 21972 20226 22024
rect 20993 22015 21051 22021
rect 20993 21981 21005 22015
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 20180 21944 20208 21972
rect 20441 21947 20499 21953
rect 20441 21944 20453 21947
rect 20180 21916 20453 21944
rect 20441 21913 20453 21916
rect 20487 21913 20499 21947
rect 20441 21907 20499 21913
rect 21008 21944 21036 21975
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 21821 22015 21879 22021
rect 21821 21981 21833 22015
rect 21867 22012 21879 22015
rect 23017 22015 23075 22021
rect 21867 21984 22094 22012
rect 21867 21981 21879 21984
rect 21821 21975 21879 21981
rect 21836 21944 21864 21975
rect 21008 21916 21864 21944
rect 21008 21888 21036 21916
rect 20530 21876 20536 21888
rect 20088 21848 20536 21876
rect 20530 21836 20536 21848
rect 20588 21876 20594 21888
rect 20641 21879 20699 21885
rect 20641 21876 20653 21879
rect 20588 21848 20653 21876
rect 20588 21836 20594 21848
rect 20641 21845 20653 21848
rect 20687 21845 20699 21879
rect 20641 21839 20699 21845
rect 20990 21836 20996 21888
rect 21048 21836 21054 21888
rect 22066 21876 22094 21984
rect 23017 21981 23029 22015
rect 23063 22012 23075 22015
rect 23198 22012 23204 22024
rect 23063 21984 23204 22012
rect 23063 21981 23075 21984
rect 23017 21975 23075 21981
rect 23198 21972 23204 21984
rect 23256 21972 23262 22024
rect 22462 21876 22468 21888
rect 22066 21848 22468 21876
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 1104 21786 35236 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 35236 21786
rect 1104 21712 35236 21734
rect 1578 21632 1584 21684
rect 1636 21632 1642 21684
rect 5994 21632 6000 21684
rect 6052 21672 6058 21684
rect 6457 21675 6515 21681
rect 6457 21672 6469 21675
rect 6052 21644 6469 21672
rect 6052 21632 6058 21644
rect 6457 21641 6469 21644
rect 6503 21641 6515 21675
rect 8662 21672 8668 21684
rect 6457 21635 6515 21641
rect 8220 21644 8668 21672
rect 1596 21604 1624 21632
rect 4065 21607 4123 21613
rect 4065 21604 4077 21607
rect 1596 21576 4077 21604
rect 4065 21573 4077 21576
rect 4111 21573 4123 21607
rect 4065 21567 4123 21573
rect 4798 21564 4804 21616
rect 4856 21564 4862 21616
rect 8220 21604 8248 21644
rect 8662 21632 8668 21644
rect 8720 21632 8726 21684
rect 9858 21672 9864 21684
rect 8956 21644 9864 21672
rect 8220 21576 8326 21604
rect 5626 21536 5632 21548
rect 5276 21508 5632 21536
rect 3602 21428 3608 21480
rect 3660 21468 3666 21480
rect 3789 21471 3847 21477
rect 3789 21468 3801 21471
rect 3660 21440 3801 21468
rect 3660 21428 3666 21440
rect 3789 21437 3801 21440
rect 3835 21468 3847 21471
rect 5276 21468 5304 21508
rect 5626 21496 5632 21508
rect 5684 21536 5690 21548
rect 6638 21545 6644 21548
rect 6089 21539 6147 21545
rect 6089 21536 6101 21539
rect 5684 21508 6101 21536
rect 5684 21496 5690 21508
rect 6089 21505 6101 21508
rect 6135 21505 6147 21539
rect 6632 21536 6644 21545
rect 6599 21508 6644 21536
rect 6089 21499 6147 21505
rect 6632 21499 6644 21508
rect 6638 21496 6644 21499
rect 6696 21496 6702 21548
rect 6733 21539 6791 21545
rect 6733 21505 6745 21539
rect 6779 21505 6791 21539
rect 6733 21499 6791 21505
rect 3835 21440 5304 21468
rect 3835 21437 3847 21440
rect 3789 21431 3847 21437
rect 5810 21428 5816 21480
rect 5868 21468 5874 21480
rect 6748 21468 6776 21499
rect 6914 21496 6920 21548
rect 6972 21496 6978 21548
rect 7926 21496 7932 21548
rect 7984 21496 7990 21548
rect 8665 21539 8723 21545
rect 8665 21505 8677 21539
rect 8711 21536 8723 21539
rect 8956 21536 8984 21644
rect 9858 21632 9864 21644
rect 9916 21632 9922 21684
rect 10229 21675 10287 21681
rect 10229 21641 10241 21675
rect 10275 21672 10287 21675
rect 10318 21672 10324 21684
rect 10275 21644 10324 21672
rect 10275 21641 10287 21644
rect 10229 21635 10287 21641
rect 10318 21632 10324 21644
rect 10376 21672 10382 21684
rect 11241 21675 11299 21681
rect 10376 21644 11100 21672
rect 10376 21632 10382 21644
rect 9401 21607 9459 21613
rect 9401 21573 9413 21607
rect 9447 21604 9459 21607
rect 9674 21604 9680 21616
rect 9447 21576 9680 21604
rect 9447 21573 9459 21576
rect 9401 21567 9459 21573
rect 9674 21564 9680 21576
rect 9732 21564 9738 21616
rect 9968 21576 10732 21604
rect 9968 21548 9996 21576
rect 8711 21508 8984 21536
rect 8711 21505 8723 21508
rect 8665 21499 8723 21505
rect 5868 21440 7144 21468
rect 5868 21428 5874 21440
rect 6825 21403 6883 21409
rect 6825 21369 6837 21403
rect 6871 21369 6883 21403
rect 7116 21400 7144 21440
rect 8864 21400 8892 21508
rect 9950 21496 9956 21548
rect 10008 21496 10014 21548
rect 10704 21545 10732 21576
rect 10778 21564 10784 21616
rect 10836 21604 10842 21616
rect 10873 21607 10931 21613
rect 10873 21604 10885 21607
rect 10836 21576 10885 21604
rect 10836 21564 10842 21576
rect 10873 21573 10885 21576
rect 10919 21573 10931 21607
rect 10873 21567 10931 21573
rect 11072 21545 11100 21644
rect 11241 21641 11253 21675
rect 11287 21672 11299 21675
rect 12526 21672 12532 21684
rect 11287 21644 12532 21672
rect 11287 21641 11299 21644
rect 11241 21635 11299 21641
rect 12526 21632 12532 21644
rect 12584 21632 12590 21684
rect 12636 21644 13952 21672
rect 12636 21613 12664 21644
rect 12621 21607 12679 21613
rect 12621 21573 12633 21607
rect 12667 21573 12679 21607
rect 12621 21567 12679 21573
rect 12986 21564 12992 21616
rect 13044 21604 13050 21616
rect 13044 21576 13676 21604
rect 13044 21564 13050 21576
rect 10689 21539 10747 21545
rect 10689 21505 10701 21539
rect 10735 21505 10747 21539
rect 10042 21428 10048 21480
rect 10100 21428 10106 21480
rect 10152 21477 10364 21502
rect 10689 21499 10747 21505
rect 10965 21539 11023 21545
rect 10965 21505 10977 21539
rect 11011 21505 11023 21539
rect 10965 21499 11023 21505
rect 11057 21539 11115 21545
rect 11057 21505 11069 21539
rect 11103 21505 11115 21539
rect 11057 21499 11115 21505
rect 10152 21474 10379 21477
rect 7116 21372 8892 21400
rect 6825 21363 6883 21369
rect 6840 21332 6868 21363
rect 9766 21360 9772 21412
rect 9824 21360 9830 21412
rect 9858 21360 9864 21412
rect 9916 21360 9922 21412
rect 10152 21344 10180 21474
rect 10321 21471 10379 21474
rect 10321 21437 10333 21471
rect 10367 21437 10379 21471
rect 10321 21431 10379 21437
rect 10410 21428 10416 21480
rect 10468 21428 10474 21480
rect 10597 21471 10655 21477
rect 10597 21437 10609 21471
rect 10643 21468 10655 21471
rect 10870 21468 10876 21480
rect 10643 21440 10876 21468
rect 10643 21437 10655 21440
rect 10597 21431 10655 21437
rect 10870 21428 10876 21440
rect 10928 21428 10934 21480
rect 10980 21468 11008 21499
rect 11238 21496 11244 21548
rect 11296 21496 11302 21548
rect 12713 21539 12771 21545
rect 11256 21468 11284 21496
rect 10980 21440 11284 21468
rect 8386 21332 8392 21344
rect 6840 21304 8392 21332
rect 8386 21292 8392 21304
rect 8444 21292 8450 21344
rect 10134 21292 10140 21344
rect 10192 21332 10198 21344
rect 10980 21332 11008 21440
rect 11606 21428 11612 21480
rect 11664 21468 11670 21480
rect 11793 21471 11851 21477
rect 11793 21468 11805 21471
rect 11664 21440 11805 21468
rect 11664 21428 11670 21440
rect 11793 21437 11805 21440
rect 11839 21437 11851 21471
rect 12268 21468 12296 21522
rect 12713 21505 12725 21539
rect 12759 21505 12771 21539
rect 12713 21499 12771 21505
rect 12728 21468 12756 21499
rect 12802 21496 12808 21548
rect 12860 21536 12866 21548
rect 13648 21545 13676 21576
rect 13814 21564 13820 21616
rect 13872 21564 13878 21616
rect 13633 21539 13691 21545
rect 12860 21508 13400 21536
rect 12860 21496 12866 21508
rect 12268 21440 12756 21468
rect 11793 21431 11851 21437
rect 12894 21428 12900 21480
rect 12952 21428 12958 21480
rect 13372 21477 13400 21508
rect 13633 21505 13645 21539
rect 13679 21505 13691 21539
rect 13633 21499 13691 21505
rect 13725 21539 13783 21545
rect 13725 21505 13737 21539
rect 13771 21536 13783 21539
rect 13832 21536 13860 21564
rect 13771 21508 13860 21536
rect 13771 21505 13783 21508
rect 13725 21499 13783 21505
rect 12989 21471 13047 21477
rect 12989 21437 13001 21471
rect 13035 21437 13047 21471
rect 12989 21431 13047 21437
rect 13357 21471 13415 21477
rect 13357 21437 13369 21471
rect 13403 21437 13415 21471
rect 13357 21431 13415 21437
rect 10192 21304 11008 21332
rect 12912 21332 12940 21428
rect 13004 21400 13032 21431
rect 13262 21400 13268 21412
rect 13004 21372 13268 21400
rect 13262 21360 13268 21372
rect 13320 21360 13326 21412
rect 13372 21400 13400 21431
rect 13814 21428 13820 21480
rect 13872 21428 13878 21480
rect 13924 21477 13952 21644
rect 14550 21632 14556 21684
rect 14608 21672 14614 21684
rect 16025 21675 16083 21681
rect 16025 21672 16037 21675
rect 14608 21644 16037 21672
rect 14608 21632 14614 21644
rect 16025 21641 16037 21644
rect 16071 21672 16083 21675
rect 16206 21672 16212 21684
rect 16071 21644 16212 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 16206 21632 16212 21644
rect 16264 21632 16270 21684
rect 16390 21632 16396 21684
rect 16448 21632 16454 21684
rect 16666 21632 16672 21684
rect 16724 21672 16730 21684
rect 16761 21675 16819 21681
rect 16761 21672 16773 21675
rect 16724 21644 16773 21672
rect 16724 21632 16730 21644
rect 16761 21641 16773 21644
rect 16807 21641 16819 21675
rect 16761 21635 16819 21641
rect 17402 21632 17408 21684
rect 17460 21672 17466 21684
rect 18049 21675 18107 21681
rect 18049 21672 18061 21675
rect 17460 21644 18061 21672
rect 17460 21632 17466 21644
rect 18049 21641 18061 21644
rect 18095 21641 18107 21675
rect 18049 21635 18107 21641
rect 20990 21632 20996 21684
rect 21048 21632 21054 21684
rect 21082 21632 21088 21684
rect 21140 21632 21146 21684
rect 21637 21675 21695 21681
rect 21637 21641 21649 21675
rect 21683 21672 21695 21675
rect 21726 21672 21732 21684
rect 21683 21644 21732 21672
rect 21683 21641 21695 21644
rect 21637 21635 21695 21641
rect 21726 21632 21732 21644
rect 21784 21632 21790 21684
rect 23017 21675 23075 21681
rect 23017 21641 23029 21675
rect 23063 21672 23075 21675
rect 23198 21672 23204 21684
rect 23063 21644 23204 21672
rect 23063 21641 23075 21644
rect 23017 21635 23075 21641
rect 23198 21632 23204 21644
rect 23256 21632 23262 21684
rect 15749 21607 15807 21613
rect 15749 21573 15761 21607
rect 15795 21604 15807 21607
rect 16408 21604 16436 21632
rect 17497 21607 17555 21613
rect 17497 21604 17509 21607
rect 15795 21576 16436 21604
rect 15795 21573 15807 21576
rect 15749 21567 15807 21573
rect 14182 21496 14188 21548
rect 14240 21536 14246 21548
rect 14461 21539 14519 21545
rect 14461 21536 14473 21539
rect 14240 21508 14473 21536
rect 14240 21496 14246 21508
rect 14461 21505 14473 21508
rect 14507 21505 14519 21539
rect 14461 21499 14519 21505
rect 15378 21496 15384 21548
rect 15436 21496 15442 21548
rect 15562 21496 15568 21548
rect 15620 21496 15626 21548
rect 15930 21496 15936 21548
rect 15988 21496 15994 21548
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21536 16267 21539
rect 16408 21536 16436 21576
rect 16868 21576 17509 21604
rect 16868 21548 16896 21576
rect 17497 21573 17509 21576
rect 17543 21604 17555 21607
rect 17586 21604 17592 21616
rect 17543 21576 17592 21604
rect 17543 21573 17555 21576
rect 17497 21567 17555 21573
rect 17586 21564 17592 21576
rect 17644 21564 17650 21616
rect 17697 21607 17755 21613
rect 17697 21604 17709 21607
rect 17696 21573 17709 21604
rect 17743 21573 17755 21607
rect 21100 21604 21128 21632
rect 21177 21607 21235 21613
rect 21177 21604 21189 21607
rect 21100 21576 21189 21604
rect 17696 21567 17755 21573
rect 21177 21573 21189 21576
rect 21223 21573 21235 21607
rect 21177 21567 21235 21573
rect 16255 21508 16436 21536
rect 16255 21505 16267 21508
rect 16209 21499 16267 21505
rect 16850 21496 16856 21548
rect 16908 21536 16914 21548
rect 17037 21539 17095 21545
rect 17037 21536 17049 21539
rect 16908 21508 17049 21536
rect 16908 21496 16914 21508
rect 17037 21505 17049 21508
rect 17083 21505 17095 21539
rect 17696 21536 17724 21567
rect 22462 21564 22468 21616
rect 22520 21564 22526 21616
rect 22554 21564 22560 21616
rect 22612 21564 22618 21616
rect 17957 21539 18015 21545
rect 17957 21536 17969 21539
rect 17037 21499 17095 21505
rect 17328 21508 17969 21536
rect 13909 21471 13967 21477
rect 13909 21437 13921 21471
rect 13955 21468 13967 21471
rect 14366 21468 14372 21480
rect 13955 21440 14372 21468
rect 13955 21437 13967 21440
rect 13909 21431 13967 21437
rect 14366 21428 14372 21440
rect 14424 21428 14430 21480
rect 15289 21471 15347 21477
rect 15289 21437 15301 21471
rect 15335 21468 15347 21471
rect 15654 21468 15660 21480
rect 15335 21440 15660 21468
rect 15335 21437 15347 21440
rect 15289 21431 15347 21437
rect 15654 21428 15660 21440
rect 15712 21428 15718 21480
rect 14093 21403 14151 21409
rect 13372 21372 13952 21400
rect 13924 21344 13952 21372
rect 14093 21369 14105 21403
rect 14139 21400 14151 21403
rect 15948 21400 15976 21496
rect 16393 21471 16451 21477
rect 16393 21437 16405 21471
rect 16439 21468 16451 21471
rect 16945 21471 17003 21477
rect 16945 21468 16957 21471
rect 16439 21440 16957 21468
rect 16439 21437 16451 21440
rect 16393 21431 16451 21437
rect 16945 21437 16957 21440
rect 16991 21437 17003 21471
rect 16945 21431 17003 21437
rect 14139 21372 15976 21400
rect 16960 21400 16988 21431
rect 17328 21400 17356 21508
rect 17696 21506 17740 21508
rect 17957 21505 17969 21508
rect 18003 21505 18015 21539
rect 17957 21499 18015 21505
rect 18233 21539 18291 21545
rect 18233 21505 18245 21539
rect 18279 21505 18291 21539
rect 18233 21499 18291 21505
rect 17586 21428 17592 21480
rect 17644 21468 17650 21480
rect 18248 21468 18276 21499
rect 20714 21496 20720 21548
rect 20772 21536 20778 21548
rect 20901 21539 20959 21545
rect 20901 21536 20913 21539
rect 20772 21508 20913 21536
rect 20772 21496 20778 21508
rect 20901 21505 20913 21508
rect 20947 21505 20959 21539
rect 20901 21499 20959 21505
rect 17644 21440 18276 21468
rect 17644 21428 17650 21440
rect 16960 21372 17356 21400
rect 14139 21369 14151 21372
rect 14093 21363 14151 21369
rect 17402 21360 17408 21412
rect 17460 21400 17466 21412
rect 20916 21400 20944 21499
rect 20990 21496 20996 21548
rect 21048 21536 21054 21548
rect 21085 21539 21143 21545
rect 21085 21536 21097 21539
rect 21048 21508 21097 21536
rect 21048 21496 21054 21508
rect 21085 21505 21097 21508
rect 21131 21536 21143 21539
rect 22005 21539 22063 21545
rect 22005 21536 22017 21539
rect 21131 21508 22017 21536
rect 21131 21505 21143 21508
rect 21085 21499 21143 21505
rect 22005 21505 22017 21508
rect 22051 21505 22063 21539
rect 22005 21499 22063 21505
rect 22189 21539 22247 21545
rect 22189 21505 22201 21539
rect 22235 21536 22247 21539
rect 22281 21539 22339 21545
rect 22281 21536 22293 21539
rect 22235 21508 22293 21536
rect 22235 21505 22247 21508
rect 22189 21499 22247 21505
rect 22281 21505 22293 21508
rect 22327 21505 22339 21539
rect 22572 21536 22600 21564
rect 22741 21539 22799 21545
rect 22741 21536 22753 21539
rect 22572 21508 22753 21536
rect 22281 21499 22339 21505
rect 22741 21505 22753 21508
rect 22787 21536 22799 21539
rect 23290 21536 23296 21548
rect 22787 21508 23296 21536
rect 22787 21505 22799 21508
rect 22741 21499 22799 21505
rect 23290 21496 23296 21508
rect 23348 21496 23354 21548
rect 21266 21428 21272 21480
rect 21324 21468 21330 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 21324 21440 21496 21468
rect 21324 21428 21330 21440
rect 21468 21409 21496 21440
rect 21560 21440 21833 21468
rect 21453 21403 21511 21409
rect 17460 21372 17724 21400
rect 20916 21372 21404 21400
rect 17460 21360 17466 21372
rect 13722 21332 13728 21344
rect 12912 21304 13728 21332
rect 10192 21292 10198 21304
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 13906 21292 13912 21344
rect 13964 21292 13970 21344
rect 17696 21341 17724 21372
rect 17681 21335 17739 21341
rect 17681 21301 17693 21335
rect 17727 21301 17739 21335
rect 17681 21295 17739 21301
rect 17865 21335 17923 21341
rect 17865 21301 17877 21335
rect 17911 21332 17923 21335
rect 18138 21332 18144 21344
rect 17911 21304 18144 21332
rect 17911 21301 17923 21304
rect 17865 21295 17923 21301
rect 18138 21292 18144 21304
rect 18196 21292 18202 21344
rect 18230 21292 18236 21344
rect 18288 21292 18294 21344
rect 21376 21332 21404 21372
rect 21453 21369 21465 21403
rect 21499 21369 21511 21403
rect 21453 21363 21511 21369
rect 21560 21332 21588 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 23017 21471 23075 21477
rect 23017 21437 23029 21471
rect 23063 21468 23075 21471
rect 23063 21440 23244 21468
rect 23063 21437 23075 21440
rect 23017 21431 23075 21437
rect 23216 21344 23244 21440
rect 21376 21304 21588 21332
rect 22649 21335 22707 21341
rect 22649 21301 22661 21335
rect 22695 21332 22707 21335
rect 22830 21332 22836 21344
rect 22695 21304 22836 21332
rect 22695 21301 22707 21304
rect 22649 21295 22707 21301
rect 22830 21292 22836 21304
rect 22888 21292 22894 21344
rect 23198 21292 23204 21344
rect 23256 21292 23262 21344
rect 1104 21242 35248 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 35248 21242
rect 1104 21168 35248 21190
rect 4798 21088 4804 21140
rect 4856 21128 4862 21140
rect 4893 21131 4951 21137
rect 4893 21128 4905 21131
rect 4856 21100 4905 21128
rect 4856 21088 4862 21100
rect 4893 21097 4905 21100
rect 4939 21097 4951 21131
rect 4893 21091 4951 21097
rect 5353 21131 5411 21137
rect 5353 21097 5365 21131
rect 5399 21128 5411 21131
rect 5442 21128 5448 21140
rect 5399 21100 5448 21128
rect 5399 21097 5411 21100
rect 5353 21091 5411 21097
rect 5368 21060 5396 21091
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 10137 21131 10195 21137
rect 10137 21097 10149 21131
rect 10183 21128 10195 21131
rect 10873 21131 10931 21137
rect 10183 21100 10824 21128
rect 10183 21097 10195 21100
rect 10137 21091 10195 21097
rect 4816 21032 5396 21060
rect 4816 20933 4844 21032
rect 6178 21020 6184 21072
rect 6236 21060 6242 21072
rect 6546 21060 6552 21072
rect 6236 21032 6552 21060
rect 6236 21020 6242 21032
rect 6546 21020 6552 21032
rect 6604 21020 6610 21072
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 10226 21060 10232 21072
rect 9364 21032 10232 21060
rect 9364 21020 9370 21032
rect 10226 21020 10232 21032
rect 10284 21020 10290 21072
rect 10796 21060 10824 21100
rect 10873 21097 10885 21131
rect 10919 21128 10931 21131
rect 12986 21128 12992 21140
rect 10919 21100 12992 21128
rect 10919 21097 10931 21100
rect 10873 21091 10931 21097
rect 12986 21088 12992 21100
rect 13044 21088 13050 21140
rect 13078 21088 13084 21140
rect 13136 21088 13142 21140
rect 13262 21088 13268 21140
rect 13320 21128 13326 21140
rect 13538 21128 13544 21140
rect 13320 21100 13544 21128
rect 13320 21088 13326 21100
rect 13538 21088 13544 21100
rect 13596 21088 13602 21140
rect 13725 21131 13783 21137
rect 13725 21097 13737 21131
rect 13771 21128 13783 21131
rect 13906 21128 13912 21140
rect 13771 21100 13912 21128
rect 13771 21097 13783 21100
rect 13725 21091 13783 21097
rect 13906 21088 13912 21100
rect 13964 21088 13970 21140
rect 14366 21088 14372 21140
rect 14424 21088 14430 21140
rect 14550 21088 14556 21140
rect 14608 21088 14614 21140
rect 15010 21088 15016 21140
rect 15068 21088 15074 21140
rect 15562 21088 15568 21140
rect 15620 21088 15626 21140
rect 16393 21131 16451 21137
rect 16393 21097 16405 21131
rect 16439 21128 16451 21131
rect 16850 21128 16856 21140
rect 16439 21100 16856 21128
rect 16439 21097 16451 21100
rect 16393 21091 16451 21097
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 18230 21088 18236 21140
rect 18288 21128 18294 21140
rect 18417 21131 18475 21137
rect 18417 21128 18429 21131
rect 18288 21100 18429 21128
rect 18288 21088 18294 21100
rect 18417 21097 18429 21100
rect 18463 21097 18475 21131
rect 18417 21091 18475 21097
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20257 21131 20315 21137
rect 20257 21128 20269 21131
rect 20036 21100 20269 21128
rect 20036 21088 20042 21100
rect 20257 21097 20269 21100
rect 20303 21097 20315 21131
rect 20257 21091 20315 21097
rect 20530 21088 20536 21140
rect 20588 21088 20594 21140
rect 22830 21088 22836 21140
rect 22888 21088 22894 21140
rect 24118 21088 24124 21140
rect 24176 21088 24182 21140
rect 11330 21060 11336 21072
rect 10796 21032 11336 21060
rect 11330 21020 11336 21032
rect 11388 21020 11394 21072
rect 5350 20952 5356 21004
rect 5408 20992 5414 21004
rect 7285 20995 7343 21001
rect 7285 20992 7297 20995
rect 5408 20964 7297 20992
rect 5408 20952 5414 20964
rect 7285 20961 7297 20964
rect 7331 20961 7343 20995
rect 7285 20955 7343 20961
rect 8938 20952 8944 21004
rect 8996 20992 9002 21004
rect 9490 20992 9496 21004
rect 8996 20964 9496 20992
rect 8996 20952 9002 20964
rect 9490 20952 9496 20964
rect 9548 20952 9554 21004
rect 10870 20992 10876 21004
rect 9784 20964 10364 20992
rect 9784 20936 9812 20964
rect 4801 20927 4859 20933
rect 4801 20893 4813 20927
rect 4847 20893 4859 20927
rect 4801 20887 4859 20893
rect 6270 20884 6276 20936
rect 6328 20884 6334 20936
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 7009 20927 7067 20933
rect 7009 20924 7021 20927
rect 6788 20896 7021 20924
rect 6788 20884 6794 20896
rect 7009 20893 7021 20896
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 9398 20884 9404 20936
rect 9456 20884 9462 20936
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 9861 20927 9919 20933
rect 9861 20893 9873 20927
rect 9907 20924 9919 20927
rect 9950 20924 9956 20936
rect 9907 20896 9956 20924
rect 9907 20893 9919 20896
rect 9861 20887 9919 20893
rect 5994 20816 6000 20868
rect 6052 20856 6058 20868
rect 6748 20856 6776 20884
rect 6052 20828 6776 20856
rect 6052 20816 6058 20828
rect 8662 20816 8668 20868
rect 8720 20856 8726 20868
rect 9033 20859 9091 20865
rect 9033 20856 9045 20859
rect 8720 20828 9045 20856
rect 8720 20816 8726 20828
rect 9033 20825 9045 20828
rect 9079 20825 9091 20859
rect 9033 20819 9091 20825
rect 9048 20788 9076 20819
rect 9490 20788 9496 20800
rect 9048 20760 9496 20788
rect 9490 20748 9496 20760
rect 9548 20748 9554 20800
rect 9585 20791 9643 20797
rect 9585 20757 9597 20791
rect 9631 20788 9643 20791
rect 9876 20788 9904 20887
rect 9950 20884 9956 20896
rect 10008 20884 10014 20936
rect 10134 20884 10140 20936
rect 10192 20924 10198 20936
rect 10336 20933 10364 20964
rect 10520 20964 10876 20992
rect 10520 20933 10548 20964
rect 10870 20952 10876 20964
rect 10928 20952 10934 21004
rect 10962 20952 10968 21004
rect 11020 20952 11026 21004
rect 13004 20992 13032 21088
rect 13004 20964 14320 20992
rect 10229 20927 10287 20933
rect 10229 20924 10241 20927
rect 10192 20896 10241 20924
rect 10192 20884 10198 20896
rect 10229 20893 10241 20896
rect 10275 20893 10287 20927
rect 10229 20887 10287 20893
rect 10321 20927 10379 20933
rect 10321 20893 10333 20927
rect 10367 20893 10379 20927
rect 10321 20887 10379 20893
rect 10505 20927 10563 20933
rect 10505 20893 10517 20927
rect 10551 20893 10563 20927
rect 10505 20887 10563 20893
rect 10689 20927 10747 20933
rect 10689 20893 10701 20927
rect 10735 20924 10747 20927
rect 10980 20924 11008 20952
rect 10735 20896 11008 20924
rect 13081 20927 13139 20933
rect 10735 20893 10747 20896
rect 10689 20887 10747 20893
rect 13081 20893 13093 20927
rect 13127 20924 13139 20927
rect 13262 20924 13268 20936
rect 13127 20896 13268 20924
rect 13127 20893 13139 20896
rect 13081 20887 13139 20893
rect 13262 20884 13268 20896
rect 13320 20884 13326 20936
rect 13449 20927 13507 20933
rect 13449 20893 13461 20927
rect 13495 20924 13507 20927
rect 13538 20924 13544 20936
rect 13495 20896 13544 20924
rect 13495 20893 13507 20896
rect 13449 20887 13507 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 14182 20924 14188 20936
rect 13648 20896 14188 20924
rect 10597 20859 10655 20865
rect 9968 20828 10548 20856
rect 9968 20800 9996 20828
rect 9631 20760 9904 20788
rect 9631 20757 9643 20760
rect 9585 20751 9643 20757
rect 9950 20748 9956 20800
rect 10008 20748 10014 20800
rect 10045 20791 10103 20797
rect 10045 20757 10057 20791
rect 10091 20788 10103 20791
rect 10318 20788 10324 20800
rect 10091 20760 10324 20788
rect 10091 20757 10103 20760
rect 10045 20751 10103 20757
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 10520 20788 10548 20828
rect 10597 20825 10609 20859
rect 10643 20856 10655 20859
rect 10965 20859 11023 20865
rect 10965 20856 10977 20859
rect 10643 20828 10977 20856
rect 10643 20825 10655 20828
rect 10597 20819 10655 20825
rect 10965 20825 10977 20828
rect 11011 20825 11023 20859
rect 10965 20819 11023 20825
rect 11149 20859 11207 20865
rect 11149 20825 11161 20859
rect 11195 20856 11207 20859
rect 11238 20856 11244 20868
rect 11195 20828 11244 20856
rect 11195 20825 11207 20828
rect 11149 20819 11207 20825
rect 11238 20816 11244 20828
rect 11296 20816 11302 20868
rect 11333 20859 11391 20865
rect 11333 20825 11345 20859
rect 11379 20825 11391 20859
rect 13648 20856 13676 20896
rect 14182 20884 14188 20896
rect 14240 20884 14246 20936
rect 14292 20933 14320 20964
rect 14384 20933 14412 21088
rect 14918 20952 14924 21004
rect 14976 20952 14982 21004
rect 14277 20927 14335 20933
rect 14277 20893 14289 20927
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20893 14427 20927
rect 15028 20924 15056 21088
rect 15378 20952 15384 21004
rect 15436 20952 15442 21004
rect 16022 20952 16028 21004
rect 16080 20952 16086 21004
rect 19978 20992 19984 21004
rect 19812 20964 19984 20992
rect 15289 20927 15347 20933
rect 15289 20924 15301 20927
rect 15028 20896 15301 20924
rect 14369 20887 14427 20893
rect 15289 20893 15301 20896
rect 15335 20893 15347 20927
rect 15289 20887 15347 20893
rect 15654 20884 15660 20936
rect 15712 20924 15718 20936
rect 16209 20927 16267 20933
rect 16209 20924 16221 20927
rect 15712 20896 16221 20924
rect 15712 20884 15718 20896
rect 16209 20893 16221 20896
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 17678 20884 17684 20936
rect 17736 20924 17742 20936
rect 17957 20927 18015 20933
rect 17957 20924 17969 20927
rect 17736 20896 17969 20924
rect 17736 20884 17742 20896
rect 17957 20893 17969 20896
rect 18003 20893 18015 20927
rect 17957 20887 18015 20893
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20893 18107 20927
rect 18049 20887 18107 20893
rect 13722 20865 13728 20868
rect 11333 20819 11391 20825
rect 13280 20828 13676 20856
rect 13709 20859 13728 20865
rect 11348 20788 11376 20819
rect 13280 20797 13308 20828
rect 13709 20825 13721 20859
rect 13709 20819 13728 20825
rect 13722 20816 13728 20819
rect 13780 20816 13786 20868
rect 13909 20859 13967 20865
rect 13909 20825 13921 20859
rect 13955 20825 13967 20859
rect 13909 20819 13967 20825
rect 15013 20859 15071 20865
rect 15013 20825 15025 20859
rect 15059 20825 15071 20859
rect 18064 20856 18092 20887
rect 18138 20884 18144 20936
rect 18196 20924 18202 20936
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18196 20896 18429 20924
rect 18196 20884 18202 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 19248 20905 19306 20911
rect 19248 20871 19260 20905
rect 19294 20871 19306 20905
rect 19426 20884 19432 20936
rect 19484 20924 19490 20936
rect 19812 20933 19840 20964
rect 19978 20952 19984 20964
rect 20036 20992 20042 21004
rect 22741 20995 22799 21001
rect 20036 20964 20668 20992
rect 20036 20952 20042 20964
rect 19521 20927 19579 20933
rect 19521 20924 19533 20927
rect 19484 20896 19533 20924
rect 19484 20884 19490 20896
rect 19521 20893 19533 20896
rect 19567 20893 19579 20927
rect 19521 20887 19579 20893
rect 19797 20927 19855 20933
rect 19797 20893 19809 20927
rect 19843 20893 19855 20927
rect 19797 20887 19855 20893
rect 20070 20884 20076 20936
rect 20128 20924 20134 20936
rect 20640 20933 20668 20964
rect 22741 20961 22753 20995
rect 22787 20992 22799 20995
rect 22848 20992 22876 21088
rect 22787 20964 22876 20992
rect 23201 20995 23259 21001
rect 22787 20961 22799 20964
rect 22741 20955 22799 20961
rect 23201 20961 23213 20995
rect 23247 20992 23259 20995
rect 24673 20995 24731 21001
rect 24673 20992 24685 20995
rect 23247 20964 24685 20992
rect 23247 20961 23259 20964
rect 23201 20955 23259 20961
rect 24673 20961 24685 20964
rect 24719 20961 24731 20995
rect 24673 20955 24731 20961
rect 20349 20927 20407 20933
rect 20349 20924 20361 20927
rect 20128 20896 20361 20924
rect 20128 20884 20134 20896
rect 20349 20893 20361 20896
rect 20395 20893 20407 20927
rect 20349 20887 20407 20893
rect 20625 20927 20683 20933
rect 20625 20893 20637 20927
rect 20671 20893 20683 20927
rect 20625 20887 20683 20893
rect 22833 20927 22891 20933
rect 22833 20893 22845 20927
rect 22879 20924 22891 20927
rect 22879 20896 23244 20924
rect 22879 20893 22891 20896
rect 22833 20887 22891 20893
rect 19248 20868 19306 20871
rect 15013 20819 15071 20825
rect 17972 20828 18092 20856
rect 10520 20760 11376 20788
rect 13265 20791 13323 20797
rect 13265 20757 13277 20791
rect 13311 20757 13323 20791
rect 13265 20751 13323 20757
rect 13354 20748 13360 20800
rect 13412 20788 13418 20800
rect 13924 20788 13952 20819
rect 13412 20760 13952 20788
rect 13412 20748 13418 20760
rect 13998 20748 14004 20800
rect 14056 20788 14062 20800
rect 15028 20788 15056 20819
rect 17972 20800 18000 20828
rect 19242 20816 19248 20868
rect 19300 20816 19306 20868
rect 20441 20859 20499 20865
rect 20441 20856 20453 20859
rect 19904 20828 20453 20856
rect 14056 20760 15056 20788
rect 14056 20748 14062 20760
rect 17954 20748 17960 20800
rect 18012 20748 18018 20800
rect 18601 20791 18659 20797
rect 18601 20757 18613 20791
rect 18647 20788 18659 20791
rect 19150 20788 19156 20800
rect 18647 20760 19156 20788
rect 18647 20757 18659 20760
rect 18601 20751 18659 20757
rect 19150 20748 19156 20760
rect 19208 20788 19214 20800
rect 19904 20797 19932 20828
rect 20441 20825 20453 20828
rect 20487 20825 20499 20859
rect 20441 20819 20499 20825
rect 23216 20800 23244 20896
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 24176 20896 24409 20924
rect 24176 20884 24182 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24397 20887 24455 20893
rect 33137 20927 33195 20933
rect 33137 20893 33149 20927
rect 33183 20893 33195 20927
rect 33137 20887 33195 20893
rect 25130 20816 25136 20868
rect 25188 20816 25194 20868
rect 19337 20791 19395 20797
rect 19337 20788 19349 20791
rect 19208 20760 19349 20788
rect 19208 20748 19214 20760
rect 19337 20757 19349 20760
rect 19383 20757 19395 20791
rect 19337 20751 19395 20757
rect 19705 20791 19763 20797
rect 19705 20757 19717 20791
rect 19751 20788 19763 20791
rect 19889 20791 19947 20797
rect 19889 20788 19901 20791
rect 19751 20760 19901 20788
rect 19751 20757 19763 20760
rect 19705 20751 19763 20757
rect 19889 20757 19901 20760
rect 19935 20757 19947 20791
rect 19889 20751 19947 20757
rect 23198 20748 23204 20800
rect 23256 20748 23262 20800
rect 26145 20791 26203 20797
rect 26145 20757 26157 20791
rect 26191 20788 26203 20791
rect 33152 20788 33180 20887
rect 34330 20816 34336 20868
rect 34388 20816 34394 20868
rect 26191 20760 33180 20788
rect 26191 20757 26203 20760
rect 26145 20751 26203 20757
rect 1104 20698 35236 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 35236 20698
rect 1104 20624 35236 20646
rect 9306 20544 9312 20596
rect 9364 20544 9370 20596
rect 9674 20544 9680 20596
rect 9732 20544 9738 20596
rect 9766 20544 9772 20596
rect 9824 20584 9830 20596
rect 10229 20587 10287 20593
rect 10229 20584 10241 20587
rect 9824 20556 10241 20584
rect 9824 20544 9830 20556
rect 10229 20553 10241 20556
rect 10275 20553 10287 20587
rect 10229 20547 10287 20553
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 10410 20584 10416 20596
rect 10367 20556 10416 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 8662 20516 8668 20528
rect 7958 20488 8668 20516
rect 8662 20476 8668 20488
rect 8720 20476 8726 20528
rect 8849 20519 8907 20525
rect 8849 20485 8861 20519
rect 8895 20516 8907 20519
rect 8938 20516 8944 20528
rect 8895 20488 8944 20516
rect 8895 20485 8907 20488
rect 8849 20479 8907 20485
rect 8938 20476 8944 20488
rect 8996 20476 9002 20528
rect 6825 20451 6883 20457
rect 6825 20417 6837 20451
rect 6871 20448 6883 20451
rect 7098 20448 7104 20460
rect 6871 20420 7104 20448
rect 6871 20417 6883 20420
rect 6825 20411 6883 20417
rect 7098 20408 7104 20420
rect 7156 20408 7162 20460
rect 7282 20408 7288 20460
rect 7340 20408 7346 20460
rect 9217 20451 9275 20457
rect 9217 20417 9229 20451
rect 9263 20448 9275 20451
rect 9324 20448 9352 20544
rect 9692 20516 9720 20544
rect 10336 20516 10364 20547
rect 10410 20544 10416 20556
rect 10468 20544 10474 20596
rect 10502 20544 10508 20596
rect 10560 20584 10566 20596
rect 10597 20587 10655 20593
rect 10597 20584 10609 20587
rect 10560 20556 10609 20584
rect 10560 20544 10566 20556
rect 10597 20553 10609 20556
rect 10643 20584 10655 20587
rect 12342 20584 12348 20596
rect 10643 20556 12348 20584
rect 10643 20553 10655 20556
rect 10597 20547 10655 20553
rect 9692 20488 10364 20516
rect 9263 20420 9352 20448
rect 9263 20417 9275 20420
rect 9217 20411 9275 20417
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 9824 20420 10517 20448
rect 9824 20408 9830 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 10505 20411 10563 20417
rect 8941 20383 8999 20389
rect 8941 20349 8953 20383
rect 8987 20380 8999 20383
rect 9309 20383 9367 20389
rect 8987 20352 9168 20380
rect 8987 20349 8999 20352
rect 8941 20343 8999 20349
rect 9140 20256 9168 20352
rect 9309 20349 9321 20383
rect 9355 20380 9367 20383
rect 9490 20380 9496 20392
rect 9355 20352 9496 20380
rect 9355 20349 9367 20352
rect 9309 20343 9367 20349
rect 9490 20340 9496 20352
rect 9548 20340 9554 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 9861 20383 9919 20389
rect 9861 20380 9873 20383
rect 9732 20352 9873 20380
rect 9732 20340 9738 20352
rect 9861 20349 9873 20352
rect 9907 20349 9919 20383
rect 9861 20343 9919 20349
rect 9953 20383 10011 20389
rect 9953 20349 9965 20383
rect 9999 20349 10011 20383
rect 9953 20343 10011 20349
rect 10045 20383 10103 20389
rect 10045 20349 10057 20383
rect 10091 20380 10103 20383
rect 10226 20380 10232 20392
rect 10091 20352 10232 20380
rect 10091 20349 10103 20352
rect 10045 20343 10103 20349
rect 9968 20312 9996 20343
rect 10226 20340 10232 20352
rect 10284 20380 10290 20392
rect 10612 20380 10640 20547
rect 12342 20544 12348 20556
rect 12400 20584 12406 20596
rect 14918 20584 14924 20596
rect 12400 20556 14924 20584
rect 12400 20544 12406 20556
rect 14918 20544 14924 20556
rect 14976 20544 14982 20596
rect 18230 20544 18236 20596
rect 18288 20544 18294 20596
rect 18874 20544 18880 20596
rect 18932 20544 18938 20596
rect 18969 20587 19027 20593
rect 18969 20553 18981 20587
rect 19015 20584 19027 20587
rect 19426 20584 19432 20596
rect 19015 20556 19432 20584
rect 19015 20553 19027 20556
rect 18969 20547 19027 20553
rect 19426 20544 19432 20556
rect 19484 20544 19490 20596
rect 19705 20587 19763 20593
rect 19705 20553 19717 20587
rect 19751 20584 19763 20587
rect 19978 20584 19984 20596
rect 19751 20556 19984 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 25041 20587 25099 20593
rect 25041 20553 25053 20587
rect 25087 20584 25099 20587
rect 25130 20584 25136 20596
rect 25087 20556 25136 20584
rect 25087 20553 25099 20556
rect 25041 20547 25099 20553
rect 25130 20544 25136 20556
rect 25188 20544 25194 20596
rect 25406 20544 25412 20596
rect 25464 20544 25470 20596
rect 10778 20476 10784 20528
rect 10836 20516 10842 20528
rect 12713 20519 12771 20525
rect 12713 20516 12725 20519
rect 10836 20488 12725 20516
rect 10836 20476 10842 20488
rect 12713 20485 12725 20488
rect 12759 20516 12771 20519
rect 12894 20516 12900 20528
rect 12759 20488 12900 20516
rect 12759 20485 12771 20488
rect 12713 20479 12771 20485
rect 12894 20476 12900 20488
rect 12952 20516 12958 20528
rect 15102 20516 15108 20528
rect 12952 20488 15108 20516
rect 12952 20476 12958 20488
rect 15102 20476 15108 20488
rect 15160 20476 15166 20528
rect 10689 20451 10747 20457
rect 10689 20417 10701 20451
rect 10735 20417 10747 20451
rect 10689 20411 10747 20417
rect 10284 20352 10640 20380
rect 10704 20380 10732 20411
rect 11698 20408 11704 20460
rect 11756 20448 11762 20460
rect 12529 20451 12587 20457
rect 12529 20448 12541 20451
rect 11756 20420 12541 20448
rect 11756 20408 11762 20420
rect 12529 20417 12541 20420
rect 12575 20448 12587 20451
rect 12802 20448 12808 20460
rect 12575 20420 12808 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 12802 20408 12808 20420
rect 12860 20408 12866 20460
rect 12989 20451 13047 20457
rect 12989 20417 13001 20451
rect 13035 20449 13047 20451
rect 13173 20451 13231 20457
rect 13035 20421 13124 20449
rect 13035 20417 13047 20421
rect 12989 20411 13047 20417
rect 11606 20380 11612 20392
rect 10704 20352 11612 20380
rect 10284 20340 10290 20352
rect 10704 20312 10732 20352
rect 11606 20340 11612 20352
rect 11664 20380 11670 20392
rect 13096 20380 13124 20421
rect 13173 20417 13185 20451
rect 13219 20417 13231 20451
rect 13173 20411 13231 20417
rect 15473 20451 15531 20457
rect 15473 20417 15485 20451
rect 15519 20448 15531 20451
rect 15654 20448 15660 20460
rect 15519 20420 15660 20448
rect 15519 20417 15531 20420
rect 15473 20411 15531 20417
rect 11664 20352 13124 20380
rect 11664 20340 11670 20352
rect 9968 20284 10732 20312
rect 10870 20272 10876 20324
rect 10928 20272 10934 20324
rect 12250 20312 12256 20324
rect 11992 20284 12256 20312
rect 9122 20204 9128 20256
rect 9180 20204 9186 20256
rect 9493 20247 9551 20253
rect 9493 20213 9505 20247
rect 9539 20244 9551 20247
rect 11992 20244 12020 20284
rect 12250 20272 12256 20284
rect 12308 20272 12314 20324
rect 12897 20315 12955 20321
rect 12897 20281 12909 20315
rect 12943 20312 12955 20315
rect 13188 20312 13216 20411
rect 15654 20408 15660 20420
rect 15712 20408 15718 20460
rect 15841 20451 15899 20457
rect 15841 20417 15853 20451
rect 15887 20448 15899 20451
rect 16022 20448 16028 20460
rect 15887 20420 16028 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20448 18107 20451
rect 18248 20448 18276 20544
rect 19150 20516 19156 20528
rect 19076 20488 19156 20516
rect 19076 20457 19104 20488
rect 19150 20476 19156 20488
rect 19208 20516 19214 20528
rect 19613 20519 19671 20525
rect 19613 20516 19625 20519
rect 19208 20488 19625 20516
rect 19208 20476 19214 20488
rect 19613 20485 19625 20488
rect 19659 20485 19671 20519
rect 19613 20479 19671 20485
rect 18095 20420 18276 20448
rect 19061 20451 19119 20457
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 19061 20417 19073 20451
rect 19107 20417 19119 20451
rect 19061 20411 19119 20417
rect 19429 20451 19487 20457
rect 19429 20417 19441 20451
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20349 16543 20383
rect 16485 20343 16543 20349
rect 12943 20284 13216 20312
rect 16500 20312 16528 20343
rect 17678 20340 17684 20392
rect 17736 20340 17742 20392
rect 17773 20383 17831 20389
rect 17773 20349 17785 20383
rect 17819 20380 17831 20383
rect 17954 20380 17960 20392
rect 17819 20352 17960 20380
rect 17819 20349 17831 20352
rect 17773 20343 17831 20349
rect 17954 20340 17960 20352
rect 18012 20340 18018 20392
rect 18138 20340 18144 20392
rect 18196 20340 18202 20392
rect 18601 20383 18659 20389
rect 18601 20380 18613 20383
rect 18340 20352 18613 20380
rect 18230 20312 18236 20324
rect 16500 20284 18236 20312
rect 12943 20281 12955 20284
rect 12897 20275 12955 20281
rect 9539 20216 12020 20244
rect 9539 20213 9551 20216
rect 9493 20207 9551 20213
rect 12158 20204 12164 20256
rect 12216 20244 12222 20256
rect 12912 20244 12940 20275
rect 18230 20272 18236 20284
rect 18288 20272 18294 20324
rect 18340 20321 18368 20352
rect 18601 20349 18613 20352
rect 18647 20380 18659 20383
rect 19242 20380 19248 20392
rect 18647 20352 19248 20380
rect 18647 20349 18659 20352
rect 18601 20343 18659 20349
rect 19242 20340 19248 20352
rect 19300 20380 19306 20392
rect 19444 20380 19472 20411
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 19576 20420 19717 20448
rect 19576 20408 19582 20420
rect 19705 20417 19717 20420
rect 19751 20448 19763 20451
rect 19978 20448 19984 20460
rect 19751 20420 19984 20448
rect 19751 20417 19763 20420
rect 19705 20411 19763 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 24949 20451 25007 20457
rect 24949 20417 24961 20451
rect 24995 20448 25007 20451
rect 25424 20448 25452 20544
rect 24995 20420 25452 20448
rect 24995 20417 25007 20420
rect 24949 20411 25007 20417
rect 19300 20352 19472 20380
rect 19300 20340 19306 20352
rect 18325 20315 18383 20321
rect 18325 20281 18337 20315
rect 18371 20281 18383 20315
rect 18325 20275 18383 20281
rect 12216 20216 12940 20244
rect 13173 20247 13231 20253
rect 12216 20204 12222 20216
rect 13173 20213 13185 20247
rect 13219 20244 13231 20247
rect 13354 20244 13360 20256
rect 13219 20216 13360 20244
rect 13219 20213 13231 20216
rect 13173 20207 13231 20213
rect 13354 20204 13360 20216
rect 13412 20204 13418 20256
rect 1104 20154 35248 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 35248 20154
rect 1104 20080 35248 20102
rect 6270 20000 6276 20052
rect 6328 20000 6334 20052
rect 9306 20000 9312 20052
rect 9364 20000 9370 20052
rect 9766 20000 9772 20052
rect 9824 20000 9830 20052
rect 10318 20000 10324 20052
rect 10376 20040 10382 20052
rect 10781 20043 10839 20049
rect 10781 20040 10793 20043
rect 10376 20012 10793 20040
rect 10376 20000 10382 20012
rect 10781 20009 10793 20012
rect 10827 20009 10839 20043
rect 10781 20003 10839 20009
rect 11057 20043 11115 20049
rect 11057 20009 11069 20043
rect 11103 20009 11115 20043
rect 11057 20003 11115 20009
rect 5810 19864 5816 19916
rect 5868 19904 5874 19916
rect 6288 19904 6316 20000
rect 9324 19972 9352 20000
rect 10594 19972 10600 19984
rect 9324 19944 9444 19972
rect 5868 19876 6316 19904
rect 8956 19876 9352 19904
rect 5868 19864 5874 19876
rect 8956 19848 8984 19876
rect 934 19796 940 19848
rect 992 19836 998 19848
rect 1397 19839 1455 19845
rect 1397 19836 1409 19839
rect 992 19808 1409 19836
rect 992 19796 998 19808
rect 1397 19805 1409 19808
rect 1443 19805 1455 19839
rect 1397 19799 1455 19805
rect 5721 19839 5779 19845
rect 5721 19805 5733 19839
rect 5767 19836 5779 19839
rect 5994 19836 6000 19848
rect 5767 19808 6000 19836
rect 5767 19805 5779 19808
rect 5721 19799 5779 19805
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 6086 19796 6092 19848
rect 6144 19796 6150 19848
rect 6270 19796 6276 19848
rect 6328 19796 6334 19848
rect 7098 19796 7104 19848
rect 7156 19796 7162 19848
rect 7282 19796 7288 19848
rect 7340 19836 7346 19848
rect 7469 19839 7527 19845
rect 7469 19836 7481 19839
rect 7340 19808 7481 19836
rect 7340 19796 7346 19808
rect 7469 19805 7481 19808
rect 7515 19805 7527 19839
rect 7469 19799 7527 19805
rect 8938 19796 8944 19848
rect 8996 19796 9002 19848
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9214 19836 9220 19848
rect 9171 19808 9220 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 9214 19796 9220 19808
rect 9272 19796 9278 19848
rect 9324 19845 9352 19876
rect 9416 19845 9444 19944
rect 9508 19944 10600 19972
rect 9508 19845 9536 19944
rect 10594 19932 10600 19944
rect 10652 19932 10658 19984
rect 11072 19972 11100 20003
rect 11606 20000 11612 20052
rect 11664 20000 11670 20052
rect 12710 20040 12716 20052
rect 12452 20012 12716 20040
rect 11790 19972 11796 19984
rect 11072 19944 11796 19972
rect 10137 19907 10195 19913
rect 10137 19873 10149 19907
rect 10183 19904 10195 19907
rect 10226 19904 10232 19916
rect 10183 19876 10232 19904
rect 10183 19873 10195 19876
rect 10137 19867 10195 19873
rect 10226 19864 10232 19876
rect 10284 19864 10290 19916
rect 11072 19904 11100 19944
rect 11790 19932 11796 19944
rect 11848 19972 11854 19984
rect 12452 19981 12480 20012
rect 12710 20000 12716 20012
rect 12768 20040 12774 20052
rect 12989 20043 13047 20049
rect 12989 20040 13001 20043
rect 12768 20012 13001 20040
rect 12768 20000 12774 20012
rect 12989 20009 13001 20012
rect 13035 20009 13047 20043
rect 12989 20003 13047 20009
rect 12437 19975 12495 19981
rect 12437 19972 12449 19975
rect 11848 19944 12449 19972
rect 11848 19932 11854 19944
rect 12437 19941 12449 19944
rect 12483 19941 12495 19975
rect 12437 19935 12495 19941
rect 12526 19932 12532 19984
rect 12584 19932 12590 19984
rect 12897 19975 12955 19981
rect 12897 19941 12909 19975
rect 12943 19972 12955 19975
rect 13262 19972 13268 19984
rect 12943 19944 13268 19972
rect 12943 19941 12955 19944
rect 12897 19935 12955 19941
rect 13262 19932 13268 19944
rect 13320 19972 13326 19984
rect 13320 19944 13584 19972
rect 13320 19932 13326 19944
rect 12342 19904 12348 19916
rect 10612 19876 11100 19904
rect 11532 19876 12348 19904
rect 10612 19848 10640 19876
rect 9309 19839 9367 19845
rect 9309 19805 9321 19839
rect 9355 19805 9367 19839
rect 9309 19799 9367 19805
rect 9401 19839 9459 19845
rect 9401 19805 9413 19839
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9493 19839 9551 19845
rect 9493 19805 9505 19839
rect 9539 19805 9551 19839
rect 9493 19799 9551 19805
rect 10505 19839 10563 19845
rect 10505 19805 10517 19839
rect 10551 19805 10563 19839
rect 10505 19799 10563 19805
rect 5077 19771 5135 19777
rect 5077 19737 5089 19771
rect 5123 19768 5135 19771
rect 7300 19768 7328 19796
rect 5123 19740 7328 19768
rect 8297 19771 8355 19777
rect 5123 19737 5135 19740
rect 5077 19731 5135 19737
rect 8297 19737 8309 19771
rect 8343 19768 8355 19771
rect 9508 19768 9536 19799
rect 8343 19740 9536 19768
rect 10229 19771 10287 19777
rect 8343 19737 8355 19740
rect 8297 19731 8355 19737
rect 10229 19737 10241 19771
rect 10275 19737 10287 19771
rect 10520 19768 10548 19799
rect 10594 19796 10600 19848
rect 10652 19796 10658 19848
rect 10873 19839 10931 19845
rect 10873 19805 10885 19839
rect 10919 19805 10931 19839
rect 10873 19799 10931 19805
rect 10888 19768 10916 19799
rect 11146 19796 11152 19848
rect 11204 19796 11210 19848
rect 11532 19845 11560 19876
rect 12342 19864 12348 19876
rect 12400 19864 12406 19916
rect 12802 19864 12808 19916
rect 12860 19904 12866 19916
rect 13081 19907 13139 19913
rect 13081 19904 13093 19907
rect 12860 19876 13093 19904
rect 12860 19864 12866 19876
rect 13081 19873 13093 19876
rect 13127 19873 13139 19907
rect 13081 19867 13139 19873
rect 11517 19839 11575 19845
rect 11517 19805 11529 19839
rect 11563 19805 11575 19839
rect 11974 19836 11980 19848
rect 11517 19799 11575 19805
rect 11716 19808 11980 19836
rect 11716 19768 11744 19808
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12158 19796 12164 19848
rect 12216 19796 12222 19848
rect 12618 19796 12624 19848
rect 12676 19836 12682 19848
rect 13556 19845 13584 19944
rect 16942 19932 16948 19984
rect 17000 19932 17006 19984
rect 13630 19864 13636 19916
rect 13688 19904 13694 19916
rect 14277 19907 14335 19913
rect 14277 19904 14289 19907
rect 13688 19876 14289 19904
rect 13688 19864 13694 19876
rect 14277 19873 14289 19876
rect 14323 19873 14335 19907
rect 14277 19867 14335 19873
rect 12989 19839 13047 19845
rect 12989 19836 13001 19839
rect 12676 19808 13001 19836
rect 12676 19796 12682 19808
rect 12989 19805 13001 19808
rect 13035 19805 13047 19839
rect 12989 19799 13047 19805
rect 13265 19839 13323 19845
rect 13265 19805 13277 19839
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 13725 19839 13783 19845
rect 13725 19805 13737 19839
rect 13771 19805 13783 19839
rect 13725 19799 13783 19805
rect 10520 19740 11744 19768
rect 11793 19771 11851 19777
rect 10229 19731 10287 19737
rect 11793 19737 11805 19771
rect 11839 19768 11851 19771
rect 12066 19768 12072 19780
rect 11839 19740 12072 19768
rect 11839 19737 11851 19740
rect 11793 19731 11851 19737
rect 1581 19703 1639 19709
rect 1581 19669 1593 19703
rect 1627 19700 1639 19703
rect 4614 19700 4620 19712
rect 1627 19672 4620 19700
rect 1627 19669 1639 19672
rect 1581 19663 1639 19669
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 8110 19660 8116 19712
rect 8168 19700 8174 19712
rect 9122 19700 9128 19712
rect 8168 19672 9128 19700
rect 8168 19660 8174 19672
rect 9122 19660 9128 19672
rect 9180 19700 9186 19712
rect 10244 19700 10272 19731
rect 12066 19728 12072 19740
rect 12124 19768 12130 19780
rect 13280 19768 13308 19799
rect 13740 19768 13768 19799
rect 14090 19796 14096 19848
rect 14148 19836 14154 19848
rect 14369 19839 14427 19845
rect 14369 19836 14381 19839
rect 14148 19808 14381 19836
rect 14148 19796 14154 19808
rect 14369 19805 14381 19808
rect 14415 19805 14427 19839
rect 14369 19799 14427 19805
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19836 15255 19839
rect 18046 19836 18052 19848
rect 15243 19808 18052 19836
rect 15243 19805 15255 19808
rect 15197 19799 15255 19805
rect 18046 19796 18052 19808
rect 18104 19796 18110 19848
rect 19429 19839 19487 19845
rect 19429 19836 19441 19839
rect 18248 19808 19441 19836
rect 18248 19780 18276 19808
rect 19429 19805 19441 19808
rect 19475 19805 19487 19839
rect 19429 19799 19487 19805
rect 12124 19740 13308 19768
rect 13464 19740 13768 19768
rect 16577 19771 16635 19777
rect 12124 19728 12130 19740
rect 11054 19700 11060 19712
rect 9180 19672 11060 19700
rect 9180 19660 9186 19672
rect 11054 19660 11060 19672
rect 11112 19660 11118 19712
rect 11238 19660 11244 19712
rect 11296 19700 11302 19712
rect 11333 19703 11391 19709
rect 11333 19700 11345 19703
rect 11296 19672 11345 19700
rect 11296 19660 11302 19672
rect 11333 19669 11345 19672
rect 11379 19669 11391 19703
rect 11333 19663 11391 19669
rect 11606 19660 11612 19712
rect 11664 19700 11670 19712
rect 12253 19703 12311 19709
rect 12253 19700 12265 19703
rect 11664 19672 12265 19700
rect 11664 19660 11670 19672
rect 12253 19669 12265 19672
rect 12299 19700 12311 19703
rect 12342 19700 12348 19712
rect 12299 19672 12348 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 12342 19660 12348 19672
rect 12400 19660 12406 19712
rect 13464 19709 13492 19740
rect 16577 19737 16589 19771
rect 16623 19768 16635 19771
rect 16666 19768 16672 19780
rect 16623 19740 16672 19768
rect 16623 19737 16635 19740
rect 16577 19731 16635 19737
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 18230 19728 18236 19780
rect 18288 19728 18294 19780
rect 18966 19728 18972 19780
rect 19024 19768 19030 19780
rect 19245 19771 19303 19777
rect 19245 19768 19257 19771
rect 19024 19740 19257 19768
rect 19024 19728 19030 19740
rect 19245 19737 19257 19740
rect 19291 19737 19303 19771
rect 19245 19731 19303 19737
rect 13449 19703 13507 19709
rect 13449 19669 13461 19703
rect 13495 19700 13507 19703
rect 13538 19700 13544 19712
rect 13495 19672 13544 19700
rect 13495 19669 13507 19672
rect 13449 19663 13507 19669
rect 13538 19660 13544 19672
rect 13596 19660 13602 19712
rect 17034 19660 17040 19712
rect 17092 19660 17098 19712
rect 19426 19660 19432 19712
rect 19484 19700 19490 19712
rect 19613 19703 19671 19709
rect 19613 19700 19625 19703
rect 19484 19672 19625 19700
rect 19484 19660 19490 19672
rect 19613 19669 19625 19672
rect 19659 19669 19671 19703
rect 19613 19663 19671 19669
rect 1104 19610 35236 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 35236 19610
rect 1104 19536 35236 19558
rect 5905 19499 5963 19505
rect 5905 19465 5917 19499
rect 5951 19496 5963 19499
rect 6270 19496 6276 19508
rect 5951 19468 6276 19496
rect 5951 19465 5963 19468
rect 5905 19459 5963 19465
rect 6270 19456 6276 19468
rect 6328 19496 6334 19508
rect 8110 19496 8116 19508
rect 6328 19468 8116 19496
rect 6328 19456 6334 19468
rect 8110 19456 8116 19468
rect 8168 19456 8174 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 12069 19499 12127 19505
rect 11756 19468 12020 19496
rect 11756 19456 11762 19468
rect 5721 19431 5779 19437
rect 5721 19397 5733 19431
rect 5767 19428 5779 19431
rect 5810 19428 5816 19440
rect 5767 19400 5816 19428
rect 5767 19397 5779 19400
rect 5721 19391 5779 19397
rect 5810 19388 5816 19400
rect 5868 19388 5874 19440
rect 7469 19431 7527 19437
rect 6196 19400 7144 19428
rect 3602 19320 3608 19372
rect 3660 19360 3666 19372
rect 5902 19360 5908 19372
rect 3660 19332 5908 19360
rect 3660 19320 3666 19332
rect 5902 19320 5908 19332
rect 5960 19320 5966 19372
rect 6196 19369 6224 19400
rect 6181 19363 6239 19369
rect 6181 19329 6193 19363
rect 6227 19329 6239 19363
rect 7116 19360 7144 19400
rect 7469 19397 7481 19431
rect 7515 19428 7527 19431
rect 9674 19428 9680 19440
rect 7515 19400 9680 19428
rect 7515 19397 7527 19400
rect 7469 19391 7527 19397
rect 9674 19388 9680 19400
rect 9732 19428 9738 19440
rect 10870 19428 10876 19440
rect 9732 19400 10876 19428
rect 9732 19388 9738 19400
rect 10870 19388 10876 19400
rect 10928 19388 10934 19440
rect 7653 19363 7711 19369
rect 7653 19360 7665 19363
rect 7116 19346 7665 19360
rect 7130 19332 7665 19346
rect 6181 19323 6239 19329
rect 7653 19329 7665 19332
rect 7699 19329 7711 19363
rect 7653 19323 7711 19329
rect 8018 19320 8024 19372
rect 8076 19320 8082 19372
rect 10594 19360 10600 19372
rect 9490 19334 9496 19346
rect 9445 19306 9496 19334
rect 6641 19295 6699 19301
rect 6641 19261 6653 19295
rect 6687 19261 6699 19295
rect 9490 19294 9496 19306
rect 9548 19334 9554 19346
rect 9600 19334 10600 19360
rect 9548 19332 10600 19334
rect 9548 19306 9628 19332
rect 10594 19320 10600 19332
rect 10652 19320 10658 19372
rect 11054 19320 11060 19372
rect 11112 19320 11118 19372
rect 11146 19320 11152 19372
rect 11204 19360 11210 19372
rect 11698 19360 11704 19372
rect 11204 19332 11704 19360
rect 11204 19320 11210 19332
rect 11698 19320 11704 19332
rect 11756 19350 11762 19372
rect 11992 19369 12020 19468
rect 12069 19465 12081 19499
rect 12115 19465 12127 19499
rect 12069 19459 12127 19465
rect 12084 19428 12112 19459
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 12308 19468 13768 19496
rect 12308 19456 12314 19468
rect 12618 19428 12624 19440
rect 12084 19400 12204 19428
rect 11793 19363 11851 19369
rect 11793 19350 11805 19363
rect 11756 19329 11805 19350
rect 11839 19329 11851 19363
rect 11756 19323 11851 19329
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19329 12035 19363
rect 11977 19323 12035 19329
rect 11756 19322 11836 19323
rect 11756 19320 11762 19322
rect 9548 19294 9554 19306
rect 6641 19255 6699 19261
rect 9493 19261 9505 19294
rect 9539 19261 9551 19294
rect 12176 19292 12204 19400
rect 12544 19400 12624 19428
rect 12250 19320 12256 19372
rect 12308 19320 12314 19372
rect 12342 19320 12348 19372
rect 12400 19360 12406 19372
rect 12544 19369 12572 19400
rect 12618 19388 12624 19400
rect 12676 19388 12682 19440
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 12400 19332 12449 19360
rect 12400 19320 12406 19332
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12437 19323 12495 19329
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 12710 19320 12716 19372
rect 12768 19320 12774 19372
rect 13538 19320 13544 19372
rect 13596 19320 13602 19372
rect 13740 19369 13768 19468
rect 17034 19456 17040 19508
rect 17092 19456 17098 19508
rect 17954 19456 17960 19508
rect 18012 19496 18018 19508
rect 18233 19499 18291 19505
rect 18233 19496 18245 19499
rect 18012 19468 18245 19496
rect 18012 19456 18018 19468
rect 18233 19465 18245 19468
rect 18279 19465 18291 19499
rect 18233 19459 18291 19465
rect 19978 19456 19984 19508
rect 20036 19456 20042 19508
rect 13725 19363 13783 19369
rect 13725 19329 13737 19363
rect 13771 19329 13783 19363
rect 13725 19323 13783 19329
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 15378 19360 15384 19372
rect 13955 19332 15384 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 15378 19320 15384 19332
rect 15436 19320 15442 19372
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16632 19332 16773 19360
rect 16632 19320 16638 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19360 17003 19363
rect 17052 19360 17080 19456
rect 17586 19428 17592 19440
rect 17328 19400 17592 19428
rect 17328 19369 17356 19400
rect 17586 19388 17592 19400
rect 17644 19428 17650 19440
rect 18785 19431 18843 19437
rect 17644 19400 18092 19428
rect 17644 19388 17650 19400
rect 18064 19369 18092 19400
rect 18432 19400 18736 19428
rect 16991 19332 17080 19360
rect 17313 19363 17371 19369
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17773 19363 17831 19369
rect 17773 19360 17785 19363
rect 17313 19323 17371 19329
rect 17420 19332 17785 19360
rect 12897 19295 12955 19301
rect 12176 19264 12434 19292
rect 9493 19255 9551 19261
rect 6086 19184 6092 19236
rect 6144 19224 6150 19236
rect 6454 19224 6460 19236
rect 6144 19196 6460 19224
rect 6144 19184 6150 19196
rect 6454 19184 6460 19196
rect 6512 19224 6518 19236
rect 6656 19224 6684 19255
rect 8018 19224 8024 19236
rect 6512 19196 8024 19224
rect 6512 19184 6518 19196
rect 8018 19184 8024 19196
rect 8076 19184 8082 19236
rect 12406 19224 12434 19264
rect 12897 19261 12909 19295
rect 12943 19292 12955 19295
rect 12989 19295 13047 19301
rect 12989 19292 13001 19295
rect 12943 19264 13001 19292
rect 12943 19261 12955 19264
rect 12897 19255 12955 19261
rect 12989 19261 13001 19264
rect 13035 19261 13047 19295
rect 12989 19255 13047 19261
rect 13188 19264 13584 19292
rect 12526 19224 12532 19236
rect 12406 19196 12532 19224
rect 12526 19184 12532 19196
rect 12584 19224 12590 19236
rect 12621 19227 12679 19233
rect 12621 19224 12633 19227
rect 12584 19196 12633 19224
rect 12584 19184 12590 19196
rect 12621 19193 12633 19196
rect 12667 19224 12679 19227
rect 13188 19224 13216 19264
rect 13556 19236 13584 19264
rect 17126 19252 17132 19304
rect 17184 19292 17190 19304
rect 17221 19295 17279 19301
rect 17221 19292 17233 19295
rect 17184 19264 17233 19292
rect 17184 19252 17190 19264
rect 17221 19261 17233 19264
rect 17267 19292 17279 19295
rect 17420 19292 17448 19332
rect 17773 19329 17785 19332
rect 17819 19329 17831 19363
rect 17773 19323 17831 19329
rect 17865 19363 17923 19369
rect 17865 19329 17877 19363
rect 17911 19329 17923 19363
rect 17865 19323 17923 19329
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19329 18107 19363
rect 18049 19323 18107 19329
rect 17267 19264 17448 19292
rect 17681 19295 17739 19301
rect 17267 19261 17279 19264
rect 17221 19255 17279 19261
rect 17681 19261 17693 19295
rect 17727 19292 17739 19295
rect 17880 19292 17908 19323
rect 18230 19320 18236 19372
rect 18288 19360 18294 19372
rect 18432 19369 18460 19400
rect 18417 19363 18475 19369
rect 18417 19360 18429 19363
rect 18288 19332 18429 19360
rect 18288 19320 18294 19332
rect 18417 19329 18429 19332
rect 18463 19329 18475 19363
rect 18417 19323 18475 19329
rect 18506 19320 18512 19372
rect 18564 19360 18570 19372
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 18564 19332 18613 19360
rect 18564 19320 18570 19332
rect 18601 19329 18613 19332
rect 18647 19329 18659 19363
rect 18708 19360 18736 19400
rect 18785 19397 18797 19431
rect 18831 19428 18843 19431
rect 18831 19400 19840 19428
rect 18831 19397 18843 19400
rect 18785 19391 18843 19397
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 18708 19332 19073 19360
rect 18601 19323 18659 19329
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 17727 19264 17908 19292
rect 18616 19292 18644 19323
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19521 19363 19579 19369
rect 19521 19360 19533 19363
rect 19484 19332 19533 19360
rect 19484 19320 19490 19332
rect 19521 19329 19533 19332
rect 19567 19329 19579 19363
rect 19521 19323 19579 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19360 19671 19363
rect 19702 19360 19708 19372
rect 19659 19332 19708 19360
rect 19659 19329 19671 19332
rect 19613 19323 19671 19329
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 19812 19369 19840 19400
rect 19797 19363 19855 19369
rect 19797 19329 19809 19363
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 18966 19292 18972 19304
rect 18616 19264 18972 19292
rect 17727 19261 17739 19264
rect 17681 19255 17739 19261
rect 12667 19196 13216 19224
rect 12667 19193 12679 19196
rect 12621 19187 12679 19193
rect 13262 19184 13268 19236
rect 13320 19184 13326 19236
rect 13538 19184 13544 19236
rect 13596 19184 13602 19236
rect 16758 19184 16764 19236
rect 16816 19184 16822 19236
rect 16942 19184 16948 19236
rect 17000 19224 17006 19236
rect 17037 19227 17095 19233
rect 17037 19224 17049 19227
rect 17000 19196 17049 19224
rect 17000 19184 17006 19196
rect 17037 19193 17049 19196
rect 17083 19193 17095 19227
rect 17037 19187 17095 19193
rect 17788 19168 17816 19264
rect 18966 19252 18972 19264
rect 19024 19252 19030 19304
rect 5905 19159 5963 19165
rect 5905 19125 5917 19159
rect 5951 19156 5963 19159
rect 5994 19156 6000 19168
rect 5951 19128 6000 19156
rect 5951 19125 5963 19128
rect 5905 19119 5963 19125
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 13446 19116 13452 19168
rect 13504 19116 13510 19168
rect 17770 19116 17776 19168
rect 17828 19116 17834 19168
rect 19334 19116 19340 19168
rect 19392 19116 19398 19168
rect 1104 19066 35248 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 35248 19066
rect 1104 18992 35248 19014
rect 8018 18912 8024 18964
rect 8076 18912 8082 18964
rect 8386 18912 8392 18964
rect 8444 18912 8450 18964
rect 15473 18955 15531 18961
rect 15473 18921 15485 18955
rect 15519 18952 15531 18955
rect 17126 18952 17132 18964
rect 15519 18924 17132 18952
rect 15519 18921 15531 18924
rect 15473 18915 15531 18921
rect 17126 18912 17132 18924
rect 17184 18912 17190 18964
rect 17218 18912 17224 18964
rect 17276 18912 17282 18964
rect 17678 18912 17684 18964
rect 17736 18912 17742 18964
rect 19334 18912 19340 18964
rect 19392 18912 19398 18964
rect 5258 18844 5264 18896
rect 5316 18884 5322 18896
rect 5994 18884 6000 18896
rect 5316 18856 6000 18884
rect 5316 18844 5322 18856
rect 5994 18844 6000 18856
rect 6052 18884 6058 18896
rect 6052 18856 6868 18884
rect 6052 18844 6058 18856
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 3881 18819 3939 18825
rect 3881 18816 3893 18819
rect 3660 18788 3893 18816
rect 3660 18776 3666 18788
rect 3881 18785 3893 18788
rect 3927 18785 3939 18819
rect 3881 18779 3939 18785
rect 4157 18819 4215 18825
rect 4157 18785 4169 18819
rect 4203 18816 4215 18819
rect 4798 18816 4804 18828
rect 4203 18788 4804 18816
rect 4203 18785 4215 18788
rect 4157 18779 4215 18785
rect 4798 18776 4804 18788
rect 4856 18776 4862 18828
rect 5905 18819 5963 18825
rect 5905 18785 5917 18819
rect 5951 18816 5963 18819
rect 6454 18816 6460 18828
rect 5951 18788 6460 18816
rect 5951 18785 5963 18788
rect 5905 18779 5963 18785
rect 6454 18776 6460 18788
rect 6512 18776 6518 18828
rect 5810 18708 5816 18760
rect 5868 18748 5874 18760
rect 6840 18757 6868 18856
rect 8036 18816 8064 18912
rect 7484 18788 8064 18816
rect 6641 18751 6699 18757
rect 6641 18748 6653 18751
rect 5868 18720 6653 18748
rect 5868 18708 5874 18720
rect 6641 18717 6653 18720
rect 6687 18717 6699 18751
rect 6641 18711 6699 18717
rect 6825 18751 6883 18757
rect 6825 18717 6837 18751
rect 6871 18717 6883 18751
rect 6825 18711 6883 18717
rect 7098 18708 7104 18760
rect 7156 18708 7162 18760
rect 7484 18757 7512 18788
rect 8110 18776 8116 18828
rect 8168 18776 8174 18828
rect 14369 18819 14427 18825
rect 14369 18785 14381 18819
rect 14415 18816 14427 18819
rect 14734 18816 14740 18828
rect 14415 18788 14740 18816
rect 14415 18785 14427 18788
rect 14369 18779 14427 18785
rect 14734 18776 14740 18788
rect 14792 18776 14798 18828
rect 16942 18776 16948 18828
rect 17000 18776 17006 18828
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 7558 18708 7564 18760
rect 7616 18708 7622 18760
rect 7892 18751 7950 18757
rect 7892 18748 7904 18751
rect 7668 18720 7904 18748
rect 4890 18640 4896 18692
rect 4948 18640 4954 18692
rect 6273 18683 6331 18689
rect 6273 18649 6285 18683
rect 6319 18680 6331 18683
rect 7006 18680 7012 18692
rect 6319 18652 7012 18680
rect 6319 18649 6331 18652
rect 6273 18643 6331 18649
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 7116 18680 7144 18708
rect 7668 18680 7696 18720
rect 7892 18717 7904 18720
rect 7938 18717 7950 18751
rect 7892 18711 7950 18717
rect 7116 18652 7696 18680
rect 7742 18640 7748 18692
rect 7800 18640 7806 18692
rect 7558 18572 7564 18624
rect 7616 18612 7622 18624
rect 8128 18612 8156 18776
rect 15013 18751 15071 18757
rect 15013 18748 15025 18751
rect 14476 18720 15025 18748
rect 14476 18624 14504 18720
rect 15013 18717 15025 18720
rect 15059 18717 15071 18751
rect 15013 18711 15071 18717
rect 15028 18680 15056 18711
rect 15286 18708 15292 18760
rect 15344 18748 15350 18760
rect 15841 18751 15899 18757
rect 15841 18748 15853 18751
rect 15344 18720 15853 18748
rect 15344 18708 15350 18720
rect 15841 18717 15853 18720
rect 15887 18717 15899 18751
rect 15841 18711 15899 18717
rect 16666 18708 16672 18760
rect 16724 18748 16730 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16724 18720 16865 18748
rect 16724 18708 16730 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 15565 18683 15623 18689
rect 15565 18680 15577 18683
rect 15028 18652 15577 18680
rect 15565 18649 15577 18652
rect 15611 18649 15623 18683
rect 15565 18643 15623 18649
rect 15749 18683 15807 18689
rect 15749 18649 15761 18683
rect 15795 18649 15807 18683
rect 17144 18680 17172 18912
rect 17586 18844 17592 18896
rect 17644 18844 17650 18896
rect 17604 18748 17632 18844
rect 19352 18816 19380 18912
rect 20073 18887 20131 18893
rect 20073 18853 20085 18887
rect 20119 18884 20131 18887
rect 20119 18856 20576 18884
rect 20119 18853 20131 18856
rect 20073 18847 20131 18853
rect 20548 18825 20576 18856
rect 20990 18844 20996 18896
rect 21048 18844 21054 18896
rect 19613 18819 19671 18825
rect 19613 18816 19625 18819
rect 19352 18788 19625 18816
rect 19613 18785 19625 18788
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 20533 18819 20591 18825
rect 20533 18785 20545 18819
rect 20579 18816 20591 18819
rect 20714 18816 20720 18828
rect 20579 18788 20720 18816
rect 20579 18785 20591 18788
rect 20533 18779 20591 18785
rect 20714 18776 20720 18788
rect 20772 18776 20778 18828
rect 17862 18748 17868 18760
rect 17604 18720 17868 18748
rect 17862 18708 17868 18720
rect 17920 18708 17926 18760
rect 19334 18708 19340 18760
rect 19392 18748 19398 18760
rect 19702 18748 19708 18760
rect 19392 18720 19708 18748
rect 19392 18708 19398 18720
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18748 20683 18751
rect 20806 18748 20812 18760
rect 20671 18720 20812 18748
rect 20671 18717 20683 18720
rect 20625 18711 20683 18717
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 33134 18708 33140 18760
rect 33192 18708 33198 18760
rect 17589 18683 17647 18689
rect 17589 18680 17601 18683
rect 17144 18652 17601 18680
rect 15749 18643 15807 18649
rect 17589 18649 17601 18652
rect 17635 18649 17647 18683
rect 17589 18643 17647 18649
rect 7616 18584 8156 18612
rect 7616 18572 7622 18584
rect 10318 18572 10324 18624
rect 10376 18612 10382 18624
rect 12618 18612 12624 18624
rect 10376 18584 12624 18612
rect 10376 18572 10382 18584
rect 12618 18572 12624 18584
rect 12676 18572 12682 18624
rect 12986 18572 12992 18624
rect 13044 18612 13050 18624
rect 13630 18612 13636 18624
rect 13044 18584 13636 18612
rect 13044 18572 13050 18584
rect 13630 18572 13636 18584
rect 13688 18572 13694 18624
rect 14458 18572 14464 18624
rect 14516 18572 14522 18624
rect 14550 18572 14556 18624
rect 14608 18612 14614 18624
rect 15105 18615 15163 18621
rect 15105 18612 15117 18615
rect 14608 18584 15117 18612
rect 14608 18572 14614 18584
rect 15105 18581 15117 18584
rect 15151 18612 15163 18615
rect 15764 18612 15792 18643
rect 17770 18640 17776 18692
rect 17828 18640 17834 18692
rect 34333 18683 34391 18689
rect 34333 18649 34345 18683
rect 34379 18680 34391 18683
rect 34882 18680 34888 18692
rect 34379 18652 34888 18680
rect 34379 18649 34391 18652
rect 34333 18643 34391 18649
rect 34882 18640 34888 18652
rect 34940 18640 34946 18692
rect 15151 18584 15792 18612
rect 15841 18615 15899 18621
rect 15151 18581 15163 18584
rect 15105 18575 15163 18581
rect 15841 18581 15853 18615
rect 15887 18612 15899 18615
rect 17788 18612 17816 18640
rect 15887 18584 17816 18612
rect 15887 18581 15899 18584
rect 15841 18575 15899 18581
rect 1104 18522 35236 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 35236 18522
rect 1104 18448 35236 18470
rect 4890 18368 4896 18420
rect 4948 18408 4954 18420
rect 4985 18411 5043 18417
rect 4985 18408 4997 18411
rect 4948 18380 4997 18408
rect 4948 18368 4954 18380
rect 4985 18377 4997 18380
rect 5031 18377 5043 18411
rect 4985 18371 5043 18377
rect 5442 18368 5448 18420
rect 5500 18368 5506 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 5997 18411 6055 18417
rect 5997 18408 6009 18411
rect 5960 18380 6009 18408
rect 5960 18368 5966 18380
rect 5997 18377 6009 18380
rect 6043 18377 6055 18411
rect 7742 18408 7748 18420
rect 5997 18371 6055 18377
rect 7024 18380 7748 18408
rect 4893 18275 4951 18281
rect 4893 18241 4905 18275
rect 4939 18272 4951 18275
rect 5460 18272 5488 18368
rect 7024 18340 7052 18380
rect 7742 18368 7748 18380
rect 7800 18368 7806 18420
rect 9398 18408 9404 18420
rect 8312 18380 9404 18408
rect 8312 18349 8340 18380
rect 9398 18368 9404 18380
rect 9456 18408 9462 18420
rect 12986 18408 12992 18420
rect 9456 18380 12992 18408
rect 9456 18368 9462 18380
rect 12986 18368 12992 18380
rect 13044 18368 13050 18420
rect 13096 18380 14228 18408
rect 13096 18349 13124 18380
rect 6932 18312 7052 18340
rect 8297 18343 8355 18349
rect 6932 18281 6960 18312
rect 8297 18309 8309 18343
rect 8343 18309 8355 18343
rect 10045 18343 10103 18349
rect 8297 18303 8355 18309
rect 8864 18312 9720 18340
rect 4939 18244 5488 18272
rect 6917 18275 6975 18281
rect 4939 18241 4951 18244
rect 4893 18235 4951 18241
rect 6917 18241 6929 18275
rect 6963 18241 6975 18275
rect 6917 18235 6975 18241
rect 7006 18232 7012 18284
rect 7064 18272 7070 18284
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 7064 18244 7481 18272
rect 7064 18232 7070 18244
rect 7469 18241 7481 18244
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 8864 18204 8892 18312
rect 8938 18232 8944 18284
rect 8996 18272 9002 18284
rect 9692 18281 9720 18312
rect 10045 18309 10057 18343
rect 10091 18340 10103 18343
rect 13081 18343 13139 18349
rect 13081 18340 13093 18343
rect 10091 18312 13093 18340
rect 10091 18309 10103 18312
rect 10045 18303 10103 18309
rect 13081 18309 13093 18312
rect 13127 18309 13139 18343
rect 14093 18343 14151 18349
rect 14093 18340 14105 18343
rect 13081 18303 13139 18309
rect 13556 18312 14105 18340
rect 9493 18275 9551 18281
rect 9493 18272 9505 18275
rect 8996 18244 9505 18272
rect 8996 18232 9002 18244
rect 9493 18241 9505 18244
rect 9539 18241 9551 18275
rect 9493 18235 9551 18241
rect 9677 18275 9735 18281
rect 9677 18241 9689 18275
rect 9723 18241 9735 18275
rect 9677 18235 9735 18241
rect 10597 18275 10655 18281
rect 10597 18241 10609 18275
rect 10643 18272 10655 18275
rect 10962 18272 10968 18284
rect 10643 18244 10968 18272
rect 10643 18241 10655 18244
rect 10597 18235 10655 18241
rect 9030 18204 9036 18216
rect 8864 18176 9036 18204
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 9508 18204 9536 18235
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18272 11391 18275
rect 11379 18244 12512 18272
rect 11379 18241 11391 18244
rect 11333 18235 11391 18241
rect 9858 18204 9864 18216
rect 9508 18176 9864 18204
rect 9858 18164 9864 18176
rect 9916 18164 9922 18216
rect 10686 18164 10692 18216
rect 10744 18164 10750 18216
rect 12484 18204 12512 18244
rect 12618 18232 12624 18284
rect 12676 18232 12682 18284
rect 12805 18275 12863 18281
rect 12805 18241 12817 18275
rect 12851 18241 12863 18275
rect 12805 18235 12863 18241
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18272 13231 18275
rect 13262 18272 13268 18284
rect 13219 18244 13268 18272
rect 13219 18241 13231 18244
rect 13173 18235 13231 18241
rect 12820 18204 12848 18235
rect 13262 18232 13268 18244
rect 13320 18272 13326 18284
rect 13556 18281 13584 18312
rect 14093 18309 14105 18312
rect 14139 18309 14151 18343
rect 14200 18340 14228 18380
rect 14458 18368 14464 18420
rect 14516 18368 14522 18420
rect 14550 18368 14556 18420
rect 14608 18368 14614 18420
rect 15194 18368 15200 18420
rect 15252 18368 15258 18420
rect 15933 18411 15991 18417
rect 15304 18380 15700 18408
rect 14568 18340 14596 18368
rect 15304 18340 15332 18380
rect 15672 18340 15700 18380
rect 15933 18377 15945 18411
rect 15979 18408 15991 18411
rect 16574 18408 16580 18420
rect 15979 18380 16580 18408
rect 15979 18377 15991 18380
rect 15933 18371 15991 18377
rect 16574 18368 16580 18380
rect 16632 18368 16638 18420
rect 17862 18368 17868 18420
rect 17920 18368 17926 18420
rect 16209 18343 16267 18349
rect 16209 18340 16221 18343
rect 14200 18312 14596 18340
rect 14752 18312 15332 18340
rect 14093 18303 14151 18309
rect 14752 18284 14780 18312
rect 13541 18275 13599 18281
rect 13541 18272 13553 18275
rect 13320 18244 13553 18272
rect 13320 18232 13326 18244
rect 13541 18241 13553 18244
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 14001 18275 14059 18281
rect 14001 18241 14013 18275
rect 14047 18241 14059 18275
rect 14277 18275 14335 18281
rect 14277 18272 14289 18275
rect 14001 18235 14059 18241
rect 14108 18244 14289 18272
rect 13449 18207 13507 18213
rect 13449 18204 13461 18207
rect 12484 18176 13461 18204
rect 13449 18173 13461 18176
rect 13495 18204 13507 18207
rect 14016 18204 14044 18235
rect 13495 18176 14044 18204
rect 13495 18173 13507 18176
rect 13449 18167 13507 18173
rect 9309 18139 9367 18145
rect 9309 18105 9321 18139
rect 9355 18136 9367 18139
rect 9766 18136 9772 18148
rect 9355 18108 9772 18136
rect 9355 18105 9367 18108
rect 9309 18099 9367 18105
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 9953 18139 10011 18145
rect 9953 18105 9965 18139
rect 9999 18136 10011 18139
rect 9999 18108 11100 18136
rect 9999 18105 10011 18108
rect 9953 18099 10011 18105
rect 11072 18068 11100 18108
rect 12618 18096 12624 18148
rect 12676 18136 12682 18148
rect 14108 18136 14136 18244
rect 14277 18241 14289 18244
rect 14323 18241 14335 18275
rect 14277 18235 14335 18241
rect 14458 18232 14464 18284
rect 14516 18272 14522 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14516 18244 14565 18272
rect 14516 18232 14522 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 14734 18232 14740 18284
rect 14792 18232 14798 18284
rect 14826 18232 14832 18284
rect 14884 18232 14890 18284
rect 14921 18275 14979 18281
rect 14921 18241 14933 18275
rect 14967 18272 14979 18275
rect 15102 18272 15108 18284
rect 14967 18244 15108 18272
rect 14967 18241 14979 18244
rect 14921 18235 14979 18241
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 15304 18281 15332 18312
rect 15396 18312 15608 18340
rect 15672 18312 16221 18340
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18241 15347 18275
rect 15289 18235 15347 18241
rect 15396 18204 15424 18312
rect 15580 18284 15608 18312
rect 16209 18309 16221 18312
rect 16255 18309 16267 18343
rect 16209 18303 16267 18309
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 14476 18176 15424 18204
rect 12676 18108 14136 18136
rect 12676 18096 12682 18108
rect 14274 18096 14280 18148
rect 14332 18136 14338 18148
rect 14476 18136 14504 18176
rect 14332 18108 14504 18136
rect 14332 18096 14338 18108
rect 14550 18096 14556 18148
rect 14608 18136 14614 18148
rect 15488 18136 15516 18235
rect 15562 18232 15568 18284
rect 15620 18232 15626 18284
rect 15654 18232 15660 18284
rect 15712 18272 15718 18284
rect 17037 18275 17095 18281
rect 17037 18272 17049 18275
rect 15712 18244 17049 18272
rect 15712 18232 15718 18244
rect 17037 18241 17049 18244
rect 17083 18272 17095 18275
rect 17497 18275 17555 18281
rect 17497 18272 17509 18275
rect 17083 18244 17509 18272
rect 17083 18241 17095 18244
rect 17037 18235 17095 18241
rect 17497 18241 17509 18244
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 17681 18275 17739 18281
rect 17681 18241 17693 18275
rect 17727 18241 17739 18275
rect 17681 18235 17739 18241
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 14608 18108 15516 18136
rect 16224 18176 16957 18204
rect 14608 18096 14614 18108
rect 13814 18068 13820 18080
rect 11072 18040 13820 18068
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 16224 18068 16252 18176
rect 16945 18173 16957 18176
rect 16991 18204 17003 18207
rect 17696 18204 17724 18235
rect 16991 18176 17724 18204
rect 16991 18173 17003 18176
rect 16945 18167 17003 18173
rect 17405 18139 17463 18145
rect 17405 18105 17417 18139
rect 17451 18136 17463 18139
rect 18506 18136 18512 18148
rect 17451 18108 18512 18136
rect 17451 18105 17463 18108
rect 17405 18099 17463 18105
rect 18506 18096 18512 18108
rect 18564 18096 18570 18148
rect 13955 18040 16252 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 1104 17978 35248 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 35248 17978
rect 1104 17904 35248 17926
rect 5902 17824 5908 17876
rect 5960 17864 5966 17876
rect 6181 17867 6239 17873
rect 6181 17864 6193 17867
rect 5960 17836 6193 17864
rect 5960 17824 5966 17836
rect 6181 17833 6193 17836
rect 6227 17833 6239 17867
rect 6181 17827 6239 17833
rect 10597 17867 10655 17873
rect 10597 17833 10609 17867
rect 10643 17864 10655 17867
rect 10686 17864 10692 17876
rect 10643 17836 10692 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 10686 17824 10692 17836
rect 10744 17824 10750 17876
rect 10962 17824 10968 17876
rect 11020 17824 11026 17876
rect 14645 17867 14703 17873
rect 14645 17833 14657 17867
rect 14691 17864 14703 17867
rect 15286 17864 15292 17876
rect 14691 17836 15292 17864
rect 14691 17833 14703 17836
rect 14645 17827 14703 17833
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 18693 17867 18751 17873
rect 18693 17833 18705 17867
rect 18739 17864 18751 17867
rect 19334 17864 19340 17876
rect 18739 17836 19340 17864
rect 18739 17833 18751 17836
rect 18693 17827 18751 17833
rect 19334 17824 19340 17836
rect 19392 17824 19398 17876
rect 20070 17824 20076 17876
rect 20128 17824 20134 17876
rect 20806 17824 20812 17876
rect 20864 17824 20870 17876
rect 23198 17824 23204 17876
rect 23256 17824 23262 17876
rect 24118 17824 24124 17876
rect 24176 17824 24182 17876
rect 9861 17799 9919 17805
rect 9861 17765 9873 17799
rect 9907 17765 9919 17799
rect 9861 17759 9919 17765
rect 3602 17688 3608 17740
rect 3660 17728 3666 17740
rect 3881 17731 3939 17737
rect 3881 17728 3893 17731
rect 3660 17700 3893 17728
rect 3660 17688 3666 17700
rect 3881 17697 3893 17700
rect 3927 17697 3939 17731
rect 9876 17728 9904 17759
rect 10318 17756 10324 17808
rect 10376 17756 10382 17808
rect 12529 17799 12587 17805
rect 10428 17768 11192 17796
rect 9876 17700 10364 17728
rect 3881 17691 3939 17697
rect 934 17620 940 17672
rect 992 17660 998 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 992 17632 1409 17660
rect 992 17620 998 17632
rect 1397 17629 1409 17632
rect 1443 17629 1455 17663
rect 1397 17623 1455 17629
rect 7006 17620 7012 17672
rect 7064 17620 7070 17672
rect 7392 17660 7512 17670
rect 7742 17660 7748 17672
rect 7116 17642 7748 17660
rect 7116 17632 7420 17642
rect 7484 17632 7748 17642
rect 4157 17595 4215 17601
rect 4157 17592 4169 17595
rect 1596 17564 4169 17592
rect 1596 17533 1624 17564
rect 4157 17561 4169 17564
rect 4203 17561 4215 17595
rect 4157 17555 4215 17561
rect 4890 17552 4896 17604
rect 4948 17552 4954 17604
rect 5905 17595 5963 17601
rect 5905 17561 5917 17595
rect 5951 17592 5963 17595
rect 7116 17592 7144 17632
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 9214 17660 9220 17672
rect 7944 17632 9220 17660
rect 5951 17564 7144 17592
rect 7944 17578 7972 17632
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 9677 17663 9735 17669
rect 9677 17629 9689 17663
rect 9723 17629 9735 17663
rect 9677 17623 9735 17629
rect 5951 17561 5963 17564
rect 5905 17555 5963 17561
rect 8938 17552 8944 17604
rect 8996 17552 9002 17604
rect 9125 17595 9183 17601
rect 9125 17561 9137 17595
rect 9171 17592 9183 17595
rect 9493 17595 9551 17601
rect 9171 17564 9444 17592
rect 9171 17561 9183 17564
rect 9125 17555 9183 17561
rect 9416 17536 9444 17564
rect 9493 17561 9505 17595
rect 9539 17592 9551 17595
rect 9692 17592 9720 17623
rect 9766 17620 9772 17672
rect 9824 17620 9830 17672
rect 10336 17669 10364 17700
rect 9861 17663 9919 17669
rect 9861 17629 9873 17663
rect 9907 17660 9919 17663
rect 10321 17663 10379 17669
rect 9907 17632 10272 17660
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 9539 17564 9720 17592
rect 9784 17592 9812 17620
rect 10244 17604 10272 17632
rect 10321 17629 10333 17663
rect 10367 17629 10379 17663
rect 10321 17623 10379 17629
rect 9953 17595 10011 17601
rect 9953 17592 9965 17595
rect 9784 17564 9965 17592
rect 9539 17561 9551 17564
rect 9493 17555 9551 17561
rect 1581 17527 1639 17533
rect 1581 17493 1593 17527
rect 1627 17493 1639 17527
rect 1581 17487 1639 17493
rect 9030 17484 9036 17536
rect 9088 17524 9094 17536
rect 9217 17527 9275 17533
rect 9217 17524 9229 17527
rect 9088 17496 9229 17524
rect 9088 17484 9094 17496
rect 9217 17493 9229 17496
rect 9263 17493 9275 17527
rect 9217 17487 9275 17493
rect 9306 17484 9312 17536
rect 9364 17484 9370 17536
rect 9398 17484 9404 17536
rect 9456 17524 9462 17536
rect 9582 17524 9588 17536
rect 9456 17496 9588 17524
rect 9456 17484 9462 17496
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 9692 17524 9720 17564
rect 9953 17561 9965 17564
rect 9999 17561 10011 17595
rect 9953 17555 10011 17561
rect 10226 17552 10232 17604
rect 10284 17592 10290 17604
rect 10428 17592 10456 17768
rect 10505 17731 10563 17737
rect 10505 17697 10517 17731
rect 10551 17728 10563 17731
rect 10778 17728 10784 17740
rect 10551 17700 10784 17728
rect 10551 17697 10563 17700
rect 10505 17691 10563 17697
rect 10778 17688 10784 17700
rect 10836 17728 10842 17740
rect 10836 17700 11008 17728
rect 10836 17688 10842 17700
rect 10980 17669 11008 17700
rect 11164 17669 11192 17768
rect 12529 17765 12541 17799
rect 12575 17796 12587 17799
rect 13170 17796 13176 17808
rect 12575 17768 13176 17796
rect 12575 17765 12587 17768
rect 12529 17759 12587 17765
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 15841 17799 15899 17805
rect 15841 17765 15853 17799
rect 15887 17796 15899 17799
rect 16666 17796 16672 17808
rect 15887 17768 16672 17796
rect 15887 17765 15899 17768
rect 15841 17759 15899 17765
rect 16666 17756 16672 17768
rect 16724 17756 16730 17808
rect 18417 17799 18475 17805
rect 18417 17765 18429 17799
rect 18463 17796 18475 17799
rect 18601 17799 18659 17805
rect 18601 17796 18613 17799
rect 18463 17768 18613 17796
rect 18463 17765 18475 17768
rect 18417 17759 18475 17765
rect 18601 17765 18613 17768
rect 18647 17765 18659 17799
rect 18601 17759 18659 17765
rect 20438 17756 20444 17808
rect 20496 17796 20502 17808
rect 20990 17796 20996 17808
rect 20496 17768 20996 17796
rect 20496 17756 20502 17768
rect 20990 17756 20996 17768
rect 21048 17796 21054 17808
rect 23569 17799 23627 17805
rect 23569 17796 23581 17799
rect 21048 17768 21220 17796
rect 21048 17756 21054 17768
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17728 11851 17731
rect 14829 17731 14887 17737
rect 14829 17728 14841 17731
rect 11839 17700 12296 17728
rect 11839 17697 11851 17700
rect 11793 17691 11851 17697
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 10704 17632 10885 17660
rect 10284 17564 10456 17592
rect 10597 17595 10655 17601
rect 10284 17552 10290 17564
rect 10597 17561 10609 17595
rect 10643 17561 10655 17595
rect 10597 17555 10655 17561
rect 10704 17592 10732 17632
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 10873 17623 10931 17629
rect 10965 17663 11023 17669
rect 10965 17629 10977 17663
rect 11011 17629 11023 17663
rect 10965 17623 11023 17629
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17629 11207 17663
rect 11149 17623 11207 17629
rect 11333 17663 11391 17669
rect 11333 17629 11345 17663
rect 11379 17629 11391 17663
rect 11333 17623 11391 17629
rect 11348 17592 11376 17623
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 12268 17669 12296 17700
rect 14476 17700 14841 17728
rect 14476 17672 14504 17700
rect 14829 17697 14841 17700
rect 14875 17697 14887 17731
rect 14829 17691 14887 17697
rect 15194 17688 15200 17740
rect 15252 17728 15258 17740
rect 21192 17737 21220 17768
rect 22848 17768 23581 17796
rect 15381 17731 15439 17737
rect 15381 17728 15393 17731
rect 15252 17700 15393 17728
rect 15252 17688 15258 17700
rect 15381 17697 15393 17700
rect 15427 17697 15439 17731
rect 18785 17731 18843 17737
rect 15381 17691 15439 17697
rect 18432 17700 18736 17728
rect 12161 17663 12219 17669
rect 12161 17660 12173 17663
rect 11664 17632 12173 17660
rect 11664 17620 11670 17632
rect 12161 17629 12173 17632
rect 12207 17629 12219 17663
rect 12161 17623 12219 17629
rect 12253 17663 12311 17669
rect 12253 17629 12265 17663
rect 12299 17660 12311 17663
rect 12299 17632 12480 17660
rect 12299 17629 12311 17632
rect 12253 17623 12311 17629
rect 11885 17595 11943 17601
rect 11885 17592 11897 17595
rect 10704 17564 11897 17592
rect 10612 17524 10640 17555
rect 10704 17536 10732 17564
rect 11885 17561 11897 17564
rect 11931 17561 11943 17595
rect 11885 17555 11943 17561
rect 12069 17595 12127 17601
rect 12069 17561 12081 17595
rect 12115 17561 12127 17595
rect 12069 17555 12127 17561
rect 9692 17496 10640 17524
rect 10686 17484 10692 17536
rect 10744 17484 10750 17536
rect 10781 17527 10839 17533
rect 10781 17493 10793 17527
rect 10827 17524 10839 17527
rect 11330 17524 11336 17536
rect 10827 17496 11336 17524
rect 10827 17493 10839 17496
rect 10781 17487 10839 17493
rect 11330 17484 11336 17496
rect 11388 17484 11394 17536
rect 11422 17484 11428 17536
rect 11480 17524 11486 17536
rect 12084 17524 12112 17555
rect 12452 17536 12480 17632
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 14642 17620 14648 17672
rect 14700 17620 14706 17672
rect 14734 17620 14740 17672
rect 14792 17620 14798 17672
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17629 15071 17663
rect 15013 17623 15071 17629
rect 15473 17663 15531 17669
rect 15473 17629 15485 17663
rect 15519 17660 15531 17663
rect 15562 17660 15568 17672
rect 15519 17632 15568 17660
rect 15519 17629 15531 17632
rect 15473 17623 15531 17629
rect 12526 17552 12532 17604
rect 12584 17552 12590 17604
rect 14550 17552 14556 17604
rect 14608 17592 14614 17604
rect 14752 17592 14780 17620
rect 15028 17592 15056 17623
rect 15562 17620 15568 17632
rect 15620 17620 15626 17672
rect 15654 17620 15660 17672
rect 15712 17620 15718 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 18432 17669 18460 17700
rect 18233 17663 18291 17669
rect 18233 17660 18245 17663
rect 18104 17632 18245 17660
rect 18104 17620 18110 17632
rect 18233 17629 18245 17632
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17660 18567 17663
rect 18555 17632 18644 17660
rect 18555 17629 18567 17632
rect 18509 17623 18567 17629
rect 15194 17592 15200 17604
rect 14608 17564 14964 17592
rect 15028 17564 15200 17592
rect 14608 17552 14614 17564
rect 11480 17496 12112 17524
rect 12161 17527 12219 17533
rect 11480 17484 11486 17496
rect 12161 17493 12173 17527
rect 12207 17524 12219 17527
rect 12250 17524 12256 17536
rect 12207 17496 12256 17524
rect 12207 17493 12219 17496
rect 12161 17487 12219 17493
rect 12250 17484 12256 17496
rect 12308 17524 12314 17536
rect 12345 17527 12403 17533
rect 12345 17524 12357 17527
rect 12308 17496 12357 17524
rect 12308 17484 12314 17496
rect 12345 17493 12357 17496
rect 12391 17493 12403 17527
rect 12345 17487 12403 17493
rect 12434 17484 12440 17536
rect 12492 17484 12498 17536
rect 14461 17527 14519 17533
rect 14461 17493 14473 17527
rect 14507 17524 14519 17527
rect 14826 17524 14832 17536
rect 14507 17496 14832 17524
rect 14507 17493 14519 17496
rect 14461 17487 14519 17493
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 14936 17533 14964 17564
rect 15194 17552 15200 17564
rect 15252 17592 15258 17604
rect 15672 17592 15700 17620
rect 18432 17592 18460 17623
rect 15252 17564 15700 17592
rect 18064 17564 18460 17592
rect 15252 17552 15258 17564
rect 18064 17536 18092 17564
rect 18616 17536 18644 17632
rect 18708 17592 18736 17700
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 18969 17731 19027 17737
rect 18969 17728 18981 17731
rect 18831 17700 18981 17728
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 18969 17697 18981 17700
rect 19015 17697 19027 17731
rect 21085 17731 21143 17737
rect 21085 17728 21097 17731
rect 18969 17691 19027 17697
rect 20364 17700 21097 17728
rect 18874 17620 18880 17672
rect 18932 17620 18938 17672
rect 20364 17669 20392 17700
rect 20916 17672 20944 17700
rect 21085 17697 21097 17700
rect 21131 17697 21143 17731
rect 21085 17691 21143 17697
rect 21177 17731 21235 17737
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 22002 17688 22008 17740
rect 22060 17728 22066 17740
rect 22848 17737 22876 17768
rect 23569 17765 23581 17768
rect 23615 17765 23627 17799
rect 23569 17759 23627 17765
rect 22833 17731 22891 17737
rect 22833 17728 22845 17731
rect 22060 17700 22845 17728
rect 22060 17688 22066 17700
rect 22833 17697 22845 17700
rect 22879 17697 22891 17731
rect 22833 17691 22891 17697
rect 23109 17731 23167 17737
rect 23109 17697 23121 17731
rect 23155 17728 23167 17731
rect 24673 17731 24731 17737
rect 24673 17728 24685 17731
rect 23155 17700 24685 17728
rect 23155 17697 23167 17700
rect 23109 17691 23167 17697
rect 24673 17697 24685 17700
rect 24719 17697 24731 17731
rect 24673 17691 24731 17697
rect 19061 17663 19119 17669
rect 19061 17629 19073 17663
rect 19107 17629 19119 17663
rect 20257 17663 20315 17669
rect 20257 17660 20269 17663
rect 19061 17623 19119 17629
rect 20180 17632 20269 17660
rect 19076 17592 19104 17623
rect 18708 17564 19104 17592
rect 20180 17536 20208 17632
rect 20257 17629 20269 17632
rect 20303 17629 20315 17663
rect 20257 17623 20315 17629
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 20438 17620 20444 17672
rect 20496 17620 20502 17672
rect 20622 17669 20628 17672
rect 20598 17663 20628 17669
rect 20598 17629 20610 17663
rect 20598 17623 20628 17629
rect 20622 17620 20628 17623
rect 20680 17620 20686 17672
rect 20714 17620 20720 17672
rect 20772 17620 20778 17672
rect 20898 17620 20904 17672
rect 20956 17620 20962 17672
rect 20993 17663 21051 17669
rect 20993 17629 21005 17663
rect 21039 17660 21051 17663
rect 21039 17632 21128 17660
rect 21039 17629 21051 17632
rect 20993 17623 21051 17629
rect 14921 17527 14979 17533
rect 14921 17493 14933 17527
rect 14967 17493 14979 17527
rect 14921 17487 14979 17493
rect 18046 17484 18052 17536
rect 18104 17484 18110 17536
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 20162 17484 20168 17536
rect 20220 17524 20226 17536
rect 21100 17524 21128 17632
rect 21266 17620 21272 17672
rect 21324 17620 21330 17672
rect 22741 17663 22799 17669
rect 22741 17629 22753 17663
rect 22787 17660 22799 17663
rect 23385 17663 23443 17669
rect 23385 17660 23397 17663
rect 22787 17632 23397 17660
rect 22787 17629 22799 17632
rect 22741 17623 22799 17629
rect 23124 17536 23152 17632
rect 23385 17629 23397 17632
rect 23431 17629 23443 17663
rect 23385 17623 23443 17629
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 23290 17552 23296 17604
rect 23348 17592 23354 17604
rect 23676 17592 23704 17623
rect 24118 17620 24124 17672
rect 24176 17660 24182 17672
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 24176 17632 24409 17660
rect 24176 17620 24182 17632
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 24397 17623 24455 17629
rect 23348 17564 23704 17592
rect 23348 17552 23354 17564
rect 25130 17552 25136 17604
rect 25188 17552 25194 17604
rect 21174 17524 21180 17536
rect 20220 17496 21180 17524
rect 20220 17484 20226 17496
rect 21174 17484 21180 17496
rect 21232 17484 21238 17536
rect 23106 17484 23112 17536
rect 23164 17484 23170 17536
rect 26145 17527 26203 17533
rect 26145 17493 26157 17527
rect 26191 17524 26203 17527
rect 33134 17524 33140 17536
rect 26191 17496 33140 17524
rect 26191 17493 26203 17496
rect 26145 17487 26203 17493
rect 33134 17484 33140 17496
rect 33192 17484 33198 17536
rect 1104 17434 35236 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 35236 17434
rect 1104 17360 35236 17382
rect 4890 17280 4896 17332
rect 4948 17320 4954 17332
rect 4985 17323 5043 17329
rect 4985 17320 4997 17323
rect 4948 17292 4997 17320
rect 4948 17280 4954 17292
rect 4985 17289 4997 17292
rect 5031 17289 5043 17323
rect 4985 17283 5043 17289
rect 5442 17280 5448 17332
rect 5500 17280 5506 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 5997 17323 6055 17329
rect 5997 17320 6009 17323
rect 5960 17292 6009 17320
rect 5960 17280 5966 17292
rect 5997 17289 6009 17292
rect 6043 17289 6055 17323
rect 5997 17283 6055 17289
rect 9030 17280 9036 17332
rect 9088 17320 9094 17332
rect 9088 17292 9352 17320
rect 9088 17280 9094 17292
rect 4706 17144 4712 17196
rect 4764 17184 4770 17196
rect 4893 17187 4951 17193
rect 4893 17184 4905 17187
rect 4764 17156 4905 17184
rect 4764 17144 4770 17156
rect 4893 17153 4905 17156
rect 4939 17184 4951 17187
rect 5460 17184 5488 17280
rect 8021 17255 8079 17261
rect 8021 17221 8033 17255
rect 8067 17252 8079 17255
rect 8938 17252 8944 17264
rect 8067 17224 8944 17252
rect 8067 17221 8079 17224
rect 8021 17215 8079 17221
rect 8938 17212 8944 17224
rect 8996 17252 9002 17264
rect 9125 17255 9183 17261
rect 9125 17252 9137 17255
rect 8996 17224 9137 17252
rect 8996 17212 9002 17224
rect 9125 17221 9137 17224
rect 9171 17221 9183 17255
rect 9324 17252 9352 17292
rect 9582 17280 9588 17332
rect 9640 17320 9646 17332
rect 9677 17323 9735 17329
rect 9677 17320 9689 17323
rect 9640 17292 9689 17320
rect 9640 17280 9646 17292
rect 9677 17289 9689 17292
rect 9723 17289 9735 17323
rect 9677 17283 9735 17289
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 11422 17320 11428 17332
rect 9907 17292 11428 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 11422 17280 11428 17292
rect 11480 17280 11486 17332
rect 13170 17280 13176 17332
rect 13228 17280 13234 17332
rect 13446 17280 13452 17332
rect 13504 17280 13510 17332
rect 14826 17280 14832 17332
rect 14884 17280 14890 17332
rect 15105 17323 15163 17329
rect 15105 17289 15117 17323
rect 15151 17320 15163 17323
rect 15194 17320 15200 17332
rect 15151 17292 15200 17320
rect 15151 17289 15163 17292
rect 15105 17283 15163 17289
rect 15194 17280 15200 17292
rect 15252 17280 15258 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 20824 17292 21465 17320
rect 9324 17224 9628 17252
rect 9125 17215 9183 17221
rect 4939 17156 5488 17184
rect 4939 17153 4951 17156
rect 4893 17147 4951 17153
rect 8754 17144 8760 17196
rect 8812 17144 8818 17196
rect 8846 17144 8852 17196
rect 8904 17144 8910 17196
rect 9030 17144 9036 17196
rect 9088 17144 9094 17196
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17184 9275 17187
rect 9398 17184 9404 17196
rect 9263 17156 9404 17184
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 9398 17144 9404 17156
rect 9456 17144 9462 17196
rect 9600 17193 9628 17224
rect 12250 17212 12256 17264
rect 12308 17212 12314 17264
rect 12526 17261 12532 17264
rect 12469 17255 12532 17261
rect 12469 17221 12481 17255
rect 12515 17221 12532 17255
rect 12469 17215 12532 17221
rect 12526 17212 12532 17215
rect 12584 17252 12590 17264
rect 12584 17224 13124 17252
rect 12584 17212 12590 17224
rect 13096 17196 13124 17224
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9585 17147 9643 17153
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 8662 17116 8668 17128
rect 8435 17088 8668 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 8662 17076 8668 17088
rect 8720 17076 8726 17128
rect 8864 17116 8892 17144
rect 9306 17116 9312 17128
rect 8864 17088 9312 17116
rect 9306 17076 9312 17088
rect 9364 17116 9370 17128
rect 9508 17116 9536 17147
rect 9858 17144 9864 17196
rect 9916 17144 9922 17196
rect 13078 17144 13084 17196
rect 13136 17144 13142 17196
rect 13188 17193 13216 17280
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17153 13231 17187
rect 13173 17147 13231 17153
rect 13357 17187 13415 17193
rect 13357 17153 13369 17187
rect 13403 17153 13415 17187
rect 13464 17184 13492 17280
rect 14844 17252 14872 17280
rect 18874 17252 18880 17264
rect 14844 17224 15240 17252
rect 13633 17187 13691 17193
rect 13633 17184 13645 17187
rect 13464 17156 13645 17184
rect 13357 17147 13415 17153
rect 13633 17153 13645 17156
rect 13679 17153 13691 17187
rect 13633 17147 13691 17153
rect 9364 17088 9536 17116
rect 9364 17076 9370 17088
rect 9674 17076 9680 17128
rect 9732 17116 9738 17128
rect 12250 17116 12256 17128
rect 9732 17088 12256 17116
rect 9732 17076 9738 17088
rect 12250 17076 12256 17088
rect 12308 17076 12314 17128
rect 12434 17076 12440 17128
rect 12492 17076 12498 17128
rect 13262 17116 13268 17128
rect 12636 17088 13268 17116
rect 9214 17008 9220 17060
rect 9272 17008 9278 17060
rect 9401 17051 9459 17057
rect 9401 17017 9413 17051
rect 9447 17048 9459 17051
rect 10686 17048 10692 17060
rect 9447 17020 10692 17048
rect 9447 17017 9459 17020
rect 9401 17011 9459 17017
rect 10686 17008 10692 17020
rect 10744 17008 10750 17060
rect 8478 16940 8484 16992
rect 8536 16940 8542 16992
rect 8570 16940 8576 16992
rect 8628 16989 8634 16992
rect 8628 16983 8668 16989
rect 8656 16949 8668 16983
rect 9232 16980 9260 17008
rect 10594 16980 10600 16992
rect 9232 16952 10600 16980
rect 8628 16943 8668 16949
rect 8628 16940 8634 16943
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 12452 16989 12480 17076
rect 12636 17057 12664 17088
rect 13262 17076 13268 17088
rect 13320 17116 13326 17128
rect 13372 17116 13400 17147
rect 14918 17144 14924 17196
rect 14976 17184 14982 17196
rect 15013 17187 15071 17193
rect 15013 17184 15025 17187
rect 14976 17156 15025 17184
rect 14976 17144 14982 17156
rect 15013 17153 15025 17156
rect 15059 17184 15071 17187
rect 15102 17184 15108 17196
rect 15059 17156 15108 17184
rect 15059 17153 15071 17156
rect 15013 17147 15071 17153
rect 15102 17144 15108 17156
rect 15160 17144 15166 17196
rect 15212 17193 15240 17224
rect 17972 17224 18880 17252
rect 17972 17196 18000 17224
rect 18874 17212 18880 17224
rect 18932 17212 18938 17264
rect 20824 17196 20852 17292
rect 21453 17289 21465 17292
rect 21499 17289 21511 17323
rect 21453 17283 21511 17289
rect 22002 17280 22008 17332
rect 22060 17280 22066 17332
rect 23109 17323 23167 17329
rect 23109 17289 23121 17323
rect 23155 17320 23167 17323
rect 23290 17320 23296 17332
rect 23155 17292 23296 17320
rect 23155 17289 23167 17292
rect 23109 17283 23167 17289
rect 23290 17280 23296 17292
rect 23348 17280 23354 17332
rect 24857 17323 24915 17329
rect 24857 17289 24869 17323
rect 24903 17320 24915 17323
rect 25130 17320 25136 17332
rect 24903 17292 25136 17320
rect 24903 17289 24915 17292
rect 24857 17283 24915 17289
rect 25130 17280 25136 17292
rect 25188 17280 25194 17332
rect 25317 17323 25375 17329
rect 25317 17289 25329 17323
rect 25363 17320 25375 17323
rect 25406 17320 25412 17332
rect 25363 17292 25412 17320
rect 25363 17289 25375 17292
rect 25317 17283 25375 17289
rect 20916 17224 21128 17252
rect 20916 17196 20944 17224
rect 15197 17187 15255 17193
rect 15197 17153 15209 17187
rect 15243 17153 15255 17187
rect 15197 17147 15255 17153
rect 17954 17144 17960 17196
rect 18012 17144 18018 17196
rect 18598 17144 18604 17196
rect 18656 17144 18662 17196
rect 20717 17187 20775 17193
rect 20717 17184 20729 17187
rect 20640 17156 20729 17184
rect 13320 17088 13400 17116
rect 13541 17119 13599 17125
rect 13320 17076 13326 17088
rect 13541 17085 13553 17119
rect 13587 17116 13599 17119
rect 18046 17116 18052 17128
rect 13587 17088 18052 17116
rect 13587 17085 13599 17088
rect 13541 17079 13599 17085
rect 18046 17076 18052 17088
rect 18104 17076 18110 17128
rect 18325 17119 18383 17125
rect 18325 17085 18337 17119
rect 18371 17116 18383 17119
rect 18509 17119 18567 17125
rect 18509 17116 18521 17119
rect 18371 17088 18521 17116
rect 18371 17085 18383 17088
rect 18325 17079 18383 17085
rect 18509 17085 18521 17088
rect 18555 17085 18567 17119
rect 18509 17079 18567 17085
rect 12621 17051 12679 17057
rect 12621 17017 12633 17051
rect 12667 17017 12679 17051
rect 14550 17048 14556 17060
rect 12621 17011 12679 17017
rect 13464 17020 14556 17048
rect 13464 16992 13492 17020
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 18616 17048 18644 17144
rect 20640 17128 20668 17156
rect 20717 17153 20729 17156
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 20806 17144 20812 17196
rect 20864 17144 20870 17196
rect 20898 17144 20904 17196
rect 20956 17144 20962 17196
rect 20990 17144 20996 17196
rect 21048 17144 21054 17196
rect 21100 17193 21128 17224
rect 21174 17212 21180 17264
rect 21232 17212 21238 17264
rect 21269 17255 21327 17261
rect 21269 17221 21281 17255
rect 21315 17252 21327 17255
rect 21315 17224 22048 17252
rect 21315 17221 21327 17224
rect 21269 17215 21327 17221
rect 21085 17187 21143 17193
rect 21085 17153 21097 17187
rect 21131 17153 21143 17187
rect 21192 17184 21220 17212
rect 22020 17193 22048 17224
rect 21361 17187 21419 17193
rect 21361 17184 21373 17187
rect 21192 17156 21373 17184
rect 21085 17147 21143 17153
rect 21361 17153 21373 17156
rect 21407 17153 21419 17187
rect 21361 17147 21419 17153
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17153 21879 17187
rect 21821 17147 21879 17153
rect 22005 17187 22063 17193
rect 22005 17153 22017 17187
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 24765 17187 24823 17193
rect 24765 17153 24777 17187
rect 24811 17184 24823 17187
rect 25332 17184 25360 17283
rect 25406 17280 25412 17292
rect 25464 17280 25470 17332
rect 24811 17156 25360 17184
rect 24811 17153 24823 17156
rect 24765 17147 24823 17153
rect 20622 17076 20628 17128
rect 20680 17076 20686 17128
rect 21836 17116 21864 17147
rect 21192 17088 21864 17116
rect 15672 17020 18644 17048
rect 15672 16992 15700 17020
rect 21192 16992 21220 17088
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16949 12495 16983
rect 12437 16943 12495 16949
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 13722 16940 13728 16992
rect 13780 16940 13786 16992
rect 15654 16940 15660 16992
rect 15712 16940 15718 16992
rect 18877 16983 18935 16989
rect 18877 16949 18889 16983
rect 18923 16980 18935 16983
rect 19334 16980 19340 16992
rect 18923 16952 19340 16980
rect 18923 16949 18935 16952
rect 18877 16943 18935 16949
rect 19334 16940 19340 16952
rect 19392 16940 19398 16992
rect 21174 16940 21180 16992
rect 21232 16940 21238 16992
rect 1104 16890 35248 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 35248 16890
rect 1104 16816 35248 16838
rect 8754 16736 8760 16788
rect 8812 16776 8818 16788
rect 10137 16779 10195 16785
rect 8812 16748 10088 16776
rect 8812 16736 8818 16748
rect 8021 16711 8079 16717
rect 8021 16677 8033 16711
rect 8067 16708 8079 16711
rect 8478 16708 8484 16720
rect 8067 16680 8484 16708
rect 8067 16677 8079 16680
rect 8021 16671 8079 16677
rect 8478 16668 8484 16680
rect 8536 16708 8542 16720
rect 10060 16708 10088 16748
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10226 16776 10232 16788
rect 10183 16748 10232 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10226 16736 10232 16748
rect 10284 16736 10290 16788
rect 10321 16779 10379 16785
rect 10321 16745 10333 16779
rect 10367 16776 10379 16779
rect 10778 16776 10784 16788
rect 10367 16748 10784 16776
rect 10367 16745 10379 16748
rect 10321 16739 10379 16745
rect 10778 16736 10784 16748
rect 10836 16736 10842 16788
rect 12621 16779 12679 16785
rect 12621 16745 12633 16779
rect 12667 16776 12679 16779
rect 12710 16776 12716 16788
rect 12667 16748 12716 16776
rect 12667 16745 12679 16748
rect 12621 16739 12679 16745
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 13446 16776 13452 16788
rect 12860 16748 13452 16776
rect 12860 16736 12866 16748
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 13722 16736 13728 16788
rect 13780 16736 13786 16788
rect 14277 16779 14335 16785
rect 14277 16745 14289 16779
rect 14323 16745 14335 16779
rect 14277 16739 14335 16745
rect 13740 16708 13768 16736
rect 14185 16711 14243 16717
rect 14185 16708 14197 16711
rect 8536 16680 9628 16708
rect 10060 16680 12388 16708
rect 13740 16680 14197 16708
rect 8536 16668 8542 16680
rect 3602 16600 3608 16652
rect 3660 16640 3666 16652
rect 3881 16643 3939 16649
rect 3881 16640 3893 16643
rect 3660 16612 3893 16640
rect 3660 16600 3666 16612
rect 3881 16609 3893 16612
rect 3927 16609 3939 16643
rect 3881 16603 3939 16609
rect 4157 16643 4215 16649
rect 4157 16609 4169 16643
rect 4203 16640 4215 16643
rect 4614 16640 4620 16652
rect 4203 16612 4620 16640
rect 4203 16609 4215 16612
rect 4157 16603 4215 16609
rect 4614 16600 4620 16612
rect 4672 16600 4678 16652
rect 8570 16600 8576 16652
rect 8628 16640 8634 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8628 16612 8953 16640
rect 8628 16600 8634 16612
rect 8941 16609 8953 16612
rect 8987 16640 8999 16643
rect 9490 16640 9496 16652
rect 8987 16612 9496 16640
rect 8987 16609 8999 16612
rect 8941 16603 8999 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9600 16640 9628 16680
rect 9600 16612 9904 16640
rect 6362 16532 6368 16584
rect 6420 16532 6426 16584
rect 6822 16532 6828 16584
rect 6880 16532 6886 16584
rect 9309 16575 9367 16581
rect 9309 16541 9321 16575
rect 9355 16541 9367 16575
rect 9309 16535 9367 16541
rect 9401 16575 9459 16581
rect 9401 16541 9413 16575
rect 9447 16572 9459 16575
rect 9600 16572 9628 16612
rect 9447 16544 9628 16572
rect 9876 16572 9904 16612
rect 9950 16600 9956 16652
rect 10008 16640 10014 16652
rect 10226 16640 10232 16652
rect 10008 16612 10232 16640
rect 10008 16600 10014 16612
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10428 16629 10456 16680
rect 10428 16601 10548 16629
rect 10520 16582 10548 16601
rect 10520 16581 10640 16582
rect 10520 16575 10661 16581
rect 9876 16544 10456 16572
rect 10520 16554 10615 16575
rect 9447 16541 9459 16544
rect 9401 16535 9459 16541
rect 4614 16464 4620 16516
rect 4672 16464 4678 16516
rect 5905 16507 5963 16513
rect 5905 16473 5917 16507
rect 5951 16504 5963 16507
rect 6840 16504 6868 16532
rect 5951 16476 6868 16504
rect 5951 16473 5963 16476
rect 5905 16467 5963 16473
rect 8938 16464 8944 16516
rect 8996 16504 9002 16516
rect 9033 16507 9091 16513
rect 9033 16504 9045 16507
rect 8996 16476 9045 16504
rect 8996 16464 9002 16476
rect 9033 16473 9045 16476
rect 9079 16473 9091 16507
rect 9324 16504 9352 16535
rect 9490 16504 9496 16516
rect 9324 16476 9496 16504
rect 9033 16467 9091 16473
rect 9490 16464 9496 16476
rect 9548 16464 9554 16516
rect 10318 16513 10324 16516
rect 10305 16507 10324 16513
rect 10305 16473 10317 16507
rect 10305 16467 10324 16473
rect 10318 16464 10324 16467
rect 10376 16464 10382 16516
rect 9398 16396 9404 16448
rect 9456 16436 9462 16448
rect 9585 16439 9643 16445
rect 9585 16436 9597 16439
rect 9456 16408 9597 16436
rect 9456 16396 9462 16408
rect 9585 16405 9597 16408
rect 9631 16405 9643 16439
rect 10428 16436 10456 16544
rect 10603 16541 10615 16554
rect 10649 16541 10661 16575
rect 10775 16575 10833 16581
rect 10775 16566 10787 16575
rect 10603 16535 10661 16541
rect 10704 16541 10787 16566
rect 10821 16541 10833 16575
rect 10704 16538 10833 16541
rect 10502 16464 10508 16516
rect 10560 16464 10566 16516
rect 10704 16504 10732 16538
rect 10775 16535 10833 16538
rect 12250 16532 12256 16584
rect 12308 16572 12314 16584
rect 12360 16581 12388 16680
rect 14185 16677 14197 16680
rect 14231 16677 14243 16711
rect 14292 16708 14320 16739
rect 14642 16736 14648 16788
rect 14700 16776 14706 16788
rect 14829 16779 14887 16785
rect 14829 16776 14841 16779
rect 14700 16748 14841 16776
rect 14700 16736 14706 16748
rect 14829 16745 14841 16748
rect 14875 16745 14887 16779
rect 14829 16739 14887 16745
rect 15654 16736 15660 16788
rect 15712 16736 15718 16788
rect 20806 16736 20812 16788
rect 20864 16736 20870 16788
rect 21174 16736 21180 16788
rect 21232 16736 21238 16788
rect 15470 16708 15476 16720
rect 14292 16680 15476 16708
rect 14185 16671 14243 16677
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 16485 16711 16543 16717
rect 16485 16708 16497 16711
rect 15856 16680 16497 16708
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 13909 16643 13967 16649
rect 13909 16640 13921 16643
rect 12584 16612 12940 16640
rect 12584 16600 12590 16612
rect 12912 16584 12940 16612
rect 13832 16612 13921 16640
rect 12345 16575 12403 16581
rect 12345 16572 12357 16575
rect 12308 16544 12357 16572
rect 12308 16532 12314 16544
rect 12345 16541 12357 16544
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 12618 16532 12624 16584
rect 12676 16532 12682 16584
rect 12894 16532 12900 16584
rect 12952 16532 12958 16584
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13633 16575 13691 16581
rect 13633 16572 13645 16575
rect 13412 16544 13645 16572
rect 13412 16532 13418 16544
rect 13633 16541 13645 16544
rect 13679 16572 13691 16575
rect 13722 16572 13728 16584
rect 13679 16544 13728 16572
rect 13679 16541 13691 16544
rect 13633 16535 13691 16541
rect 13722 16532 13728 16544
rect 13780 16532 13786 16584
rect 12526 16504 12532 16516
rect 10612 16476 12532 16504
rect 10612 16436 10640 16476
rect 12526 16464 12532 16476
rect 12584 16464 12590 16516
rect 13170 16464 13176 16516
rect 13228 16504 13234 16516
rect 13832 16504 13860 16612
rect 13909 16609 13921 16612
rect 13955 16609 13967 16643
rect 15856 16640 15884 16680
rect 16485 16677 16497 16680
rect 16531 16677 16543 16711
rect 17313 16711 17371 16717
rect 16485 16671 16543 16677
rect 16592 16680 16988 16708
rect 13909 16603 13967 16609
rect 14016 16612 15884 16640
rect 14016 16572 14044 16612
rect 13924 16544 14044 16572
rect 14093 16575 14151 16581
rect 13924 16513 13952 16544
rect 14093 16541 14105 16575
rect 14139 16541 14151 16575
rect 14093 16535 14151 16541
rect 13228 16476 13860 16504
rect 13228 16464 13234 16476
rect 10428 16408 10640 16436
rect 10689 16439 10747 16445
rect 9585 16399 9643 16405
rect 10689 16405 10701 16439
rect 10735 16436 10747 16439
rect 10778 16436 10784 16448
rect 10735 16408 10784 16436
rect 10735 16405 10747 16408
rect 10689 16399 10747 16405
rect 10778 16396 10784 16408
rect 10836 16396 10842 16448
rect 12805 16439 12863 16445
rect 12805 16405 12817 16439
rect 12851 16436 12863 16439
rect 13354 16436 13360 16448
rect 12851 16408 13360 16436
rect 12851 16405 12863 16408
rect 12805 16399 12863 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13832 16436 13860 16476
rect 13909 16507 13967 16513
rect 13909 16473 13921 16507
rect 13955 16473 13967 16507
rect 13909 16467 13967 16473
rect 14108 16436 14136 16535
rect 14182 16532 14188 16584
rect 14240 16572 14246 16584
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 14240 16544 14381 16572
rect 14240 16532 14246 16544
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 14550 16532 14556 16584
rect 14608 16532 14614 16584
rect 14826 16532 14832 16584
rect 14884 16572 14890 16584
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14884 16544 14933 16572
rect 14884 16532 14890 16544
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 14921 16535 14979 16541
rect 15102 16532 15108 16584
rect 15160 16532 15166 16584
rect 15856 16581 15884 16612
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16592 16640 16620 16680
rect 16448 16612 16620 16640
rect 16669 16643 16727 16649
rect 16448 16600 16454 16612
rect 16669 16609 16681 16643
rect 16715 16640 16727 16643
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16715 16612 16865 16640
rect 16715 16609 16727 16612
rect 16669 16603 16727 16609
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 16960 16640 16988 16680
rect 17313 16677 17325 16711
rect 17359 16708 17371 16711
rect 19242 16708 19248 16720
rect 17359 16680 19248 16708
rect 17359 16677 17371 16680
rect 17313 16671 17371 16677
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 18601 16643 18659 16649
rect 16960 16612 18552 16640
rect 16853 16603 16911 16609
rect 15841 16575 15899 16581
rect 15841 16541 15853 16575
rect 15887 16541 15899 16575
rect 15841 16535 15899 16541
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16541 16083 16575
rect 16025 16535 16083 16541
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16572 16175 16575
rect 16298 16572 16304 16584
rect 16163 16544 16304 16572
rect 16163 16541 16175 16544
rect 16117 16535 16175 16541
rect 15470 16464 15476 16516
rect 15528 16504 15534 16516
rect 16040 16504 16068 16535
rect 16298 16532 16304 16544
rect 16356 16572 16362 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16356 16544 16957 16572
rect 16356 16532 16362 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 18524 16572 18552 16612
rect 18601 16609 18613 16643
rect 18647 16640 18659 16643
rect 19334 16640 19340 16652
rect 18647 16612 19340 16640
rect 18647 16609 18659 16612
rect 18601 16603 18659 16609
rect 19334 16600 19340 16612
rect 19392 16640 19398 16652
rect 20824 16640 20852 16736
rect 21085 16643 21143 16649
rect 21085 16640 21097 16643
rect 19392 16612 19656 16640
rect 19392 16600 19398 16612
rect 18693 16575 18751 16581
rect 18693 16572 18705 16575
rect 18524 16544 18705 16572
rect 16945 16535 17003 16541
rect 18693 16541 18705 16544
rect 18739 16541 18751 16575
rect 18693 16535 18751 16541
rect 16209 16507 16267 16513
rect 16209 16504 16221 16507
rect 15528 16476 16221 16504
rect 15528 16464 15534 16476
rect 16209 16473 16221 16476
rect 16255 16473 16267 16507
rect 18708 16504 18736 16535
rect 18782 16532 18788 16584
rect 18840 16532 18846 16584
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19426 16572 19432 16584
rect 18923 16544 19432 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19426 16532 19432 16544
rect 19484 16572 19490 16584
rect 19628 16581 19656 16612
rect 20732 16612 20852 16640
rect 20916 16612 21097 16640
rect 19521 16575 19579 16581
rect 19521 16572 19533 16575
rect 19484 16544 19533 16572
rect 19484 16532 19490 16544
rect 19521 16541 19533 16544
rect 19567 16541 19579 16575
rect 19521 16535 19579 16541
rect 19613 16575 19671 16581
rect 19613 16541 19625 16575
rect 19659 16541 19671 16575
rect 19613 16535 19671 16541
rect 19797 16575 19855 16581
rect 19797 16541 19809 16575
rect 19843 16572 19855 16575
rect 20622 16572 20628 16584
rect 19843 16544 20628 16572
rect 19843 16541 19855 16544
rect 19797 16535 19855 16541
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 20732 16581 20760 16612
rect 20916 16584 20944 16612
rect 21085 16609 21097 16612
rect 21131 16609 21143 16643
rect 21085 16603 21143 16609
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16541 20775 16575
rect 20717 16535 20775 16541
rect 20809 16575 20867 16581
rect 20809 16541 20821 16575
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 18708 16476 19257 16504
rect 16209 16467 16267 16473
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 20162 16504 20168 16516
rect 19245 16467 19303 16473
rect 19352 16476 20168 16504
rect 13832 16408 14136 16436
rect 14642 16396 14648 16448
rect 14700 16396 14706 16448
rect 19061 16439 19119 16445
rect 19061 16405 19073 16439
rect 19107 16436 19119 16439
rect 19352 16436 19380 16476
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 20640 16504 20668 16532
rect 20824 16504 20852 16535
rect 20898 16532 20904 16584
rect 20956 16532 20962 16584
rect 20990 16532 20996 16584
rect 21048 16532 21054 16584
rect 33134 16532 33140 16584
rect 33192 16532 33198 16584
rect 21266 16504 21272 16516
rect 20640 16476 21272 16504
rect 21266 16464 21272 16476
rect 21324 16464 21330 16516
rect 34333 16507 34391 16513
rect 34333 16473 34345 16507
rect 34379 16504 34391 16507
rect 34882 16504 34888 16516
rect 34379 16476 34888 16504
rect 34379 16473 34391 16476
rect 34333 16467 34391 16473
rect 34882 16464 34888 16476
rect 34940 16464 34946 16516
rect 19107 16408 19380 16436
rect 19429 16439 19487 16445
rect 19107 16405 19119 16408
rect 19061 16399 19119 16405
rect 19429 16405 19441 16439
rect 19475 16436 19487 16439
rect 19978 16436 19984 16448
rect 19475 16408 19984 16436
rect 19475 16405 19487 16408
rect 19429 16399 19487 16405
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 1104 16346 35236 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 35236 16346
rect 1104 16272 35236 16294
rect 4525 16235 4583 16241
rect 4525 16201 4537 16235
rect 4571 16232 4583 16235
rect 4614 16232 4620 16244
rect 4571 16204 4620 16232
rect 4571 16201 4583 16204
rect 4525 16195 4583 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 4706 16192 4712 16244
rect 4764 16192 4770 16244
rect 6362 16232 6368 16244
rect 4816 16204 6368 16232
rect 4341 16167 4399 16173
rect 4341 16133 4353 16167
rect 4387 16164 4399 16167
rect 4724 16164 4752 16192
rect 4816 16173 4844 16204
rect 6362 16192 6368 16204
rect 6420 16232 6426 16244
rect 9217 16235 9275 16241
rect 6420 16204 7144 16232
rect 6420 16192 6426 16204
rect 4387 16136 4752 16164
rect 4801 16167 4859 16173
rect 4387 16133 4399 16136
rect 4341 16127 4399 16133
rect 4448 16105 4476 16136
rect 4801 16133 4813 16167
rect 4847 16133 4859 16167
rect 4801 16127 4859 16133
rect 4433 16099 4491 16105
rect 4433 16065 4445 16099
rect 4479 16096 4491 16099
rect 4479 16068 4513 16096
rect 4479 16065 4491 16068
rect 4433 16059 4491 16065
rect 5258 16056 5264 16108
rect 5316 16056 5322 16108
rect 5445 16099 5503 16105
rect 5445 16065 5457 16099
rect 5491 16096 5503 16099
rect 5813 16099 5871 16105
rect 5491 16068 5580 16096
rect 5491 16065 5503 16068
rect 5445 16059 5503 16065
rect 5552 15892 5580 16068
rect 5813 16065 5825 16099
rect 5859 16065 5871 16099
rect 5813 16059 5871 16065
rect 5997 16099 6055 16105
rect 5997 16065 6009 16099
rect 6043 16065 6055 16099
rect 5997 16059 6055 16065
rect 6181 16099 6239 16105
rect 6181 16065 6193 16099
rect 6227 16096 6239 16099
rect 6454 16096 6460 16108
rect 6227 16068 6460 16096
rect 6227 16065 6239 16068
rect 6181 16059 6239 16065
rect 5828 15960 5856 16059
rect 6012 16028 6040 16059
rect 6454 16056 6460 16068
rect 6512 16056 6518 16108
rect 6822 16056 6828 16108
rect 6880 16056 6886 16108
rect 7116 16105 7144 16204
rect 9217 16201 9229 16235
rect 9263 16232 9275 16235
rect 14461 16235 14519 16241
rect 9263 16204 13584 16232
rect 9263 16201 9275 16204
rect 9217 16195 9275 16201
rect 8478 16164 8484 16176
rect 7958 16136 8484 16164
rect 8478 16124 8484 16136
rect 8536 16124 8542 16176
rect 8570 16124 8576 16176
rect 8628 16124 8634 16176
rect 9030 16124 9036 16176
rect 9088 16164 9094 16176
rect 9309 16167 9367 16173
rect 9309 16164 9321 16167
rect 9088 16136 9321 16164
rect 9088 16124 9094 16136
rect 9309 16133 9321 16136
rect 9355 16133 9367 16167
rect 9309 16127 9367 16133
rect 9490 16124 9496 16176
rect 9548 16124 9554 16176
rect 11532 16136 12480 16164
rect 7101 16099 7159 16105
rect 7101 16065 7113 16099
rect 7147 16065 7159 16099
rect 8665 16099 8723 16105
rect 8665 16096 8677 16099
rect 7101 16059 7159 16065
rect 7944 16068 8677 16096
rect 7944 16040 7972 16068
rect 8665 16065 8677 16068
rect 8711 16065 8723 16099
rect 8665 16059 8723 16065
rect 8941 16099 8999 16105
rect 8941 16065 8953 16099
rect 8987 16096 8999 16099
rect 9508 16096 9536 16124
rect 8987 16068 9536 16096
rect 8987 16065 8999 16068
rect 8941 16059 8999 16065
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 11532 16105 11560 16136
rect 11808 16105 11836 16136
rect 11517 16099 11575 16105
rect 11517 16096 11529 16099
rect 11296 16068 11529 16096
rect 11296 16056 11302 16068
rect 11517 16065 11529 16068
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 11701 16099 11759 16105
rect 11701 16065 11713 16099
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11793 16099 11851 16105
rect 11793 16065 11805 16099
rect 11839 16065 11851 16099
rect 11793 16059 11851 16065
rect 11977 16099 12035 16105
rect 11977 16065 11989 16099
rect 12023 16096 12035 16099
rect 12158 16096 12164 16108
rect 12023 16068 12164 16096
rect 12023 16065 12035 16068
rect 11977 16059 12035 16065
rect 6012 16000 6684 16028
rect 6656 15972 6684 16000
rect 7926 15988 7932 16040
rect 7984 15988 7990 16040
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 9033 16031 9091 16037
rect 9033 16028 9045 16031
rect 8444 16000 9045 16028
rect 8444 15988 8450 16000
rect 9033 15997 9045 16000
rect 9079 15997 9091 16031
rect 9033 15991 9091 15997
rect 9677 16031 9735 16037
rect 9677 15997 9689 16031
rect 9723 16028 9735 16031
rect 10042 16028 10048 16040
rect 9723 16000 10048 16028
rect 9723 15997 9735 16000
rect 9677 15991 9735 15997
rect 6546 15960 6552 15972
rect 5828 15932 6552 15960
rect 6546 15920 6552 15932
rect 6604 15920 6610 15972
rect 6638 15920 6644 15972
rect 6696 15920 6702 15972
rect 9048 15960 9076 15991
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 11716 16028 11744 16059
rect 11992 16028 12020 16059
rect 12158 16056 12164 16068
rect 12216 16056 12222 16108
rect 12452 16096 12480 16136
rect 12728 16136 13124 16164
rect 12728 16108 12756 16136
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 12452 16094 12512 16096
rect 12544 16094 12633 16096
rect 12452 16068 12633 16094
rect 12484 16066 12572 16068
rect 12621 16065 12633 16068
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 12710 16056 12716 16108
rect 12768 16056 12774 16108
rect 12805 16099 12863 16105
rect 12805 16065 12817 16099
rect 12851 16096 12863 16099
rect 12986 16096 12992 16108
rect 12851 16068 12992 16096
rect 12851 16065 12863 16068
rect 12805 16059 12863 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 13096 16105 13124 16136
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16065 13139 16099
rect 13081 16059 13139 16065
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 13556 16105 13584 16204
rect 14461 16201 14473 16235
rect 14507 16232 14519 16235
rect 14826 16232 14832 16244
rect 14507 16204 14832 16232
rect 14507 16201 14519 16204
rect 14461 16195 14519 16201
rect 14826 16192 14832 16204
rect 14884 16192 14890 16244
rect 15378 16192 15384 16244
rect 15436 16192 15442 16244
rect 16393 16235 16451 16241
rect 16393 16201 16405 16235
rect 16439 16232 16451 16235
rect 16574 16232 16580 16244
rect 16439 16204 16580 16232
rect 16439 16201 16451 16204
rect 16393 16195 16451 16201
rect 16574 16192 16580 16204
rect 16632 16192 16638 16244
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 19978 16232 19984 16244
rect 18840 16204 19984 16232
rect 18840 16192 18846 16204
rect 19978 16192 19984 16204
rect 20036 16192 20042 16244
rect 20254 16192 20260 16244
rect 20312 16232 20318 16244
rect 20312 16204 21036 16232
rect 20312 16192 20318 16204
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 15289 16099 15347 16105
rect 15289 16096 15301 16099
rect 13771 16068 15301 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 15289 16065 15301 16068
rect 15335 16065 15347 16099
rect 15396 16096 15424 16192
rect 15657 16167 15715 16173
rect 15657 16133 15669 16167
rect 15703 16164 15715 16167
rect 16209 16167 16267 16173
rect 16209 16164 16221 16167
rect 15703 16136 16221 16164
rect 15703 16133 15715 16136
rect 15657 16127 15715 16133
rect 16209 16133 16221 16136
rect 16255 16164 16267 16167
rect 16255 16136 16712 16164
rect 16255 16133 16267 16136
rect 16209 16127 16267 16133
rect 16684 16105 16712 16136
rect 19242 16124 19248 16176
rect 19300 16164 19306 16176
rect 21008 16173 21036 16204
rect 21082 16192 21088 16244
rect 21140 16232 21146 16244
rect 21177 16235 21235 16241
rect 21177 16232 21189 16235
rect 21140 16204 21189 16232
rect 21140 16192 21146 16204
rect 21177 16201 21189 16204
rect 21223 16201 21235 16235
rect 21177 16195 21235 16201
rect 20809 16167 20867 16173
rect 20809 16164 20821 16167
rect 19300 16136 20821 16164
rect 19300 16124 19306 16136
rect 19904 16105 19932 16136
rect 15473 16099 15531 16105
rect 15473 16096 15485 16099
rect 15396 16068 15485 16096
rect 15289 16059 15347 16065
rect 15473 16065 15485 16068
rect 15519 16096 15531 16099
rect 15565 16099 15623 16105
rect 15565 16096 15577 16099
rect 15519 16068 15577 16096
rect 15519 16065 15531 16068
rect 15473 16059 15531 16065
rect 15565 16065 15577 16068
rect 15611 16065 15623 16099
rect 15565 16059 15623 16065
rect 15749 16099 15807 16105
rect 15749 16065 15761 16099
rect 15795 16065 15807 16099
rect 15749 16059 15807 16065
rect 16485 16099 16543 16105
rect 16485 16065 16497 16099
rect 16531 16065 16543 16099
rect 16485 16059 16543 16065
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16065 16727 16099
rect 16669 16059 16727 16065
rect 19889 16099 19947 16105
rect 19889 16065 19901 16099
rect 19935 16065 19947 16099
rect 19889 16059 19947 16065
rect 10468 16000 12020 16028
rect 10468 15988 10474 16000
rect 12250 15988 12256 16040
rect 12308 16028 12314 16040
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12308 16000 12909 16028
rect 12308 15988 12314 16000
rect 12897 15997 12909 16000
rect 12943 15997 12955 16031
rect 15304 16028 15332 16059
rect 15764 16028 15792 16059
rect 15304 16000 15792 16028
rect 12897 15991 12955 15997
rect 16500 15972 16528 16059
rect 20070 16056 20076 16108
rect 20128 16056 20134 16108
rect 20180 16105 20208 16136
rect 20809 16133 20821 16136
rect 20855 16133 20867 16167
rect 20809 16127 20867 16133
rect 20993 16167 21051 16173
rect 20993 16133 21005 16167
rect 21039 16133 21051 16167
rect 20993 16127 21051 16133
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 20254 16056 20260 16108
rect 20312 16096 20318 16108
rect 20349 16099 20407 16105
rect 20349 16096 20361 16099
rect 20312 16068 20361 16096
rect 20312 16056 20318 16068
rect 20349 16065 20361 16068
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 20438 16056 20444 16108
rect 20496 16056 20502 16108
rect 20530 16056 20536 16108
rect 20588 16056 20594 16108
rect 21192 16096 21220 16195
rect 23106 16192 23112 16244
rect 23164 16192 23170 16244
rect 23290 16192 23296 16244
rect 23348 16192 23354 16244
rect 23753 16235 23811 16241
rect 23753 16201 23765 16235
rect 23799 16232 23811 16235
rect 25593 16235 25651 16241
rect 23799 16204 24164 16232
rect 23799 16201 23811 16204
rect 23753 16195 23811 16201
rect 23308 16164 23336 16192
rect 24136 16173 24164 16204
rect 25593 16201 25605 16235
rect 25639 16232 25651 16235
rect 33134 16232 33140 16244
rect 25639 16204 33140 16232
rect 25639 16201 25651 16204
rect 25593 16195 25651 16201
rect 33134 16192 33140 16204
rect 33192 16192 33198 16244
rect 22480 16136 23336 16164
rect 24121 16167 24179 16173
rect 22480 16108 22508 16136
rect 24121 16133 24133 16167
rect 24167 16133 24179 16167
rect 25777 16167 25835 16173
rect 25777 16164 25789 16167
rect 25346 16136 25789 16164
rect 24121 16127 24179 16133
rect 25777 16133 25789 16136
rect 25823 16133 25835 16167
rect 25777 16127 25835 16133
rect 21453 16099 21511 16105
rect 21453 16096 21465 16099
rect 21192 16068 21465 16096
rect 21453 16065 21465 16068
rect 21499 16065 21511 16099
rect 21453 16059 21511 16065
rect 22002 16056 22008 16108
rect 22060 16056 22066 16108
rect 22462 16056 22468 16108
rect 22520 16056 22526 16108
rect 22649 16099 22707 16105
rect 22649 16065 22661 16099
rect 22695 16065 22707 16099
rect 22649 16059 22707 16065
rect 19981 16031 20039 16037
rect 19981 15997 19993 16031
rect 20027 16028 20039 16031
rect 21269 16031 21327 16037
rect 21269 16028 21281 16031
rect 20027 16000 21281 16028
rect 20027 15997 20039 16000
rect 19981 15991 20039 15997
rect 21269 15997 21281 16000
rect 21315 15997 21327 16031
rect 21269 15991 21327 15997
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 16028 21695 16031
rect 21913 16031 21971 16037
rect 21913 16028 21925 16031
rect 21683 16000 21925 16028
rect 21683 15997 21695 16000
rect 21637 15991 21695 15997
rect 21913 15997 21925 16000
rect 21959 15997 21971 16031
rect 21913 15991 21971 15997
rect 22664 16028 22692 16059
rect 22830 16056 22836 16108
rect 22888 16096 22894 16108
rect 22925 16099 22983 16105
rect 22925 16096 22937 16099
rect 22888 16068 22937 16096
rect 22888 16056 22894 16068
rect 22925 16065 22937 16068
rect 22971 16096 22983 16099
rect 23385 16099 23443 16105
rect 23385 16096 23397 16099
rect 22971 16068 23397 16096
rect 22971 16065 22983 16068
rect 22925 16059 22983 16065
rect 23385 16065 23397 16068
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 25406 16056 25412 16108
rect 25464 16096 25470 16108
rect 25869 16099 25927 16105
rect 25869 16096 25881 16099
rect 25464 16068 25881 16096
rect 25464 16056 25470 16068
rect 25869 16065 25881 16068
rect 25915 16096 25927 16099
rect 26050 16096 26056 16108
rect 25915 16068 26056 16096
rect 25915 16065 25927 16068
rect 25869 16059 25927 16065
rect 26050 16056 26056 16068
rect 26108 16096 26114 16108
rect 26145 16099 26203 16105
rect 26145 16096 26157 16099
rect 26108 16068 26157 16096
rect 26108 16056 26114 16068
rect 26145 16065 26157 16068
rect 26191 16065 26203 16099
rect 26145 16059 26203 16065
rect 23293 16031 23351 16037
rect 23293 16028 23305 16031
rect 22664 16000 23305 16028
rect 9769 15963 9827 15969
rect 9769 15960 9781 15963
rect 9048 15932 9781 15960
rect 9769 15929 9781 15932
rect 9815 15929 9827 15963
rect 9769 15923 9827 15929
rect 10226 15920 10232 15972
rect 10284 15960 10290 15972
rect 10597 15963 10655 15969
rect 10597 15960 10609 15963
rect 10284 15932 10609 15960
rect 10284 15920 10290 15932
rect 10597 15929 10609 15932
rect 10643 15929 10655 15963
rect 10597 15923 10655 15929
rect 12161 15963 12219 15969
rect 12161 15929 12173 15963
rect 12207 15960 12219 15963
rect 12986 15960 12992 15972
rect 12207 15932 12992 15960
rect 12207 15929 12219 15932
rect 12161 15923 12219 15929
rect 12986 15920 12992 15932
rect 13044 15960 13050 15972
rect 15381 15963 15439 15969
rect 13044 15932 13400 15960
rect 13044 15920 13050 15932
rect 6730 15892 6736 15904
rect 5552 15864 6736 15892
rect 6730 15852 6736 15864
rect 6788 15852 6794 15904
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 9950 15892 9956 15904
rect 9907 15864 9956 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 9950 15852 9956 15864
rect 10008 15852 10014 15904
rect 11517 15895 11575 15901
rect 11517 15861 11529 15895
rect 11563 15892 11575 15895
rect 11606 15892 11612 15904
rect 11563 15864 11612 15892
rect 11563 15861 11575 15864
rect 11517 15855 11575 15861
rect 11606 15852 11612 15864
rect 11664 15852 11670 15904
rect 12066 15852 12072 15904
rect 12124 15852 12130 15904
rect 12342 15852 12348 15904
rect 12400 15892 12406 15904
rect 12529 15895 12587 15901
rect 12529 15892 12541 15895
rect 12400 15864 12541 15892
rect 12400 15852 12406 15864
rect 12529 15861 12541 15864
rect 12575 15861 12587 15895
rect 12529 15855 12587 15861
rect 13262 15852 13268 15904
rect 13320 15852 13326 15904
rect 13372 15892 13400 15932
rect 15381 15929 15393 15963
rect 15427 15960 15439 15963
rect 16482 15960 16488 15972
rect 15427 15932 16488 15960
rect 15427 15929 15439 15932
rect 15381 15923 15439 15929
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 20717 15963 20775 15969
rect 20717 15929 20729 15963
rect 20763 15960 20775 15963
rect 20898 15960 20904 15972
rect 20763 15932 20904 15960
rect 20763 15929 20775 15932
rect 20717 15923 20775 15929
rect 20898 15920 20904 15932
rect 20956 15920 20962 15972
rect 22373 15963 22431 15969
rect 22373 15929 22385 15963
rect 22419 15960 22431 15963
rect 22664 15960 22692 16000
rect 23293 15997 23305 16000
rect 23339 15997 23351 16031
rect 23293 15991 23351 15997
rect 23845 16031 23903 16037
rect 23845 15997 23857 16031
rect 23891 16028 23903 16031
rect 24118 16028 24124 16040
rect 23891 16000 24124 16028
rect 23891 15997 23903 16000
rect 23845 15991 23903 15997
rect 24118 15988 24124 16000
rect 24176 15988 24182 16040
rect 22419 15932 22692 15960
rect 22419 15929 22431 15932
rect 22373 15923 22431 15929
rect 15654 15892 15660 15904
rect 13372 15864 15660 15892
rect 15654 15852 15660 15864
rect 15712 15852 15718 15904
rect 16209 15895 16267 15901
rect 16209 15861 16221 15895
rect 16255 15892 16267 15895
rect 16298 15892 16304 15904
rect 16255 15864 16304 15892
rect 16255 15861 16267 15864
rect 16209 15855 16267 15861
rect 16298 15852 16304 15864
rect 16356 15852 16362 15904
rect 16758 15852 16764 15904
rect 16816 15852 16822 15904
rect 1104 15802 35248 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 35248 15802
rect 1104 15728 35248 15750
rect 6178 15648 6184 15700
rect 6236 15648 6242 15700
rect 6822 15688 6828 15700
rect 6380 15660 6828 15688
rect 1394 15444 1400 15496
rect 1452 15444 1458 15496
rect 1581 15351 1639 15357
rect 1581 15317 1593 15351
rect 1627 15348 1639 15351
rect 4338 15348 4344 15360
rect 1627 15320 4344 15348
rect 1627 15317 1639 15320
rect 1581 15311 1639 15317
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 6196 15348 6224 15648
rect 6380 15493 6408 15660
rect 6822 15648 6828 15660
rect 6880 15648 6886 15700
rect 7009 15691 7067 15697
rect 7009 15657 7021 15691
rect 7055 15688 7067 15691
rect 7190 15688 7196 15700
rect 7055 15660 7196 15688
rect 7055 15657 7067 15660
rect 7009 15651 7067 15657
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8846 15688 8852 15700
rect 8527 15660 8852 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 8846 15648 8852 15660
rect 8904 15648 8910 15700
rect 10137 15691 10195 15697
rect 10137 15657 10149 15691
rect 10183 15688 10195 15691
rect 10318 15688 10324 15700
rect 10183 15660 10324 15688
rect 10183 15657 10195 15660
rect 10137 15651 10195 15657
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 11606 15648 11612 15700
rect 11664 15688 11670 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11664 15660 12357 15688
rect 11664 15648 11670 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 12345 15651 12403 15657
rect 12805 15691 12863 15697
rect 12805 15657 12817 15691
rect 12851 15688 12863 15691
rect 13170 15688 13176 15700
rect 12851 15660 13176 15688
rect 12851 15657 12863 15660
rect 12805 15651 12863 15657
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 15286 15648 15292 15700
rect 15344 15648 15350 15700
rect 15565 15691 15623 15697
rect 15565 15657 15577 15691
rect 15611 15688 15623 15691
rect 16209 15691 16267 15697
rect 15611 15660 16160 15688
rect 15611 15657 15623 15660
rect 15565 15651 15623 15657
rect 6454 15580 6460 15632
rect 6512 15580 6518 15632
rect 6638 15580 6644 15632
rect 6696 15620 6702 15632
rect 6914 15620 6920 15632
rect 6696 15592 6920 15620
rect 6696 15580 6702 15592
rect 6914 15580 6920 15592
rect 6972 15620 6978 15632
rect 10597 15623 10655 15629
rect 6972 15592 7328 15620
rect 6972 15580 6978 15592
rect 6472 15552 6500 15580
rect 6733 15555 6791 15561
rect 6733 15552 6745 15555
rect 6472 15524 6745 15552
rect 6733 15521 6745 15524
rect 6779 15552 6791 15555
rect 6779 15524 7236 15552
rect 6779 15521 6791 15524
rect 6733 15515 6791 15521
rect 6546 15493 6552 15496
rect 6365 15487 6423 15493
rect 6365 15453 6377 15487
rect 6411 15453 6423 15487
rect 6365 15447 6423 15453
rect 6512 15487 6552 15493
rect 6512 15453 6524 15487
rect 6512 15447 6552 15453
rect 6546 15444 6552 15447
rect 6604 15444 6610 15496
rect 7208 15428 7236 15524
rect 7300 15496 7328 15592
rect 10597 15589 10609 15623
rect 10643 15620 10655 15623
rect 10686 15620 10692 15632
rect 10643 15592 10692 15620
rect 10643 15589 10655 15592
rect 10597 15583 10655 15589
rect 10686 15580 10692 15592
rect 10744 15580 10750 15632
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 12710 15620 12716 15632
rect 12124 15592 12716 15620
rect 12124 15580 12130 15592
rect 12710 15580 12716 15592
rect 12768 15580 12774 15632
rect 12897 15623 12955 15629
rect 12897 15589 12909 15623
rect 12943 15620 12955 15623
rect 12986 15620 12992 15632
rect 12943 15592 12992 15620
rect 12943 15589 12955 15592
rect 12897 15583 12955 15589
rect 12986 15580 12992 15592
rect 13044 15580 13050 15632
rect 13354 15580 13360 15632
rect 13412 15580 13418 15632
rect 16132 15620 16160 15660
rect 16209 15657 16221 15691
rect 16255 15688 16267 15691
rect 16574 15688 16580 15700
rect 16255 15660 16580 15688
rect 16255 15657 16267 15660
rect 16209 15651 16267 15657
rect 16574 15648 16580 15660
rect 16632 15648 16638 15700
rect 16758 15648 16764 15700
rect 16816 15648 16822 15700
rect 20901 15691 20959 15697
rect 20901 15657 20913 15691
rect 20947 15688 20959 15691
rect 22002 15688 22008 15700
rect 20947 15660 22008 15688
rect 20947 15657 20959 15660
rect 20901 15651 20959 15657
rect 22002 15648 22008 15660
rect 22060 15648 22066 15700
rect 22373 15691 22431 15697
rect 22373 15657 22385 15691
rect 22419 15688 22431 15691
rect 22462 15688 22468 15700
rect 22419 15660 22468 15688
rect 22419 15657 22431 15660
rect 22373 15651 22431 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 23753 15691 23811 15697
rect 23753 15657 23765 15691
rect 23799 15688 23811 15691
rect 24118 15688 24124 15700
rect 23799 15660 24124 15688
rect 23799 15657 23811 15660
rect 23753 15651 23811 15657
rect 24118 15648 24124 15660
rect 24176 15648 24182 15700
rect 16390 15620 16396 15632
rect 16132 15592 16396 15620
rect 16390 15580 16396 15592
rect 16448 15580 16454 15632
rect 16482 15580 16488 15632
rect 16540 15580 16546 15632
rect 7745 15555 7803 15561
rect 7745 15521 7757 15555
rect 7791 15552 7803 15555
rect 10226 15552 10232 15564
rect 7791 15524 8248 15552
rect 7791 15521 7803 15524
rect 7745 15515 7803 15521
rect 8220 15496 8248 15524
rect 9324 15524 10232 15552
rect 7282 15444 7288 15496
rect 7340 15444 7346 15496
rect 7926 15484 7932 15496
rect 7760 15456 7932 15484
rect 7190 15376 7196 15428
rect 7248 15416 7254 15428
rect 7760 15416 7788 15456
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 8202 15444 8208 15496
rect 8260 15444 8266 15496
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8386 15484 8392 15496
rect 8343 15456 8392 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 9324 15425 9352 15524
rect 9692 15496 9720 15524
rect 10226 15512 10232 15524
rect 10284 15552 10290 15564
rect 12529 15555 12587 15561
rect 10284 15524 11928 15552
rect 10284 15512 10290 15524
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 7248 15388 7788 15416
rect 7837 15419 7895 15425
rect 7248 15376 7254 15388
rect 7837 15385 7849 15419
rect 7883 15416 7895 15419
rect 9309 15419 9367 15425
rect 9309 15416 9321 15419
rect 7883 15388 9321 15416
rect 7883 15385 7895 15388
rect 7837 15379 7895 15385
rect 9309 15385 9321 15388
rect 9355 15385 9367 15419
rect 9508 15416 9536 15447
rect 9674 15444 9680 15496
rect 9732 15444 9738 15496
rect 9766 15444 9772 15496
rect 9824 15444 9830 15496
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 10042 15484 10048 15496
rect 9907 15456 10048 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 10410 15444 10416 15496
rect 10468 15444 10474 15496
rect 10778 15444 10784 15496
rect 10836 15444 10842 15496
rect 11057 15487 11115 15493
rect 11057 15453 11069 15487
rect 11103 15453 11115 15487
rect 11057 15447 11115 15453
rect 11072 15416 11100 15447
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11900 15493 11928 15524
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 13262 15552 13268 15564
rect 12575 15524 13268 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13262 15512 13268 15524
rect 13320 15512 13326 15564
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11296 15456 11437 15484
rect 11296 15444 11302 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11885 15487 11943 15493
rect 11885 15453 11897 15487
rect 11931 15453 11943 15487
rect 11885 15447 11943 15453
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15484 12311 15487
rect 12342 15484 12348 15496
rect 12299 15456 12348 15484
rect 12299 15453 12311 15456
rect 12253 15447 12311 15453
rect 9508 15388 11100 15416
rect 9309 15379 9367 15385
rect 7852 15348 7880 15379
rect 10796 15360 10824 15388
rect 6196 15320 7880 15348
rect 10778 15308 10784 15360
rect 10836 15308 10842 15360
rect 11900 15348 11928 15447
rect 12342 15444 12348 15456
rect 12400 15444 12406 15496
rect 12894 15444 12900 15496
rect 12952 15444 12958 15496
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13372 15493 13400 15580
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 15102 15552 15108 15564
rect 13872 15524 15108 15552
rect 13872 15512 13878 15524
rect 15102 15512 15108 15524
rect 15160 15552 15166 15564
rect 15197 15555 15255 15561
rect 15197 15552 15209 15555
rect 15160 15524 15209 15552
rect 15160 15512 15166 15524
rect 15197 15521 15209 15524
rect 15243 15521 15255 15555
rect 15197 15515 15255 15521
rect 13081 15487 13139 15493
rect 13081 15484 13093 15487
rect 13044 15456 13093 15484
rect 13044 15444 13050 15456
rect 13081 15453 13093 15456
rect 13127 15453 13139 15487
rect 13081 15447 13139 15453
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15453 13231 15487
rect 13173 15447 13231 15453
rect 13357 15487 13415 15493
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13357 15447 13415 15453
rect 12360 15416 12388 15444
rect 13188 15416 13216 15447
rect 13538 15444 13544 15496
rect 13596 15484 13602 15496
rect 13596 15456 15240 15484
rect 13596 15444 13602 15456
rect 12360 15388 13216 15416
rect 13722 15376 13728 15428
rect 13780 15416 13786 15428
rect 15105 15419 15163 15425
rect 15105 15416 15117 15419
rect 13780 15388 15117 15416
rect 13780 15376 13786 15388
rect 15105 15385 15117 15388
rect 15151 15385 15163 15419
rect 15212 15416 15240 15456
rect 15378 15444 15384 15496
rect 15436 15444 15442 15496
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 16117 15487 16175 15493
rect 16117 15484 16129 15487
rect 15712 15456 16129 15484
rect 15712 15444 15718 15456
rect 16117 15453 16129 15456
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15453 16359 15487
rect 16500 15484 16528 15580
rect 16669 15487 16727 15493
rect 16669 15484 16681 15487
rect 16500 15456 16681 15484
rect 16301 15447 16359 15453
rect 16669 15453 16681 15456
rect 16715 15453 16727 15487
rect 16776 15484 16804 15648
rect 20438 15512 20444 15564
rect 20496 15552 20502 15564
rect 20714 15552 20720 15564
rect 20496 15524 20720 15552
rect 20496 15512 20502 15524
rect 20714 15512 20720 15524
rect 20772 15552 20778 15564
rect 20772 15524 21036 15552
rect 20772 15512 20778 15524
rect 16853 15487 16911 15493
rect 16853 15484 16865 15487
rect 16776 15456 16865 15484
rect 16669 15447 16727 15453
rect 16853 15453 16865 15456
rect 16899 15453 16911 15487
rect 20530 15484 20536 15496
rect 16853 15447 16911 15453
rect 19996 15456 20536 15484
rect 15841 15419 15899 15425
rect 15841 15416 15853 15419
rect 15212 15388 15853 15416
rect 15105 15379 15163 15385
rect 15841 15385 15853 15388
rect 15887 15416 15899 15419
rect 16316 15416 16344 15447
rect 15887 15388 16344 15416
rect 15887 15385 15899 15388
rect 15841 15379 15899 15385
rect 19996 15360 20024 15456
rect 20530 15444 20536 15456
rect 20588 15484 20594 15496
rect 21008 15493 21036 15524
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 20588 15456 20821 15484
rect 20588 15444 20594 15456
rect 20809 15453 20821 15456
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 12802 15348 12808 15360
rect 11900 15320 12808 15348
rect 12802 15308 12808 15320
rect 12860 15308 12866 15360
rect 13078 15308 13084 15360
rect 13136 15348 13142 15360
rect 13265 15351 13323 15357
rect 13265 15348 13277 15351
rect 13136 15320 13277 15348
rect 13136 15308 13142 15320
rect 13265 15317 13277 15320
rect 13311 15317 13323 15351
rect 13265 15311 13323 15317
rect 16025 15351 16083 15357
rect 16025 15317 16037 15351
rect 16071 15348 16083 15351
rect 16574 15348 16580 15360
rect 16071 15320 16580 15348
rect 16071 15317 16083 15320
rect 16025 15311 16083 15317
rect 16574 15308 16580 15320
rect 16632 15308 16638 15360
rect 16758 15308 16764 15360
rect 16816 15308 16822 15360
rect 19978 15308 19984 15360
rect 20036 15308 20042 15360
rect 1104 15258 35236 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 35236 15258
rect 1104 15184 35236 15206
rect 6730 15104 6736 15156
rect 6788 15104 6794 15156
rect 9490 15104 9496 15156
rect 9548 15144 9554 15156
rect 9548 15116 10824 15144
rect 9548 15104 9554 15116
rect 4338 15036 4344 15088
rect 4396 15036 4402 15088
rect 5074 15036 5080 15088
rect 5132 15036 5138 15088
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 4062 15008 4068 15020
rect 3660 14980 4068 15008
rect 3660 14968 3666 14980
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 6641 15011 6699 15017
rect 6641 14977 6653 15011
rect 6687 15008 6699 15011
rect 6748 15008 6776 15104
rect 6914 15036 6920 15088
rect 6972 15036 6978 15088
rect 8481 15079 8539 15085
rect 8481 15045 8493 15079
rect 8527 15076 8539 15079
rect 8938 15076 8944 15088
rect 8527 15048 8944 15076
rect 8527 15045 8539 15048
rect 8481 15039 8539 15045
rect 8938 15036 8944 15048
rect 8996 15036 9002 15088
rect 9674 15036 9680 15088
rect 9732 15036 9738 15088
rect 9766 15036 9772 15088
rect 9824 15076 9830 15088
rect 10229 15079 10287 15085
rect 10229 15076 10241 15079
rect 9824 15048 10241 15076
rect 9824 15036 9830 15048
rect 10229 15045 10241 15048
rect 10275 15045 10287 15079
rect 10229 15039 10287 15045
rect 10410 15036 10416 15088
rect 10468 15036 10474 15088
rect 10796 15085 10824 15116
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 13814 15144 13820 15156
rect 12584 15116 13820 15144
rect 12584 15104 12590 15116
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 16574 15104 16580 15156
rect 16632 15104 16638 15156
rect 16666 15104 16672 15156
rect 16724 15104 16730 15156
rect 16853 15147 16911 15153
rect 16853 15113 16865 15147
rect 16899 15144 16911 15147
rect 19334 15144 19340 15156
rect 16899 15116 19340 15144
rect 16899 15113 16911 15116
rect 16853 15107 16911 15113
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19705 15147 19763 15153
rect 19705 15144 19717 15147
rect 19484 15116 19717 15144
rect 19484 15104 19490 15116
rect 19705 15113 19717 15116
rect 19751 15113 19763 15147
rect 19705 15107 19763 15113
rect 10781 15079 10839 15085
rect 10781 15045 10793 15079
rect 10827 15045 10839 15079
rect 10781 15039 10839 15045
rect 11238 15036 11244 15088
rect 11296 15036 11302 15088
rect 6918 15033 6976 15036
rect 6687 14980 6776 15008
rect 6825 15011 6883 15017
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 6825 14977 6837 15011
rect 6871 14977 6883 15011
rect 6918 14999 6930 15033
rect 6964 14999 6976 15033
rect 6918 14993 6976 14999
rect 7010 15017 7068 15023
rect 7010 14983 7022 15017
rect 7056 15008 7068 15017
rect 7190 15008 7196 15020
rect 7056 14983 7196 15008
rect 7010 14980 7196 14983
rect 7010 14977 7068 14980
rect 6825 14971 6883 14977
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14909 6147 14943
rect 6089 14903 6147 14909
rect 6104 14804 6132 14903
rect 6840 14884 6868 14971
rect 7190 14968 7196 14980
rect 7248 14968 7254 15020
rect 7650 14940 7656 14952
rect 6932 14912 7656 14940
rect 6822 14832 6828 14884
rect 6880 14832 6886 14884
rect 6546 14804 6552 14816
rect 6104 14776 6552 14804
rect 6546 14764 6552 14776
rect 6604 14804 6610 14816
rect 6932 14804 6960 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7285 14875 7343 14881
rect 7285 14841 7297 14875
rect 7331 14872 7343 14875
rect 7466 14872 7472 14884
rect 7331 14844 7472 14872
rect 7331 14841 7343 14844
rect 7285 14835 7343 14841
rect 7466 14832 7472 14844
rect 7524 14872 7530 14884
rect 7760 14872 7788 14994
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 10597 15011 10655 15017
rect 10597 15008 10609 15011
rect 8720 14980 10609 15008
rect 8720 14968 8726 14980
rect 10597 14977 10609 14980
rect 10643 15008 10655 15011
rect 10686 15008 10692 15020
rect 10643 14980 10692 15008
rect 10643 14977 10655 14980
rect 10597 14971 10655 14977
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 10873 15011 10931 15017
rect 10873 14977 10885 15011
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 8202 14900 8208 14952
rect 8260 14940 8266 14952
rect 9309 14943 9367 14949
rect 9309 14940 9321 14943
rect 8260 14912 9321 14940
rect 8260 14900 8266 14912
rect 9309 14909 9321 14912
rect 9355 14940 9367 14943
rect 9766 14940 9772 14952
rect 9355 14912 9772 14940
rect 9355 14909 9367 14912
rect 9309 14903 9367 14909
rect 9766 14900 9772 14912
rect 9824 14940 9830 14952
rect 10889 14940 10917 14971
rect 10962 14968 10968 15020
rect 11020 15008 11026 15020
rect 11057 15011 11115 15017
rect 11057 15008 11069 15011
rect 11020 14980 11069 15008
rect 11020 14968 11026 14980
rect 11057 14977 11069 14980
rect 11103 15008 11115 15011
rect 12158 15008 12164 15020
rect 11103 14980 12164 15008
rect 11103 14977 11115 14980
rect 11057 14971 11115 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12710 14968 12716 15020
rect 12768 15008 12774 15020
rect 14918 15008 14924 15020
rect 12768 14980 14924 15008
rect 12768 14968 12774 14980
rect 14918 14968 14924 14980
rect 14976 15008 14982 15020
rect 15378 15008 15384 15020
rect 14976 14980 15384 15008
rect 14976 14968 14982 14980
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 14977 15623 15011
rect 16592 15008 16620 15104
rect 16684 15076 16712 15104
rect 16684 15048 16896 15076
rect 16868 15017 16896 15048
rect 19242 15036 19248 15088
rect 19300 15076 19306 15088
rect 19521 15079 19579 15085
rect 19521 15076 19533 15079
rect 19300 15048 19533 15076
rect 19300 15036 19306 15048
rect 19521 15045 19533 15048
rect 19567 15045 19579 15079
rect 19521 15039 19579 15045
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16592 14980 16681 15008
rect 15565 14971 15623 14977
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16853 15011 16911 15017
rect 16853 14977 16865 15011
rect 16899 15008 16911 15011
rect 17313 15011 17371 15017
rect 17313 15008 17325 15011
rect 16899 14980 17325 15008
rect 16899 14977 16911 14980
rect 16853 14971 16911 14977
rect 17313 14977 17325 14980
rect 17359 15008 17371 15011
rect 17957 15011 18015 15017
rect 17957 15008 17969 15011
rect 17359 14980 17969 15008
rect 17359 14977 17371 14980
rect 17313 14971 17371 14977
rect 17957 14977 17969 14980
rect 18003 14977 18015 15011
rect 18877 15011 18935 15017
rect 18877 15008 18889 15011
rect 17957 14971 18015 14977
rect 18064 14980 18889 15008
rect 9824 14912 10917 14940
rect 9824 14900 9830 14912
rect 13446 14900 13452 14952
rect 13504 14940 13510 14952
rect 15286 14940 15292 14952
rect 13504 14912 15292 14940
rect 13504 14900 13510 14912
rect 15286 14900 15292 14912
rect 15344 14940 15350 14952
rect 15580 14940 15608 14971
rect 18064 14952 18092 14980
rect 18877 14977 18889 14980
rect 18923 15008 18935 15011
rect 19337 15011 19395 15017
rect 19337 15008 19349 15011
rect 18923 14980 19349 15008
rect 18923 14977 18935 14980
rect 18877 14971 18935 14977
rect 19337 14977 19349 14980
rect 19383 14977 19395 15011
rect 19337 14971 19395 14977
rect 15344 14912 15608 14940
rect 15344 14900 15350 14912
rect 16758 14900 16764 14952
rect 16816 14940 16822 14952
rect 17221 14943 17279 14949
rect 17221 14940 17233 14943
rect 16816 14912 17233 14940
rect 16816 14900 16822 14912
rect 17221 14909 17233 14912
rect 17267 14940 17279 14943
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 17267 14912 17877 14940
rect 17267 14909 17279 14912
rect 17221 14903 17279 14909
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 18046 14900 18052 14952
rect 18104 14900 18110 14952
rect 18966 14900 18972 14952
rect 19024 14900 19030 14952
rect 19245 14943 19303 14949
rect 19245 14909 19257 14943
rect 19291 14940 19303 14943
rect 20070 14940 20076 14952
rect 19291 14912 20076 14940
rect 19291 14909 19303 14912
rect 19245 14903 19303 14909
rect 20070 14900 20076 14912
rect 20128 14900 20134 14952
rect 7524 14844 7788 14872
rect 7524 14832 7530 14844
rect 10870 14832 10876 14884
rect 10928 14872 10934 14884
rect 11422 14872 11428 14884
rect 10928 14844 11428 14872
rect 10928 14832 10934 14844
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 11974 14832 11980 14884
rect 12032 14872 12038 14884
rect 12894 14872 12900 14884
rect 12032 14844 12900 14872
rect 12032 14832 12038 14844
rect 12894 14832 12900 14844
rect 12952 14832 12958 14884
rect 17681 14875 17739 14881
rect 17681 14841 17693 14875
rect 17727 14872 17739 14875
rect 20346 14872 20352 14884
rect 17727 14844 20352 14872
rect 17727 14841 17739 14844
rect 17681 14835 17739 14841
rect 20346 14832 20352 14844
rect 20404 14872 20410 14884
rect 20990 14872 20996 14884
rect 20404 14844 20996 14872
rect 20404 14832 20410 14844
rect 20990 14832 20996 14844
rect 21048 14832 21054 14884
rect 6604 14776 6960 14804
rect 6604 14764 6610 14776
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 13538 14804 13544 14816
rect 10652 14776 13544 14804
rect 10652 14764 10658 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 15565 14807 15623 14813
rect 15565 14773 15577 14807
rect 15611 14804 15623 14807
rect 15654 14804 15660 14816
rect 15611 14776 15660 14804
rect 15611 14773 15623 14776
rect 15565 14767 15623 14773
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 18230 14764 18236 14816
rect 18288 14764 18294 14816
rect 19334 14764 19340 14816
rect 19392 14804 19398 14816
rect 20438 14804 20444 14816
rect 19392 14776 20444 14804
rect 19392 14764 19398 14776
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 1104 14714 35248 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 35248 14714
rect 1104 14640 35248 14662
rect 4706 14560 4712 14612
rect 4764 14600 4770 14612
rect 4893 14603 4951 14609
rect 4893 14600 4905 14603
rect 4764 14572 4905 14600
rect 4764 14560 4770 14572
rect 4893 14569 4905 14572
rect 4939 14569 4951 14603
rect 4893 14563 4951 14569
rect 4908 14396 4936 14563
rect 5074 14560 5080 14612
rect 5132 14600 5138 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 5132 14572 5181 14600
rect 5132 14560 5138 14572
rect 5169 14569 5181 14572
rect 5215 14569 5227 14603
rect 5169 14563 5227 14569
rect 5258 14560 5264 14612
rect 5316 14600 5322 14612
rect 6086 14600 6092 14612
rect 5316 14572 6092 14600
rect 5316 14560 5322 14572
rect 6086 14560 6092 14572
rect 6144 14600 6150 14612
rect 6822 14600 6828 14612
rect 6144 14572 6828 14600
rect 6144 14560 6150 14572
rect 6822 14560 6828 14572
rect 6880 14560 6886 14612
rect 10042 14560 10048 14612
rect 10100 14600 10106 14612
rect 10962 14600 10968 14612
rect 10100 14572 10968 14600
rect 10100 14560 10106 14572
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11790 14560 11796 14612
rect 11848 14600 11854 14612
rect 12342 14600 12348 14612
rect 11848 14572 12348 14600
rect 11848 14560 11854 14572
rect 12342 14560 12348 14572
rect 12400 14600 12406 14612
rect 12713 14603 12771 14609
rect 12713 14600 12725 14603
rect 12400 14572 12725 14600
rect 12400 14560 12406 14572
rect 12713 14569 12725 14572
rect 12759 14569 12771 14603
rect 12713 14563 12771 14569
rect 13078 14560 13084 14612
rect 13136 14600 13142 14612
rect 13357 14603 13415 14609
rect 13357 14600 13369 14603
rect 13136 14572 13369 14600
rect 13136 14560 13142 14572
rect 13357 14569 13369 14572
rect 13403 14569 13415 14603
rect 13357 14563 13415 14569
rect 13817 14603 13875 14609
rect 13817 14569 13829 14603
rect 13863 14600 13875 14603
rect 14550 14600 14556 14612
rect 13863 14572 14556 14600
rect 13863 14569 13875 14572
rect 13817 14563 13875 14569
rect 14550 14560 14556 14572
rect 14608 14600 14614 14612
rect 15381 14603 15439 14609
rect 15381 14600 15393 14603
rect 14608 14572 15393 14600
rect 14608 14560 14614 14572
rect 15381 14569 15393 14572
rect 15427 14569 15439 14603
rect 15381 14563 15439 14569
rect 15933 14603 15991 14609
rect 15933 14569 15945 14603
rect 15979 14600 15991 14603
rect 18046 14600 18052 14612
rect 15979 14572 18052 14600
rect 15979 14569 15991 14572
rect 15933 14563 15991 14569
rect 18046 14560 18052 14572
rect 18104 14560 18110 14612
rect 18230 14560 18236 14612
rect 18288 14560 18294 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19521 14603 19579 14609
rect 19521 14600 19533 14603
rect 19392 14572 19533 14600
rect 19392 14560 19398 14572
rect 19521 14569 19533 14572
rect 19567 14569 19579 14603
rect 19521 14563 19579 14569
rect 19978 14560 19984 14612
rect 20036 14560 20042 14612
rect 20625 14603 20683 14609
rect 20625 14569 20637 14603
rect 20671 14600 20683 14603
rect 22281 14603 22339 14609
rect 20671 14572 20944 14600
rect 20671 14569 20683 14572
rect 20625 14563 20683 14569
rect 5902 14492 5908 14544
rect 5960 14532 5966 14544
rect 6181 14535 6239 14541
rect 6181 14532 6193 14535
rect 5960 14504 6193 14532
rect 5960 14492 5966 14504
rect 6181 14501 6193 14504
rect 6227 14501 6239 14535
rect 14458 14532 14464 14544
rect 6181 14495 6239 14501
rect 12636 14504 14464 14532
rect 8496 14436 11376 14464
rect 8496 14408 8524 14436
rect 5077 14399 5135 14405
rect 5077 14396 5089 14399
rect 4908 14368 5089 14396
rect 5077 14365 5089 14368
rect 5123 14396 5135 14399
rect 5534 14396 5540 14408
rect 5123 14368 5540 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5534 14356 5540 14368
rect 5592 14396 5598 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 5592 14368 5825 14396
rect 5592 14356 5598 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 5813 14359 5871 14365
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 7101 14399 7159 14405
rect 7101 14365 7113 14399
rect 7147 14396 7159 14399
rect 7190 14396 7196 14408
rect 7147 14368 7196 14396
rect 7147 14365 7159 14368
rect 7101 14359 7159 14365
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 8478 14356 8484 14408
rect 8536 14356 8542 14408
rect 9953 14399 10011 14405
rect 9953 14365 9965 14399
rect 9999 14396 10011 14399
rect 10226 14396 10232 14408
rect 9999 14368 10232 14396
rect 9999 14365 10011 14368
rect 9953 14359 10011 14365
rect 10226 14356 10232 14368
rect 10284 14396 10290 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 10284 14368 10517 14396
rect 10284 14356 10290 14368
rect 10505 14365 10517 14368
rect 10551 14365 10563 14399
rect 10873 14399 10931 14405
rect 10873 14396 10885 14399
rect 10505 14359 10563 14365
rect 10612 14368 10885 14396
rect 6748 14328 6776 14356
rect 7009 14331 7067 14337
rect 7009 14328 7021 14331
rect 6748 14300 7021 14328
rect 7009 14297 7021 14300
rect 7055 14297 7067 14331
rect 7009 14291 7067 14297
rect 7561 14331 7619 14337
rect 7561 14297 7573 14331
rect 7607 14328 7619 14331
rect 7834 14328 7840 14340
rect 7607 14300 7840 14328
rect 7607 14297 7619 14300
rect 7561 14291 7619 14297
rect 7834 14288 7840 14300
rect 7892 14288 7898 14340
rect 10134 14288 10140 14340
rect 10192 14328 10198 14340
rect 10612 14328 10640 14368
rect 10873 14365 10885 14368
rect 10919 14396 10931 14399
rect 10962 14396 10968 14408
rect 10919 14368 10968 14396
rect 10919 14365 10931 14368
rect 10873 14359 10931 14365
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 11054 14356 11060 14408
rect 11112 14396 11118 14408
rect 11149 14399 11207 14405
rect 11149 14396 11161 14399
rect 11112 14368 11161 14396
rect 11112 14356 11118 14368
rect 11149 14365 11161 14368
rect 11195 14396 11207 14399
rect 11238 14396 11244 14408
rect 11195 14368 11244 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11238 14356 11244 14368
rect 11296 14356 11302 14408
rect 11348 14405 11376 14436
rect 12066 14424 12072 14476
rect 12124 14424 12130 14476
rect 12636 14464 12664 14504
rect 14458 14492 14464 14504
rect 14516 14532 14522 14544
rect 14516 14504 15056 14532
rect 14516 14492 14522 14504
rect 12452 14436 12664 14464
rect 11333 14399 11391 14405
rect 11333 14365 11345 14399
rect 11379 14365 11391 14399
rect 11333 14359 11391 14365
rect 10192 14300 10640 14328
rect 10192 14288 10198 14300
rect 10686 14288 10692 14340
rect 10744 14288 10750 14340
rect 10778 14288 10784 14340
rect 10836 14288 10842 14340
rect 11348 14328 11376 14359
rect 11422 14356 11428 14408
rect 11480 14356 11486 14408
rect 11517 14399 11575 14405
rect 11517 14365 11529 14399
rect 11563 14396 11575 14399
rect 11698 14396 11704 14408
rect 11563 14368 11704 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 11974 14356 11980 14408
rect 12032 14356 12038 14408
rect 12158 14356 12164 14408
rect 12216 14396 12222 14408
rect 12253 14399 12311 14405
rect 12253 14396 12265 14399
rect 12216 14368 12265 14396
rect 12216 14356 12222 14368
rect 12253 14365 12265 14368
rect 12299 14365 12311 14399
rect 12253 14359 12311 14365
rect 12342 14356 12348 14408
rect 12400 14356 12406 14408
rect 11348 14300 12388 14328
rect 12360 14294 12388 14300
rect 12452 14294 12480 14436
rect 12710 14424 12716 14476
rect 12768 14464 12774 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12768 14436 12817 14464
rect 12768 14424 12774 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 13446 14424 13452 14476
rect 13504 14424 13510 14476
rect 13538 14424 13544 14476
rect 13596 14464 13602 14476
rect 13596 14436 14872 14464
rect 13596 14424 13602 14436
rect 12526 14356 12532 14408
rect 12584 14356 12590 14408
rect 12894 14356 12900 14408
rect 12952 14396 12958 14408
rect 12989 14399 13047 14405
rect 12989 14396 13001 14399
rect 12952 14368 13001 14396
rect 12952 14356 12958 14368
rect 12989 14365 13001 14368
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13630 14356 13636 14408
rect 13688 14356 13694 14408
rect 13722 14356 13728 14408
rect 13780 14356 13786 14408
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 14844 14405 14872 14436
rect 15028 14405 15056 14504
rect 16390 14492 16396 14544
rect 16448 14492 16454 14544
rect 16132 14436 16344 14464
rect 16132 14408 16160 14436
rect 14829 14399 14887 14405
rect 14829 14365 14841 14399
rect 14875 14365 14887 14399
rect 14829 14359 14887 14365
rect 15013 14399 15071 14405
rect 15013 14365 15025 14399
rect 15059 14365 15071 14399
rect 15286 14396 15292 14408
rect 15013 14359 15071 14365
rect 15120 14368 15292 14396
rect 12544 14328 12572 14356
rect 12713 14331 12771 14337
rect 12713 14328 12725 14331
rect 12544 14300 12725 14328
rect 5442 14220 5448 14272
rect 5500 14220 5506 14272
rect 11057 14263 11115 14269
rect 11057 14229 11069 14263
rect 11103 14260 11115 14263
rect 11514 14260 11520 14272
rect 11103 14232 11520 14260
rect 11103 14229 11115 14232
rect 11057 14223 11115 14229
rect 11514 14220 11520 14232
rect 11572 14220 11578 14272
rect 11701 14263 11759 14269
rect 11701 14229 11713 14263
rect 11747 14260 11759 14263
rect 12250 14260 12256 14272
rect 11747 14232 12256 14260
rect 11747 14229 11759 14232
rect 11701 14223 11759 14229
rect 12250 14220 12256 14232
rect 12308 14220 12314 14272
rect 12360 14266 12480 14294
rect 12713 14297 12725 14300
rect 12759 14328 12771 14331
rect 12802 14328 12808 14340
rect 12759 14300 12808 14328
rect 12759 14297 12771 14300
rect 12713 14291 12771 14297
rect 12802 14288 12808 14300
rect 12860 14288 12866 14340
rect 13354 14288 13360 14340
rect 13412 14328 13418 14340
rect 13740 14328 13768 14356
rect 13412 14300 13768 14328
rect 13412 14288 13418 14300
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14921 14331 14979 14337
rect 14921 14328 14933 14331
rect 13872 14300 14933 14328
rect 13872 14288 13878 14300
rect 14921 14297 14933 14300
rect 14967 14297 14979 14331
rect 14921 14291 14979 14297
rect 12526 14220 12532 14272
rect 12584 14220 12590 14272
rect 13170 14220 13176 14272
rect 13228 14260 13234 14272
rect 15120 14260 15148 14368
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 15808 14399 15866 14405
rect 15808 14365 15820 14399
rect 15854 14396 15866 14399
rect 16114 14396 16120 14408
rect 15854 14368 16120 14396
rect 15854 14365 15866 14368
rect 15808 14359 15866 14365
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 16209 14399 16267 14405
rect 16209 14365 16221 14399
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16224 14328 16252 14359
rect 15212 14300 16252 14328
rect 16316 14328 16344 14436
rect 16408 14405 16436 14492
rect 16393 14399 16451 14405
rect 16393 14365 16405 14399
rect 16439 14365 16451 14399
rect 18248 14396 18276 14560
rect 20714 14492 20720 14544
rect 20772 14492 20778 14544
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19613 14467 19671 14473
rect 19613 14464 19625 14467
rect 19484 14436 19625 14464
rect 19484 14424 19490 14436
rect 19613 14433 19625 14436
rect 19659 14433 19671 14467
rect 20806 14464 20812 14476
rect 19613 14427 19671 14433
rect 20272 14436 20812 14464
rect 20272 14408 20300 14436
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 20916 14464 20944 14572
rect 22281 14569 22293 14603
rect 22327 14600 22339 14603
rect 22462 14600 22468 14612
rect 22327 14572 22468 14600
rect 22327 14569 22339 14572
rect 22281 14563 22339 14569
rect 20916 14436 21312 14464
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 18248 14368 19257 14396
rect 16393 14359 16451 14365
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19334 14356 19340 14408
rect 19392 14356 19398 14408
rect 19705 14399 19763 14405
rect 19705 14365 19717 14399
rect 19751 14365 19763 14399
rect 19705 14359 19763 14365
rect 20165 14399 20223 14405
rect 20165 14365 20177 14399
rect 20211 14396 20223 14399
rect 20254 14396 20260 14408
rect 20211 14368 20260 14396
rect 20211 14365 20223 14368
rect 20165 14359 20223 14365
rect 18782 14328 18788 14340
rect 16316 14300 18788 14328
rect 15212 14269 15240 14300
rect 18782 14288 18788 14300
rect 18840 14288 18846 14340
rect 19352 14328 19380 14356
rect 19720 14328 19748 14359
rect 20254 14356 20260 14368
rect 20312 14356 20318 14408
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20441 14399 20499 14405
rect 20441 14396 20453 14399
rect 20404 14368 20453 14396
rect 20404 14356 20410 14368
rect 20441 14365 20453 14368
rect 20487 14365 20499 14399
rect 20717 14399 20775 14405
rect 20717 14390 20729 14399
rect 20441 14359 20499 14365
rect 20548 14365 20729 14390
rect 20763 14365 20775 14399
rect 20548 14362 20775 14365
rect 20548 14328 20576 14362
rect 20717 14359 20775 14362
rect 20990 14356 20996 14408
rect 21048 14356 21054 14408
rect 21284 14405 21312 14436
rect 22388 14405 22416 14572
rect 22462 14560 22468 14572
rect 22520 14560 22526 14612
rect 22557 14603 22615 14609
rect 22557 14569 22569 14603
rect 22603 14600 22615 14603
rect 22830 14600 22836 14612
rect 22603 14572 22836 14600
rect 22603 14569 22615 14572
rect 22557 14563 22615 14569
rect 22830 14560 22836 14572
rect 22888 14560 22894 14612
rect 22554 14424 22560 14476
rect 22612 14464 22618 14476
rect 22649 14467 22707 14473
rect 22649 14464 22661 14467
rect 22612 14436 22661 14464
rect 22612 14424 22618 14436
rect 22649 14433 22661 14436
rect 22695 14433 22707 14467
rect 22649 14427 22707 14433
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 22373 14399 22431 14405
rect 22373 14365 22385 14399
rect 22419 14365 22431 14399
rect 22373 14359 22431 14365
rect 19352 14300 19748 14328
rect 20272 14300 20576 14328
rect 13228 14232 15148 14260
rect 15197 14263 15255 14269
rect 13228 14220 13234 14232
rect 15197 14229 15209 14263
rect 15243 14229 15255 14263
rect 15197 14223 15255 14229
rect 15746 14220 15752 14272
rect 15804 14220 15810 14272
rect 16393 14263 16451 14269
rect 16393 14229 16405 14263
rect 16439 14260 16451 14263
rect 17034 14260 17040 14272
rect 16439 14232 17040 14260
rect 16439 14229 16451 14232
rect 16393 14223 16451 14229
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 18874 14220 18880 14272
rect 18932 14260 18938 14272
rect 19337 14263 19395 14269
rect 19337 14260 19349 14263
rect 18932 14232 19349 14260
rect 18932 14220 18938 14232
rect 19337 14229 19349 14232
rect 19383 14229 19395 14263
rect 19337 14223 19395 14229
rect 19978 14220 19984 14272
rect 20036 14260 20042 14272
rect 20272 14269 20300 14300
rect 20806 14288 20812 14340
rect 20864 14337 20870 14340
rect 20864 14331 20886 14337
rect 20874 14297 20886 14331
rect 20864 14291 20886 14297
rect 20864 14288 20870 14291
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 20036 14232 20269 14260
rect 20036 14220 20042 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 20714 14220 20720 14272
rect 20772 14260 20778 14272
rect 21100 14260 21128 14359
rect 22462 14356 22468 14408
rect 22520 14356 22526 14408
rect 33134 14356 33140 14408
rect 33192 14356 33198 14408
rect 34333 14331 34391 14337
rect 34333 14297 34345 14331
rect 34379 14328 34391 14331
rect 34882 14328 34888 14340
rect 34379 14300 34888 14328
rect 34379 14297 34391 14300
rect 34333 14291 34391 14297
rect 34882 14288 34888 14300
rect 34940 14288 34946 14340
rect 20772 14232 21128 14260
rect 20772 14220 20778 14232
rect 21266 14220 21272 14272
rect 21324 14220 21330 14272
rect 1104 14170 35236 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 35236 14170
rect 1104 14096 35236 14118
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6362 14056 6368 14068
rect 5960 14028 6368 14056
rect 5960 14016 5966 14028
rect 6362 14016 6368 14028
rect 6420 14056 6426 14068
rect 6549 14059 6607 14065
rect 6549 14056 6561 14059
rect 6420 14028 6561 14056
rect 6420 14016 6426 14028
rect 6549 14025 6561 14028
rect 6595 14025 6607 14059
rect 6549 14019 6607 14025
rect 8938 14016 8944 14068
rect 8996 14016 9002 14068
rect 10134 14016 10140 14068
rect 10192 14056 10198 14068
rect 10192 14028 10732 14056
rect 10192 14016 10198 14028
rect 6086 13948 6092 14000
rect 6144 13948 6150 14000
rect 8956 13988 8984 14016
rect 8956 13960 9674 13988
rect 4062 13880 4068 13932
rect 4120 13880 4126 13932
rect 5442 13880 5448 13932
rect 5500 13880 5506 13932
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 7650 13880 7656 13932
rect 7708 13920 7714 13932
rect 7837 13923 7895 13929
rect 7837 13920 7849 13923
rect 7708 13892 7849 13920
rect 7708 13880 7714 13892
rect 7837 13889 7849 13892
rect 7883 13889 7895 13923
rect 7837 13883 7895 13889
rect 8662 13744 8668 13796
rect 8720 13744 8726 13796
rect 9646 13784 9674 13960
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 10284 13892 10609 13920
rect 10284 13880 10290 13892
rect 10597 13889 10609 13892
rect 10643 13889 10655 13923
rect 10704 13920 10732 14028
rect 12250 14016 12256 14068
rect 12308 14056 12314 14068
rect 13446 14056 13452 14068
rect 12308 14028 13452 14056
rect 12308 14016 12314 14028
rect 13446 14016 13452 14028
rect 13504 14016 13510 14068
rect 15286 14056 15292 14068
rect 13648 14028 14596 14056
rect 13078 13948 13084 14000
rect 13136 13988 13142 14000
rect 13648 13988 13676 14028
rect 14568 14000 14596 14028
rect 14660 14028 15292 14056
rect 13136 13960 13676 13988
rect 13136 13948 13142 13960
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10704 13892 10793 13920
rect 10597 13883 10655 13889
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 10879 13923 10937 13929
rect 10879 13889 10891 13923
rect 10925 13920 10937 13923
rect 10925 13892 11008 13920
rect 10925 13889 10937 13892
rect 10879 13883 10937 13889
rect 10980 13784 11008 13892
rect 11054 13880 11060 13932
rect 11112 13880 11118 13932
rect 13170 13880 13176 13932
rect 13228 13880 13234 13932
rect 13446 13880 13452 13932
rect 13504 13880 13510 13932
rect 13648 13929 13676 13960
rect 14550 13948 14556 14000
rect 14608 13948 14614 14000
rect 14660 13997 14688 14028
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 15746 14016 15752 14068
rect 15804 14016 15810 14068
rect 18874 14016 18880 14068
rect 18932 14016 18938 14068
rect 18966 14016 18972 14068
rect 19024 14056 19030 14068
rect 19061 14059 19119 14065
rect 19061 14056 19073 14059
rect 19024 14028 19073 14056
rect 19024 14016 19030 14028
rect 19061 14025 19073 14028
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 20254 14016 20260 14068
rect 20312 14016 20318 14068
rect 20438 14016 20444 14068
rect 20496 14056 20502 14068
rect 20496 14028 20852 14056
rect 20496 14016 20502 14028
rect 14645 13991 14703 13997
rect 14645 13957 14657 13991
rect 14691 13957 14703 13991
rect 14645 13951 14703 13957
rect 15197 13991 15255 13997
rect 15197 13957 15209 13991
rect 15243 13988 15255 13991
rect 15764 13988 15792 14016
rect 19242 13988 19248 14000
rect 15243 13960 15792 13988
rect 18984 13960 19248 13988
rect 15243 13957 15255 13960
rect 15197 13951 15255 13957
rect 13633 13923 13691 13929
rect 13633 13889 13645 13923
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 13909 13923 13967 13929
rect 13909 13920 13921 13923
rect 13780 13892 13921 13920
rect 13780 13880 13786 13892
rect 13909 13889 13921 13892
rect 13955 13920 13967 13923
rect 14090 13920 14096 13932
rect 13955 13892 14096 13920
rect 13955 13889 13967 13892
rect 13909 13883 13967 13889
rect 14090 13880 14096 13892
rect 14148 13880 14154 13932
rect 14277 13923 14335 13929
rect 14277 13889 14289 13923
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 13078 13812 13084 13864
rect 13136 13812 13142 13864
rect 14292 13852 14320 13883
rect 14366 13880 14372 13932
rect 14424 13880 14430 13932
rect 14660 13852 14688 13951
rect 14737 13923 14795 13929
rect 14737 13889 14749 13923
rect 14783 13889 14795 13923
rect 14737 13883 14795 13889
rect 14292 13824 14688 13852
rect 11698 13784 11704 13796
rect 9646 13756 11704 13784
rect 11698 13744 11704 13756
rect 11756 13744 11762 13796
rect 12710 13744 12716 13796
rect 12768 13784 12774 13796
rect 13354 13784 13360 13796
rect 12768 13756 13360 13784
rect 12768 13744 12774 13756
rect 13354 13744 13360 13756
rect 13412 13784 13418 13796
rect 13412 13756 14044 13784
rect 13412 13744 13418 13756
rect 4328 13719 4386 13725
rect 4328 13685 4340 13719
rect 4374 13716 4386 13719
rect 4706 13716 4712 13728
rect 4374 13688 4712 13716
rect 4374 13685 4386 13688
rect 4328 13679 4386 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 10686 13676 10692 13728
rect 10744 13676 10750 13728
rect 10965 13719 11023 13725
rect 10965 13685 10977 13719
rect 11011 13716 11023 13719
rect 11974 13716 11980 13728
rect 11011 13688 11980 13716
rect 11011 13685 11023 13688
rect 10965 13679 11023 13685
rect 11974 13676 11980 13688
rect 12032 13676 12038 13728
rect 12342 13676 12348 13728
rect 12400 13676 12406 13728
rect 12894 13676 12900 13728
rect 12952 13676 12958 13728
rect 13906 13676 13912 13728
rect 13964 13676 13970 13728
rect 14016 13716 14044 13756
rect 14090 13744 14096 13796
rect 14148 13784 14154 13796
rect 14752 13784 14780 13883
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15160 13892 15301 13920
rect 15160 13880 15166 13892
rect 15289 13889 15301 13892
rect 15335 13889 15347 13923
rect 15289 13883 15347 13889
rect 15565 13923 15623 13929
rect 15565 13889 15577 13923
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 15580 13852 15608 13883
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 17954 13920 17960 13932
rect 15712 13892 17960 13920
rect 15712 13880 15718 13892
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 18785 13923 18843 13929
rect 18785 13920 18797 13923
rect 18064 13892 18797 13920
rect 18064 13864 18092 13892
rect 18785 13889 18797 13892
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 15580 13824 16344 13852
rect 15381 13787 15439 13793
rect 15381 13784 15393 13787
rect 14148 13756 14780 13784
rect 14844 13756 15393 13784
rect 14148 13744 14154 13756
rect 14844 13716 14872 13756
rect 15381 13753 15393 13756
rect 15427 13753 15439 13787
rect 15381 13747 15439 13753
rect 16316 13728 16344 13824
rect 18046 13812 18052 13864
rect 18104 13812 18110 13864
rect 18800 13852 18828 13883
rect 18874 13880 18880 13932
rect 18932 13920 18938 13932
rect 18984 13929 19012 13960
rect 19242 13948 19248 13960
rect 19300 13988 19306 14000
rect 19705 13991 19763 13997
rect 19705 13988 19717 13991
rect 19300 13960 19717 13988
rect 19300 13948 19306 13960
rect 19705 13957 19717 13960
rect 19751 13988 19763 13991
rect 19889 13991 19947 13997
rect 19889 13988 19901 13991
rect 19751 13960 19901 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 19889 13957 19901 13960
rect 19935 13957 19947 13991
rect 20533 13991 20591 13997
rect 20533 13988 20545 13991
rect 19889 13951 19947 13957
rect 20088 13960 20545 13988
rect 18969 13923 19027 13929
rect 18969 13920 18981 13923
rect 18932 13892 18981 13920
rect 18932 13880 18938 13892
rect 18969 13889 18981 13892
rect 19015 13889 19027 13923
rect 19610 13920 19616 13932
rect 18969 13883 19027 13889
rect 19260 13892 19616 13920
rect 19260 13861 19288 13892
rect 19610 13880 19616 13892
rect 19668 13920 19674 13932
rect 20088 13929 20116 13960
rect 20533 13957 20545 13960
rect 20579 13957 20591 13991
rect 20533 13951 20591 13957
rect 20824 13988 20852 14028
rect 21266 14016 21272 14068
rect 21324 14016 21330 14068
rect 22462 14016 22468 14068
rect 22520 14016 22526 14068
rect 23661 14059 23719 14065
rect 23661 14025 23673 14059
rect 23707 14056 23719 14059
rect 24118 14056 24124 14068
rect 23707 14028 24124 14056
rect 23707 14025 23719 14028
rect 23661 14019 23719 14025
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 25501 14059 25559 14065
rect 25501 14025 25513 14059
rect 25547 14056 25559 14059
rect 33134 14056 33140 14068
rect 25547 14028 33140 14056
rect 25547 14025 25559 14028
rect 25501 14019 25559 14025
rect 33134 14016 33140 14028
rect 33192 14016 33198 14068
rect 21284 13988 21312 14016
rect 20824 13960 21220 13988
rect 21284 13960 21956 13988
rect 20824 13929 20852 13960
rect 21192 13929 21220 13960
rect 19797 13923 19855 13929
rect 19797 13920 19809 13923
rect 19668 13892 19809 13920
rect 19668 13880 19674 13892
rect 19797 13889 19809 13892
rect 19843 13889 19855 13923
rect 20073 13923 20131 13929
rect 20073 13920 20085 13923
rect 19797 13883 19855 13889
rect 19996 13892 20085 13920
rect 19245 13855 19303 13861
rect 19245 13852 19257 13855
rect 18800 13824 19257 13852
rect 19245 13821 19257 13824
rect 19291 13821 19303 13855
rect 19245 13815 19303 13821
rect 19337 13855 19395 13861
rect 19337 13821 19349 13855
rect 19383 13852 19395 13855
rect 19426 13852 19432 13864
rect 19383 13824 19432 13852
rect 19383 13821 19395 13824
rect 19337 13815 19395 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19444 13784 19472 13812
rect 19996 13784 20024 13892
rect 20073 13889 20085 13892
rect 20119 13889 20131 13923
rect 20349 13923 20407 13929
rect 20349 13920 20361 13923
rect 20073 13883 20131 13889
rect 20180 13892 20361 13920
rect 19444 13756 20024 13784
rect 14016 13688 14872 13716
rect 14918 13676 14924 13728
rect 14976 13676 14982 13728
rect 16298 13676 16304 13728
rect 16356 13676 16362 13728
rect 19334 13676 19340 13728
rect 19392 13716 19398 13728
rect 20180 13716 20208 13892
rect 20349 13889 20361 13892
rect 20395 13889 20407 13923
rect 20349 13883 20407 13889
rect 20809 13923 20867 13929
rect 20809 13889 20821 13923
rect 20855 13889 20867 13923
rect 20809 13883 20867 13889
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13889 21051 13923
rect 20993 13883 21051 13889
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 20717 13855 20775 13861
rect 20717 13821 20729 13855
rect 20763 13852 20775 13855
rect 21008 13852 21036 13883
rect 21284 13852 21312 13883
rect 21928 13861 21956 13960
rect 22005 13923 22063 13929
rect 22005 13889 22017 13923
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 20763 13824 21312 13852
rect 21913 13855 21971 13861
rect 20763 13821 20775 13824
rect 20717 13815 20775 13821
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 20993 13787 21051 13793
rect 20993 13753 21005 13787
rect 21039 13784 21051 13787
rect 21726 13784 21732 13796
rect 21039 13756 21732 13784
rect 21039 13753 21051 13756
rect 20993 13747 21051 13753
rect 21726 13744 21732 13756
rect 21784 13784 21790 13796
rect 22020 13784 22048 13883
rect 22373 13855 22431 13861
rect 22373 13821 22385 13855
rect 22419 13852 22431 13855
rect 22480 13852 22508 14016
rect 24029 13991 24087 13997
rect 24029 13988 24041 13991
rect 23124 13960 24041 13988
rect 22554 13880 22560 13932
rect 22612 13920 22618 13932
rect 22741 13923 22799 13929
rect 22741 13920 22753 13923
rect 22612 13892 22753 13920
rect 22612 13880 22618 13892
rect 22741 13889 22753 13892
rect 22787 13889 22799 13923
rect 22741 13883 22799 13889
rect 23124 13861 23152 13960
rect 24029 13957 24041 13960
rect 24075 13957 24087 13991
rect 25685 13991 25743 13997
rect 25685 13988 25697 13991
rect 25254 13960 25697 13988
rect 24029 13951 24087 13957
rect 25685 13957 25697 13960
rect 25731 13957 25743 13991
rect 25685 13951 25743 13957
rect 26050 13948 26056 14000
rect 26108 13948 26114 14000
rect 25777 13923 25835 13929
rect 25777 13889 25789 13923
rect 25823 13920 25835 13923
rect 26068 13920 26096 13948
rect 25823 13892 26096 13920
rect 25823 13889 25835 13892
rect 25777 13883 25835 13889
rect 22649 13855 22707 13861
rect 22649 13852 22661 13855
rect 22419 13824 22661 13852
rect 22419 13821 22431 13824
rect 22373 13815 22431 13821
rect 22649 13821 22661 13824
rect 22695 13821 22707 13855
rect 22649 13815 22707 13821
rect 23109 13855 23167 13861
rect 23109 13821 23121 13855
rect 23155 13821 23167 13855
rect 23109 13815 23167 13821
rect 23474 13812 23480 13864
rect 23532 13852 23538 13864
rect 23753 13855 23811 13861
rect 23753 13852 23765 13855
rect 23532 13824 23765 13852
rect 23532 13812 23538 13824
rect 23753 13821 23765 13824
rect 23799 13852 23811 13855
rect 24118 13852 24124 13864
rect 23799 13824 24124 13852
rect 23799 13821 23811 13824
rect 23753 13815 23811 13821
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 25038 13812 25044 13864
rect 25096 13852 25102 13864
rect 25792 13852 25820 13883
rect 25096 13824 25820 13852
rect 25096 13812 25102 13824
rect 21784 13756 22048 13784
rect 21784 13744 21790 13756
rect 19392 13688 20208 13716
rect 19392 13676 19398 13688
rect 21450 13676 21456 13728
rect 21508 13676 21514 13728
rect 1104 13626 35248 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 35248 13626
rect 1104 13552 35248 13574
rect 6362 13472 6368 13524
rect 6420 13472 6426 13524
rect 8386 13472 8392 13524
rect 8444 13472 8450 13524
rect 11793 13515 11851 13521
rect 11793 13512 11805 13515
rect 9646 13484 11805 13512
rect 8404 13444 8432 13472
rect 9646 13444 9674 13484
rect 11793 13481 11805 13484
rect 11839 13512 11851 13515
rect 12066 13512 12072 13524
rect 11839 13484 12072 13512
rect 11839 13481 11851 13484
rect 11793 13475 11851 13481
rect 12066 13472 12072 13484
rect 12124 13512 12130 13524
rect 12618 13512 12624 13524
rect 12124 13484 12624 13512
rect 12124 13472 12130 13484
rect 12618 13472 12624 13484
rect 12676 13472 12682 13524
rect 12710 13472 12716 13524
rect 12768 13472 12774 13524
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 13173 13515 13231 13521
rect 13173 13512 13185 13515
rect 12860 13484 13185 13512
rect 12860 13472 12866 13484
rect 13173 13481 13185 13484
rect 13219 13481 13231 13515
rect 13173 13475 13231 13481
rect 17954 13472 17960 13524
rect 18012 13472 18018 13524
rect 18969 13515 19027 13521
rect 18969 13481 18981 13515
rect 19015 13512 19027 13515
rect 19334 13512 19340 13524
rect 19015 13484 19340 13512
rect 19015 13481 19027 13484
rect 18969 13475 19027 13481
rect 19334 13472 19340 13484
rect 19392 13472 19398 13524
rect 19426 13472 19432 13524
rect 19484 13512 19490 13524
rect 19613 13515 19671 13521
rect 19613 13512 19625 13515
rect 19484 13484 19625 13512
rect 19484 13472 19490 13484
rect 19613 13481 19625 13484
rect 19659 13481 19671 13515
rect 19613 13475 19671 13481
rect 8404 13416 9674 13444
rect 11701 13447 11759 13453
rect 11701 13413 11713 13447
rect 11747 13413 11759 13447
rect 11701 13407 11759 13413
rect 11885 13447 11943 13453
rect 11885 13413 11897 13447
rect 11931 13444 11943 13447
rect 12342 13444 12348 13456
rect 11931 13416 12348 13444
rect 11931 13413 11943 13416
rect 11885 13407 11943 13413
rect 4062 13336 4068 13388
rect 4120 13336 4126 13388
rect 11716 13376 11744 13407
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 12989 13447 13047 13453
rect 12989 13413 13001 13447
rect 13035 13444 13047 13447
rect 13722 13444 13728 13456
rect 13035 13416 13728 13444
rect 13035 13413 13047 13416
rect 12989 13407 13047 13413
rect 13722 13404 13728 13416
rect 13780 13444 13786 13456
rect 13780 13416 14320 13444
rect 13780 13404 13786 13416
rect 11790 13376 11796 13388
rect 11716 13348 11796 13376
rect 11790 13336 11796 13348
rect 11848 13376 11854 13388
rect 11848 13348 12572 13376
rect 11848 13336 11854 13348
rect 934 13268 940 13320
rect 992 13308 998 13320
rect 1397 13311 1455 13317
rect 1397 13308 1409 13311
rect 992 13280 1409 13308
rect 992 13268 998 13280
rect 1397 13277 1409 13280
rect 1443 13277 1455 13311
rect 1397 13271 1455 13277
rect 6089 13311 6147 13317
rect 6089 13277 6101 13311
rect 6135 13308 6147 13311
rect 7098 13308 7104 13320
rect 6135 13280 7104 13308
rect 6135 13277 6147 13280
rect 6089 13271 6147 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7282 13268 7288 13320
rect 7340 13268 7346 13320
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7892 13280 7941 13308
rect 7892 13268 7898 13280
rect 7929 13277 7941 13280
rect 7975 13277 7987 13311
rect 7929 13271 7987 13277
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 11974 13268 11980 13320
rect 12032 13268 12038 13320
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 12437 13311 12495 13317
rect 12437 13308 12449 13311
rect 12207 13280 12449 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12437 13277 12449 13280
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 4341 13243 4399 13249
rect 4341 13240 4353 13243
rect 2746 13212 4353 13240
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13172 1639 13175
rect 2746 13172 2774 13212
rect 4341 13209 4353 13212
rect 4387 13209 4399 13243
rect 4341 13203 4399 13209
rect 5074 13200 5080 13252
rect 5132 13200 5138 13252
rect 10704 13240 10732 13268
rect 11698 13240 11704 13252
rect 10704 13212 11704 13240
rect 11698 13200 11704 13212
rect 11756 13240 11762 13252
rect 12176 13240 12204 13271
rect 11756 13212 12204 13240
rect 12544 13240 12572 13348
rect 12618 13336 12624 13388
rect 12676 13336 12682 13388
rect 12802 13336 12808 13388
rect 12860 13376 12866 13388
rect 12860 13348 13124 13376
rect 12860 13336 12866 13348
rect 12636 13308 12664 13336
rect 12713 13311 12771 13317
rect 12713 13308 12725 13311
rect 12636 13280 12725 13308
rect 12713 13277 12725 13280
rect 12759 13308 12771 13311
rect 12986 13308 12992 13320
rect 12759 13280 12992 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 12986 13268 12992 13280
rect 13044 13268 13050 13320
rect 13096 13317 13124 13348
rect 13081 13311 13139 13317
rect 13081 13277 13093 13311
rect 13127 13277 13139 13311
rect 13081 13271 13139 13277
rect 13357 13311 13415 13317
rect 13357 13277 13369 13311
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13372 13240 13400 13271
rect 14090 13268 14096 13320
rect 14148 13268 14154 13320
rect 14292 13317 14320 13416
rect 17972 13376 18000 13472
rect 18233 13447 18291 13453
rect 18233 13413 18245 13447
rect 18279 13444 18291 13447
rect 18874 13444 18880 13456
rect 18279 13416 18880 13444
rect 18279 13413 18291 13416
rect 18233 13407 18291 13413
rect 18874 13404 18880 13416
rect 18932 13444 18938 13456
rect 18932 13416 19564 13444
rect 18932 13404 18938 13416
rect 19245 13379 19303 13385
rect 19245 13376 19257 13379
rect 17972 13348 19257 13376
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13277 14335 13311
rect 14277 13271 14335 13277
rect 14369 13311 14427 13317
rect 14369 13277 14381 13311
rect 14415 13277 14427 13311
rect 14369 13271 14427 13277
rect 14384 13240 14412 13271
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17589 13311 17647 13317
rect 17589 13308 17601 13311
rect 17092 13280 17601 13308
rect 17092 13268 17098 13280
rect 17589 13277 17601 13280
rect 17635 13277 17647 13311
rect 17589 13271 17647 13277
rect 17773 13311 17831 13317
rect 17773 13277 17785 13311
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 12544 13212 13400 13240
rect 13648 13212 14412 13240
rect 17788 13240 17816 13271
rect 17954 13268 17960 13320
rect 18012 13268 18018 13320
rect 18800 13317 18828 13348
rect 19245 13345 19257 13348
rect 19291 13345 19303 13379
rect 19245 13339 19303 13345
rect 18785 13311 18843 13317
rect 18785 13277 18797 13311
rect 18831 13277 18843 13311
rect 18785 13271 18843 13277
rect 18969 13311 19027 13317
rect 18969 13277 18981 13311
rect 19015 13277 19027 13311
rect 18969 13271 19027 13277
rect 19429 13311 19487 13317
rect 19429 13277 19441 13311
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 18984 13240 19012 13271
rect 19444 13240 19472 13271
rect 17788 13212 17908 13240
rect 11756 13200 11762 13212
rect 1627 13144 2774 13172
rect 11425 13175 11483 13181
rect 1627 13141 1639 13144
rect 1581 13135 1639 13141
rect 11425 13141 11437 13175
rect 11471 13172 11483 13175
rect 11514 13172 11520 13184
rect 11471 13144 11520 13172
rect 11471 13141 11483 13144
rect 11425 13135 11483 13141
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 13538 13132 13544 13184
rect 13596 13172 13602 13184
rect 13648 13181 13676 13212
rect 17880 13184 17908 13212
rect 18616 13212 19472 13240
rect 19536 13240 19564 13416
rect 19628 13376 19656 13475
rect 19978 13472 19984 13524
rect 20036 13472 20042 13524
rect 22373 13515 22431 13521
rect 22373 13481 22385 13515
rect 22419 13512 22431 13515
rect 22554 13512 22560 13524
rect 22419 13484 22560 13512
rect 22419 13481 22431 13484
rect 22373 13475 22431 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 22646 13472 22652 13524
rect 22704 13472 22710 13524
rect 21637 13379 21695 13385
rect 19628 13348 20024 13376
rect 19610 13268 19616 13320
rect 19668 13308 19674 13320
rect 19996 13317 20024 13348
rect 21637 13345 21649 13379
rect 21683 13376 21695 13379
rect 21683 13348 22140 13376
rect 21683 13345 21695 13348
rect 21637 13339 21695 13345
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19668 13280 19717 13308
rect 19668 13268 19674 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 19981 13311 20039 13317
rect 19981 13277 19993 13311
rect 20027 13277 20039 13311
rect 19981 13271 20039 13277
rect 21450 13268 21456 13320
rect 21508 13308 21514 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 21508 13280 21557 13308
rect 21508 13268 21514 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 22112 13317 22140 13348
rect 22097 13311 22155 13317
rect 22097 13277 22109 13311
rect 22143 13277 22155 13311
rect 22097 13271 22155 13277
rect 19889 13243 19947 13249
rect 19889 13240 19901 13243
rect 19536 13212 19901 13240
rect 18616 13184 18644 13212
rect 19889 13209 19901 13212
rect 19935 13209 19947 13243
rect 19889 13203 19947 13209
rect 22112 13184 22140 13271
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22664 13308 22692 13472
rect 22244 13280 22692 13308
rect 22244 13268 22250 13280
rect 22373 13243 22431 13249
rect 22373 13209 22385 13243
rect 22419 13240 22431 13243
rect 22462 13240 22468 13252
rect 22419 13212 22468 13240
rect 22419 13209 22431 13212
rect 22373 13203 22431 13209
rect 22462 13200 22468 13212
rect 22520 13200 22526 13252
rect 13633 13175 13691 13181
rect 13633 13172 13645 13175
rect 13596 13144 13645 13172
rect 13596 13132 13602 13144
rect 13633 13141 13645 13144
rect 13679 13141 13691 13175
rect 13633 13135 13691 13141
rect 13998 13132 14004 13184
rect 14056 13172 14062 13184
rect 16022 13172 16028 13184
rect 14056 13144 16028 13172
rect 14056 13132 14062 13144
rect 16022 13132 16028 13144
rect 16080 13132 16086 13184
rect 17862 13132 17868 13184
rect 17920 13132 17926 13184
rect 18598 13132 18604 13184
rect 18656 13132 18662 13184
rect 22094 13132 22100 13184
rect 22152 13132 22158 13184
rect 1104 13082 35236 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 35236 13082
rect 1104 13008 35236 13030
rect 5074 12928 5080 12980
rect 5132 12968 5138 12980
rect 5169 12971 5227 12977
rect 5169 12968 5181 12971
rect 5132 12940 5181 12968
rect 5132 12928 5138 12940
rect 5169 12937 5181 12940
rect 5215 12937 5227 12971
rect 5169 12931 5227 12937
rect 5534 12928 5540 12980
rect 5592 12928 5598 12980
rect 10413 12971 10471 12977
rect 10413 12937 10425 12971
rect 10459 12968 10471 12971
rect 11241 12971 11299 12977
rect 10459 12940 11100 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12832 5135 12835
rect 5552 12832 5580 12928
rect 10321 12903 10379 12909
rect 10321 12900 10333 12903
rect 8786 12872 10333 12900
rect 10321 12869 10333 12872
rect 10367 12900 10379 12903
rect 10778 12900 10784 12912
rect 10367 12872 10784 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 10778 12860 10784 12872
rect 10836 12900 10842 12912
rect 10836 12872 11008 12900
rect 10836 12860 10842 12872
rect 5123 12804 5580 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 7282 12792 7288 12844
rect 7340 12792 7346 12844
rect 7834 12792 7840 12844
rect 7892 12792 7898 12844
rect 10226 12792 10232 12844
rect 10284 12792 10290 12844
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12733 10839 12767
rect 10781 12727 10839 12733
rect 10042 12656 10048 12708
rect 10100 12656 10106 12708
rect 10796 12696 10824 12727
rect 10870 12724 10876 12776
rect 10928 12724 10934 12776
rect 10980 12773 11008 12872
rect 11072 12773 11100 12940
rect 11241 12937 11253 12971
rect 11287 12937 11299 12971
rect 11241 12931 11299 12937
rect 11256 12844 11284 12931
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12894 12928 12900 12980
rect 12952 12928 12958 12980
rect 13998 12968 14004 12980
rect 13096 12940 14004 12968
rect 11992 12900 12020 12928
rect 12802 12900 12808 12912
rect 11532 12872 12808 12900
rect 11238 12792 11244 12844
rect 11296 12792 11302 12844
rect 11532 12841 11560 12872
rect 11517 12835 11575 12841
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 12084 12841 12112 12872
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 12912 12900 12940 12928
rect 13096 12909 13124 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14090 12928 14096 12980
rect 14148 12928 14154 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 14200 12940 14657 12968
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 12912 12872 13001 12900
rect 12989 12869 13001 12872
rect 13035 12869 13047 12903
rect 12989 12863 13047 12869
rect 13081 12903 13139 12909
rect 13081 12869 13093 12903
rect 13127 12869 13139 12903
rect 14108 12900 14136 12928
rect 13081 12863 13139 12869
rect 13740 12872 14136 12900
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12253 12835 12311 12841
rect 12253 12801 12265 12835
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 13357 12835 13415 12841
rect 13357 12801 13369 12835
rect 13403 12832 13415 12835
rect 13633 12835 13691 12841
rect 13633 12832 13645 12835
rect 13403 12804 13645 12832
rect 13403 12801 13415 12804
rect 13357 12795 13415 12801
rect 13633 12801 13645 12804
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 10965 12767 11023 12773
rect 10965 12733 10977 12767
rect 11011 12733 11023 12767
rect 10965 12727 11023 12733
rect 11057 12767 11115 12773
rect 11057 12733 11069 12767
rect 11103 12764 11115 12767
rect 11330 12764 11336 12776
rect 11103 12736 11336 12764
rect 11103 12733 11115 12736
rect 11057 12727 11115 12733
rect 11330 12724 11336 12736
rect 11388 12724 11394 12776
rect 11716 12764 11744 12792
rect 12268 12764 12296 12795
rect 11716 12736 12296 12764
rect 13541 12767 13599 12773
rect 13541 12733 13553 12767
rect 13587 12764 13599 12767
rect 13740 12764 13768 12872
rect 13817 12835 13875 12841
rect 13817 12801 13829 12835
rect 13863 12832 13875 12835
rect 13906 12832 13912 12844
rect 13863 12804 13912 12832
rect 13863 12801 13875 12804
rect 13817 12795 13875 12801
rect 13906 12792 13912 12804
rect 13964 12832 13970 12844
rect 14200 12832 14228 12940
rect 14645 12937 14657 12940
rect 14691 12937 14703 12971
rect 14645 12931 14703 12937
rect 14918 12928 14924 12980
rect 14976 12928 14982 12980
rect 16224 12940 16988 12968
rect 14936 12900 14964 12928
rect 14568 12872 14964 12900
rect 14568 12844 14596 12872
rect 16022 12860 16028 12912
rect 16080 12900 16086 12912
rect 16224 12900 16252 12940
rect 16080 12872 16252 12900
rect 16316 12872 16896 12900
rect 16080 12860 16086 12872
rect 13964 12804 14228 12832
rect 13964 12792 13970 12804
rect 14366 12792 14372 12844
rect 14424 12792 14430 12844
rect 14550 12792 14556 12844
rect 14608 12792 14614 12844
rect 14829 12835 14887 12841
rect 14829 12801 14841 12835
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 13587 12736 13768 12764
rect 14093 12767 14151 12773
rect 13587 12733 13599 12736
rect 13541 12727 13599 12733
rect 14093 12733 14105 12767
rect 14139 12733 14151 12767
rect 14384 12764 14412 12792
rect 14844 12764 14872 12795
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 16316 12841 16344 12872
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 14976 12804 15669 12832
rect 14976 12792 14982 12804
rect 15657 12801 15669 12804
rect 15703 12832 15715 12835
rect 16209 12835 16267 12841
rect 16209 12832 16221 12835
rect 15703 12830 15976 12832
rect 16132 12830 16221 12832
rect 15703 12804 16221 12830
rect 15703 12801 15715 12804
rect 15948 12802 16160 12804
rect 15657 12795 15715 12801
rect 16209 12801 16221 12804
rect 16255 12801 16267 12835
rect 16209 12795 16267 12801
rect 16301 12835 16359 12841
rect 16301 12801 16313 12835
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 16666 12792 16672 12844
rect 16724 12792 16730 12844
rect 16868 12841 16896 12872
rect 16960 12844 16988 12940
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17313 12971 17371 12977
rect 17313 12968 17325 12971
rect 17092 12940 17325 12968
rect 17092 12928 17098 12940
rect 17313 12937 17325 12940
rect 17359 12937 17371 12971
rect 17313 12931 17371 12937
rect 17957 12971 18015 12977
rect 17957 12937 17969 12971
rect 18003 12968 18015 12971
rect 18046 12968 18052 12980
rect 18003 12940 18052 12968
rect 18003 12937 18015 12940
rect 17957 12931 18015 12937
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 17126 12860 17132 12912
rect 17184 12900 17190 12912
rect 17184 12872 18368 12900
rect 17184 12860 17190 12872
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 14384 12736 14872 12764
rect 15013 12767 15071 12773
rect 14093 12727 14151 12733
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 16574 12764 16580 12776
rect 15059 12736 16580 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 11609 12699 11667 12705
rect 11609 12696 11621 12699
rect 10796 12668 11621 12696
rect 11609 12665 11621 12668
rect 11655 12665 11667 12699
rect 14108 12696 14136 12727
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 16868 12764 16896 12795
rect 16942 12792 16948 12844
rect 17000 12792 17006 12844
rect 17034 12792 17040 12844
rect 17092 12792 17098 12844
rect 17221 12835 17279 12841
rect 17221 12801 17233 12835
rect 17267 12832 17279 12835
rect 17494 12832 17500 12844
rect 17267 12804 17500 12832
rect 17267 12801 17279 12804
rect 17221 12795 17279 12801
rect 17494 12792 17500 12804
rect 17552 12832 17558 12844
rect 18233 12835 18291 12841
rect 18233 12832 18245 12835
rect 17552 12804 18245 12832
rect 17552 12792 17558 12804
rect 18233 12801 18245 12804
rect 18279 12801 18291 12835
rect 18233 12795 18291 12801
rect 17052 12764 17080 12792
rect 16868 12736 17080 12764
rect 17681 12767 17739 12773
rect 17681 12733 17693 12767
rect 17727 12733 17739 12767
rect 17681 12727 17739 12733
rect 17773 12767 17831 12773
rect 17773 12733 17785 12767
rect 17819 12764 17831 12767
rect 17862 12764 17868 12776
rect 17819 12736 17868 12764
rect 17819 12733 17831 12736
rect 17773 12727 17831 12733
rect 11609 12659 11667 12665
rect 13556 12668 14136 12696
rect 13556 12640 13584 12668
rect 16114 12656 16120 12708
rect 16172 12656 16178 12708
rect 17221 12699 17279 12705
rect 17221 12665 17233 12699
rect 17267 12696 17279 12699
rect 17696 12696 17724 12727
rect 17862 12724 17868 12736
rect 17920 12724 17926 12776
rect 17954 12724 17960 12776
rect 18012 12724 18018 12776
rect 18340 12773 18368 12872
rect 22281 12835 22339 12841
rect 22281 12801 22293 12835
rect 22327 12832 22339 12835
rect 22462 12832 22468 12844
rect 22327 12804 22468 12832
rect 22327 12801 22339 12804
rect 22281 12795 22339 12801
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12733 18383 12767
rect 18325 12727 18383 12733
rect 18598 12724 18604 12776
rect 18656 12724 18662 12776
rect 22094 12724 22100 12776
rect 22152 12764 22158 12776
rect 22189 12767 22247 12773
rect 22189 12764 22201 12767
rect 22152 12736 22201 12764
rect 22152 12724 22158 12736
rect 22189 12733 22201 12736
rect 22235 12733 22247 12767
rect 22189 12727 22247 12733
rect 17972 12696 18000 12724
rect 17267 12668 18000 12696
rect 17267 12665 17279 12668
rect 17221 12659 17279 12665
rect 10597 12631 10655 12637
rect 10597 12597 10609 12631
rect 10643 12628 10655 12631
rect 12158 12628 12164 12640
rect 10643 12600 12164 12628
rect 10643 12597 10655 12600
rect 10597 12591 10655 12597
rect 12158 12588 12164 12600
rect 12216 12588 12222 12640
rect 12253 12631 12311 12637
rect 12253 12597 12265 12631
rect 12299 12628 12311 12631
rect 12434 12628 12440 12640
rect 12299 12600 12440 12628
rect 12299 12597 12311 12600
rect 12253 12591 12311 12597
rect 12434 12588 12440 12600
rect 12492 12588 12498 12640
rect 13538 12588 13544 12640
rect 13596 12588 13602 12640
rect 13722 12588 13728 12640
rect 13780 12628 13786 12640
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 13780 12600 14013 12628
rect 13780 12588 13786 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 14001 12591 14059 12597
rect 15746 12588 15752 12640
rect 15804 12588 15810 12640
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 22649 12631 22707 12637
rect 22649 12597 22661 12631
rect 22695 12628 22707 12631
rect 23566 12628 23572 12640
rect 22695 12600 23572 12628
rect 22695 12597 22707 12600
rect 22649 12591 22707 12597
rect 23566 12588 23572 12600
rect 23624 12588 23630 12640
rect 1104 12538 35248 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 35248 12538
rect 1104 12464 35248 12486
rect 6178 12384 6184 12436
rect 6236 12424 6242 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 6236 12396 6469 12424
rect 6236 12384 6242 12396
rect 6457 12393 6469 12396
rect 6503 12393 6515 12427
rect 6457 12387 6515 12393
rect 10781 12427 10839 12433
rect 10781 12393 10793 12427
rect 10827 12424 10839 12427
rect 10870 12424 10876 12436
rect 10827 12396 10876 12424
rect 10827 12393 10839 12396
rect 10781 12387 10839 12393
rect 10870 12384 10876 12396
rect 10928 12384 10934 12436
rect 11333 12427 11391 12433
rect 11333 12393 11345 12427
rect 11379 12424 11391 12427
rect 11882 12424 11888 12436
rect 11379 12396 11888 12424
rect 11379 12393 11391 12396
rect 11333 12387 11391 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 12158 12384 12164 12436
rect 12216 12384 12222 12436
rect 14918 12424 14924 12436
rect 12728 12396 14924 12424
rect 3878 12248 3884 12300
rect 3936 12288 3942 12300
rect 4157 12291 4215 12297
rect 4157 12288 4169 12291
rect 3936 12260 4169 12288
rect 3936 12248 3942 12260
rect 4157 12257 4169 12260
rect 4203 12257 4215 12291
rect 10888 12288 10916 12384
rect 12176 12356 12204 12384
rect 12728 12356 12756 12396
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 16301 12427 16359 12433
rect 16301 12393 16313 12427
rect 16347 12424 16359 12427
rect 16574 12424 16580 12436
rect 16347 12396 16580 12424
rect 16347 12393 16359 12396
rect 16301 12387 16359 12393
rect 16546 12384 16580 12396
rect 16632 12384 16638 12436
rect 17034 12384 17040 12436
rect 17092 12384 17098 12436
rect 17862 12384 17868 12436
rect 17920 12384 17926 12436
rect 22462 12384 22468 12436
rect 22520 12384 22526 12436
rect 12176 12328 12756 12356
rect 4157 12251 4215 12257
rect 10060 12260 10824 12288
rect 10888 12260 12296 12288
rect 10060 12232 10088 12260
rect 10042 12180 10048 12232
rect 10100 12180 10106 12232
rect 10689 12223 10747 12229
rect 10689 12189 10701 12223
rect 10735 12189 10747 12223
rect 10796 12220 10824 12260
rect 10873 12223 10931 12229
rect 10873 12220 10885 12223
rect 10796 12192 10885 12220
rect 10689 12183 10747 12189
rect 10873 12189 10885 12192
rect 10919 12220 10931 12223
rect 10962 12220 10968 12232
rect 10919 12192 10968 12220
rect 10919 12189 10931 12192
rect 10873 12183 10931 12189
rect 4433 12155 4491 12161
rect 4433 12121 4445 12155
rect 4479 12152 4491 12155
rect 4706 12152 4712 12164
rect 4479 12124 4712 12152
rect 4479 12121 4491 12124
rect 4433 12115 4491 12121
rect 4706 12112 4712 12124
rect 4764 12112 4770 12164
rect 5166 12112 5172 12164
rect 5224 12112 5230 12164
rect 6181 12155 6239 12161
rect 6181 12121 6193 12155
rect 6227 12152 6239 12155
rect 7190 12152 7196 12164
rect 6227 12124 7196 12152
rect 6227 12121 6239 12124
rect 6181 12115 6239 12121
rect 7190 12112 7196 12124
rect 7248 12152 7254 12164
rect 10226 12152 10232 12164
rect 7248 12124 10232 12152
rect 7248 12112 7254 12124
rect 10226 12112 10232 12124
rect 10284 12152 10290 12164
rect 10704 12152 10732 12183
rect 10962 12180 10968 12192
rect 11020 12180 11026 12232
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11425 12223 11483 12229
rect 11425 12220 11437 12223
rect 11388 12192 11437 12220
rect 11388 12180 11394 12192
rect 11425 12189 11437 12192
rect 11471 12189 11483 12223
rect 11425 12183 11483 12189
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 11808 12229 11836 12260
rect 11609 12223 11667 12229
rect 11609 12220 11621 12223
rect 11572 12192 11621 12220
rect 11572 12180 11578 12192
rect 11609 12189 11621 12192
rect 11655 12189 11667 12223
rect 11609 12183 11667 12189
rect 11701 12223 11759 12229
rect 11701 12189 11713 12223
rect 11747 12189 11759 12223
rect 11701 12183 11759 12189
rect 11793 12223 11851 12229
rect 11793 12189 11805 12223
rect 11839 12189 11851 12223
rect 11793 12183 11851 12189
rect 10284 12124 10732 12152
rect 11716 12152 11744 12183
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 12268 12229 12296 12260
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11940 12192 11989 12220
rect 11940 12180 11946 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 12526 12180 12532 12232
rect 12584 12180 12590 12232
rect 12728 12229 12756 12328
rect 13909 12359 13967 12365
rect 13909 12325 13921 12359
rect 13955 12356 13967 12359
rect 16546 12356 16574 12384
rect 16853 12359 16911 12365
rect 16853 12356 16865 12359
rect 13955 12328 14964 12356
rect 16546 12328 16865 12356
rect 13955 12325 13967 12328
rect 13909 12319 13967 12325
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13722 12288 13728 12300
rect 13679 12260 13728 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 14277 12291 14335 12297
rect 14277 12257 14289 12291
rect 14323 12288 14335 12291
rect 14829 12291 14887 12297
rect 14829 12288 14841 12291
rect 14323 12260 14841 12288
rect 14323 12257 14335 12260
rect 14277 12251 14335 12257
rect 14829 12257 14841 12260
rect 14875 12257 14887 12291
rect 14829 12251 14887 12257
rect 12713 12223 12771 12229
rect 12713 12189 12725 12223
rect 12759 12189 12771 12223
rect 12713 12183 12771 12189
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 14182 12220 14188 12232
rect 14139 12192 14188 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 14182 12180 14188 12192
rect 14240 12180 14246 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14936 12229 14964 12328
rect 16853 12325 16865 12328
rect 16899 12325 16911 12359
rect 16853 12319 16911 12325
rect 20625 12359 20683 12365
rect 20625 12325 20637 12359
rect 20671 12356 20683 12359
rect 21634 12356 21640 12368
rect 20671 12328 21640 12356
rect 20671 12325 20683 12328
rect 20625 12319 20683 12325
rect 21634 12316 21640 12328
rect 21692 12316 21698 12368
rect 20165 12291 20223 12297
rect 20165 12288 20177 12291
rect 15028 12260 20177 12288
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14424 12192 14565 12220
rect 14424 12180 14430 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14921 12223 14979 12229
rect 14921 12189 14933 12223
rect 14967 12189 14979 12223
rect 14921 12183 14979 12189
rect 12544 12152 12572 12180
rect 11716 12124 12572 12152
rect 12621 12155 12679 12161
rect 10284 12112 10290 12124
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 15028 12152 15056 12260
rect 20165 12257 20177 12260
rect 20211 12257 20223 12291
rect 20809 12291 20867 12297
rect 20809 12288 20821 12291
rect 20165 12251 20223 12257
rect 20272 12260 20821 12288
rect 15933 12223 15991 12229
rect 15933 12220 15945 12223
rect 12667 12124 15056 12152
rect 15672 12192 15945 12220
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 15672 12096 15700 12192
rect 15933 12189 15945 12192
rect 15979 12220 15991 12223
rect 16577 12223 16635 12229
rect 16577 12220 16589 12223
rect 15979 12192 16589 12220
rect 15979 12189 15991 12192
rect 15933 12183 15991 12189
rect 16577 12189 16589 12192
rect 16623 12189 16635 12223
rect 17126 12220 17132 12232
rect 16577 12183 16635 12189
rect 16868 12192 17132 12220
rect 16868 12164 16896 12192
rect 17126 12180 17132 12192
rect 17184 12220 17190 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 17184 12192 17417 12220
rect 17184 12180 17190 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 17494 12180 17500 12232
rect 17552 12180 17558 12232
rect 20272 12229 20300 12260
rect 20809 12257 20821 12260
rect 20855 12257 20867 12291
rect 20809 12251 20867 12257
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 21729 12291 21787 12297
rect 21729 12288 21741 12291
rect 21315 12260 21741 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 21729 12257 21741 12260
rect 21775 12288 21787 12291
rect 22186 12288 22192 12300
rect 21775 12260 22192 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 17681 12223 17739 12229
rect 17681 12189 17693 12223
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20717 12223 20775 12229
rect 20717 12189 20729 12223
rect 20763 12189 20775 12223
rect 20717 12183 20775 12189
rect 20901 12223 20959 12229
rect 20901 12189 20913 12223
rect 20947 12220 20959 12223
rect 21284 12220 21312 12251
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 20947 12192 21312 12220
rect 22281 12223 22339 12229
rect 20947 12189 20959 12192
rect 20901 12183 20959 12189
rect 22281 12189 22293 12223
rect 22327 12189 22339 12223
rect 22281 12183 22339 12189
rect 24397 12223 24455 12229
rect 24397 12189 24409 12223
rect 24443 12220 24455 12223
rect 24443 12192 24992 12220
rect 24443 12189 24455 12192
rect 24397 12183 24455 12189
rect 16301 12155 16359 12161
rect 16301 12121 16313 12155
rect 16347 12152 16359 12155
rect 16758 12152 16764 12164
rect 16347 12124 16764 12152
rect 16347 12121 16359 12124
rect 16301 12115 16359 12121
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 16850 12112 16856 12164
rect 16908 12112 16914 12164
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17696 12152 17724 12183
rect 17000 12124 17724 12152
rect 17000 12112 17006 12124
rect 20732 12096 20760 12183
rect 22296 12152 22324 12183
rect 22020 12124 22324 12152
rect 22020 12096 22048 12124
rect 24964 12096 24992 12192
rect 33134 12180 33140 12232
rect 33192 12180 33198 12232
rect 34333 12155 34391 12161
rect 34333 12121 34345 12155
rect 34379 12152 34391 12155
rect 34882 12152 34888 12164
rect 34379 12124 34888 12152
rect 34379 12121 34391 12124
rect 34333 12115 34391 12121
rect 34882 12112 34888 12124
rect 34940 12112 34946 12164
rect 11606 12044 11612 12096
rect 11664 12044 11670 12096
rect 12158 12044 12164 12096
rect 12216 12044 12222 12096
rect 12342 12044 12348 12096
rect 12400 12044 12406 12096
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 15654 12044 15660 12096
rect 15712 12044 15718 12096
rect 15749 12087 15807 12093
rect 15749 12053 15761 12087
rect 15795 12084 15807 12087
rect 16114 12084 16120 12096
rect 15795 12056 16120 12084
rect 15795 12053 15807 12056
rect 15749 12047 15807 12053
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 16485 12087 16543 12093
rect 16485 12053 16497 12087
rect 16531 12084 16543 12087
rect 17494 12084 17500 12096
rect 16531 12056 17500 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 20714 12044 20720 12096
rect 20772 12044 20778 12096
rect 21818 12044 21824 12096
rect 21876 12044 21882 12096
rect 22002 12044 22008 12096
rect 22060 12044 22066 12096
rect 24394 12044 24400 12096
rect 24452 12084 24458 12096
rect 24489 12087 24547 12093
rect 24489 12084 24501 12087
rect 24452 12056 24501 12084
rect 24452 12044 24458 12056
rect 24489 12053 24501 12056
rect 24535 12053 24547 12087
rect 24489 12047 24547 12053
rect 24946 12044 24952 12096
rect 25004 12044 25010 12096
rect 1104 11994 35236 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 35236 11994
rect 1104 11920 35236 11942
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 5224 11852 5273 11880
rect 5224 11840 5230 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 5261 11843 5319 11849
rect 5534 11840 5540 11892
rect 5592 11880 5598 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 5592 11852 5641 11880
rect 5592 11840 5598 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 11606 11840 11612 11892
rect 11664 11840 11670 11892
rect 11793 11883 11851 11889
rect 11793 11849 11805 11883
rect 11839 11880 11851 11883
rect 11882 11880 11888 11892
rect 11839 11852 11888 11880
rect 11839 11849 11851 11852
rect 11793 11843 11851 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12158 11840 12164 11892
rect 12216 11840 12222 11892
rect 12434 11840 12440 11892
rect 12492 11840 12498 11892
rect 15654 11840 15660 11892
rect 15712 11840 15718 11892
rect 15746 11840 15752 11892
rect 15804 11840 15810 11892
rect 16114 11840 16120 11892
rect 16172 11840 16178 11892
rect 16301 11883 16359 11889
rect 16301 11849 16313 11883
rect 16347 11880 16359 11883
rect 16758 11880 16764 11892
rect 16347 11852 16764 11880
rect 16347 11849 16359 11852
rect 16301 11843 16359 11849
rect 16758 11840 16764 11852
rect 16816 11840 16822 11892
rect 33134 11880 33140 11892
rect 26206 11852 33140 11880
rect 5169 11747 5227 11753
rect 5169 11713 5181 11747
rect 5215 11744 5227 11747
rect 5552 11744 5580 11840
rect 5215 11716 5580 11744
rect 11624 11744 11652 11840
rect 12176 11753 12204 11840
rect 12452 11812 12480 11840
rect 12452 11784 12664 11812
rect 12636 11753 12664 11784
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 15289 11815 15347 11821
rect 15289 11812 15301 11815
rect 14240 11784 15301 11812
rect 14240 11772 14246 11784
rect 15289 11781 15301 11784
rect 15335 11781 15347 11815
rect 15489 11815 15547 11821
rect 15489 11812 15501 11815
rect 15289 11775 15347 11781
rect 15396 11784 15501 11812
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11624 11716 11989 11744
rect 5215 11713 5227 11716
rect 5169 11707 5227 11713
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12161 11747 12219 11753
rect 12161 11713 12173 11747
rect 12207 11713 12219 11747
rect 12161 11707 12219 11713
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11713 12495 11747
rect 12437 11707 12495 11713
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 14366 11744 14372 11756
rect 12667 11716 14372 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 11882 11636 11888 11688
rect 11940 11636 11946 11688
rect 11992 11676 12020 11707
rect 12452 11676 12480 11707
rect 14366 11704 14372 11716
rect 14424 11744 14430 11756
rect 15396 11744 15424 11784
rect 15489 11781 15501 11784
rect 15535 11781 15547 11815
rect 15489 11775 15547 11781
rect 14424 11716 15424 11744
rect 15764 11744 15792 11840
rect 16132 11812 16160 11840
rect 16850 11812 16856 11824
rect 16132 11784 16856 11812
rect 16850 11772 16856 11784
rect 16908 11772 16914 11824
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 23661 11815 23719 11821
rect 23661 11812 23673 11815
rect 23624 11784 23673 11812
rect 23624 11772 23630 11784
rect 23661 11781 23673 11784
rect 23707 11781 23719 11815
rect 23661 11775 23719 11781
rect 24394 11772 24400 11824
rect 24452 11772 24458 11824
rect 16117 11747 16175 11753
rect 16117 11744 16129 11747
rect 15764 11716 16129 11744
rect 14424 11704 14430 11716
rect 16117 11713 16129 11716
rect 16163 11713 16175 11747
rect 16117 11707 16175 11713
rect 16298 11704 16304 11756
rect 16356 11704 16362 11756
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 17313 11747 17371 11753
rect 17313 11744 17325 11747
rect 16724 11716 17325 11744
rect 16724 11704 16730 11716
rect 17313 11713 17325 11716
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 22097 11747 22155 11753
rect 22097 11713 22109 11747
rect 22143 11713 22155 11747
rect 22097 11707 22155 11713
rect 11992 11648 12480 11676
rect 17405 11679 17463 11685
rect 17405 11645 17417 11679
rect 17451 11676 17463 11679
rect 22002 11676 22008 11688
rect 17451 11648 22008 11676
rect 17451 11645 17463 11648
rect 17405 11639 17463 11645
rect 22002 11636 22008 11648
rect 22060 11636 22066 11688
rect 12345 11611 12403 11617
rect 12345 11577 12357 11611
rect 12391 11608 12403 11611
rect 21818 11608 21824 11620
rect 12391 11580 21824 11608
rect 12391 11577 12403 11580
rect 12345 11571 12403 11577
rect 21818 11568 21824 11580
rect 21876 11608 21882 11620
rect 22112 11608 22140 11707
rect 23290 11636 23296 11688
rect 23348 11676 23354 11688
rect 23385 11679 23443 11685
rect 23385 11676 23397 11679
rect 23348 11648 23397 11676
rect 23348 11636 23354 11648
rect 23385 11645 23397 11648
rect 23431 11645 23443 11679
rect 23385 11639 23443 11645
rect 21876 11580 22140 11608
rect 22465 11611 22523 11617
rect 21876 11568 21882 11580
rect 22465 11577 22477 11611
rect 22511 11608 22523 11611
rect 22511 11580 23520 11608
rect 22511 11577 22523 11580
rect 22465 11571 22523 11577
rect 23492 11552 23520 11580
rect 12618 11500 12624 11552
rect 12676 11500 12682 11552
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 15473 11543 15531 11549
rect 15473 11540 15485 11543
rect 14516 11512 15485 11540
rect 14516 11500 14522 11512
rect 15473 11509 15485 11512
rect 15519 11509 15531 11543
rect 15473 11503 15531 11509
rect 20625 11543 20683 11549
rect 20625 11509 20637 11543
rect 20671 11540 20683 11543
rect 20714 11540 20720 11552
rect 20671 11512 20720 11540
rect 20671 11509 20683 11512
rect 20625 11503 20683 11509
rect 20714 11500 20720 11512
rect 20772 11500 20778 11552
rect 23290 11500 23296 11552
rect 23348 11500 23354 11552
rect 23474 11500 23480 11552
rect 23532 11500 23538 11552
rect 25133 11543 25191 11549
rect 25133 11509 25145 11543
rect 25179 11540 25191 11543
rect 26206 11540 26234 11852
rect 33134 11840 33140 11852
rect 33192 11840 33198 11892
rect 25179 11512 26234 11540
rect 25179 11509 25191 11512
rect 25133 11503 25191 11509
rect 1104 11450 35248 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 35248 11450
rect 1104 11376 35248 11398
rect 6178 11296 6184 11348
rect 6236 11336 6242 11348
rect 6549 11339 6607 11345
rect 6549 11336 6561 11339
rect 6236 11308 6561 11336
rect 6236 11296 6242 11308
rect 6549 11305 6561 11308
rect 6595 11305 6607 11339
rect 6549 11299 6607 11305
rect 12158 11296 12164 11348
rect 12216 11296 12222 11348
rect 12618 11296 12624 11348
rect 12676 11296 12682 11348
rect 1581 11271 1639 11277
rect 1581 11237 1593 11271
rect 1627 11237 1639 11271
rect 1581 11231 1639 11237
rect 1596 11200 1624 11231
rect 4525 11203 4583 11209
rect 4525 11200 4537 11203
rect 1596 11172 4537 11200
rect 4525 11169 4537 11172
rect 4571 11169 4583 11203
rect 4525 11163 4583 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 7282 11200 7288 11212
rect 6319 11172 7288 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 7282 11160 7288 11172
rect 7340 11160 7346 11212
rect 1394 11092 1400 11144
rect 1452 11092 1458 11144
rect 3878 11092 3884 11144
rect 3936 11132 3942 11144
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 3936 11104 4261 11132
rect 3936 11092 3942 11104
rect 4249 11101 4261 11104
rect 4295 11101 4307 11135
rect 12176 11132 12204 11296
rect 12345 11203 12403 11209
rect 12345 11169 12357 11203
rect 12391 11200 12403 11203
rect 12636 11200 12664 11296
rect 12391 11172 12664 11200
rect 12391 11169 12403 11172
rect 12345 11163 12403 11169
rect 12253 11135 12311 11141
rect 12253 11132 12265 11135
rect 12176 11104 12265 11132
rect 4249 11095 4307 11101
rect 12253 11101 12265 11104
rect 12299 11101 12311 11135
rect 24489 11135 24547 11141
rect 24489 11132 24501 11135
rect 12253 11095 12311 11101
rect 23492 11104 24501 11132
rect 5534 11024 5540 11076
rect 5592 11024 5598 11076
rect 12342 11024 12348 11076
rect 12400 11064 12406 11076
rect 20714 11064 20720 11076
rect 12400 11036 20720 11064
rect 12400 11024 12406 11036
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 23382 10956 23388 11008
rect 23440 10996 23446 11008
rect 23492 10996 23520 11104
rect 24489 11101 24501 11104
rect 24535 11132 24547 11135
rect 24946 11132 24952 11144
rect 24535 11104 24952 11132
rect 24535 11101 24547 11104
rect 24489 11095 24547 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 24581 11067 24639 11073
rect 24581 11033 24593 11067
rect 24627 11064 24639 11067
rect 24854 11064 24860 11076
rect 24627 11036 24860 11064
rect 24627 11033 24639 11036
rect 24581 11027 24639 11033
rect 24854 11024 24860 11036
rect 24912 11024 24918 11076
rect 23440 10968 23520 10996
rect 23440 10956 23446 10968
rect 1104 10906 35236 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 35236 10906
rect 1104 10832 35236 10854
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5534 10792 5540 10804
rect 5307 10764 5540 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5534 10752 5540 10764
rect 5592 10752 5598 10804
rect 5626 10752 5632 10804
rect 5684 10752 5690 10804
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10656 5227 10659
rect 5644 10656 5672 10752
rect 12618 10684 12624 10736
rect 12676 10724 12682 10736
rect 13725 10727 13783 10733
rect 13725 10724 13737 10727
rect 12676 10696 13737 10724
rect 12676 10684 12682 10696
rect 13725 10693 13737 10696
rect 13771 10693 13783 10727
rect 13725 10687 13783 10693
rect 14458 10684 14464 10736
rect 14516 10684 14522 10736
rect 23474 10684 23480 10736
rect 23532 10724 23538 10736
rect 23753 10727 23811 10733
rect 23753 10724 23765 10727
rect 23532 10696 23765 10724
rect 23532 10684 23538 10696
rect 23753 10693 23765 10696
rect 23799 10693 23811 10727
rect 23753 10687 23811 10693
rect 5215 10628 5672 10656
rect 5215 10625 5227 10628
rect 5169 10619 5227 10625
rect 24854 10616 24860 10668
rect 24912 10616 24918 10668
rect 13449 10591 13507 10597
rect 13449 10588 13461 10591
rect 13280 10560 13461 10588
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 13280 10461 13308 10560
rect 13449 10557 13461 10560
rect 13495 10557 13507 10591
rect 13449 10551 13507 10557
rect 23290 10548 23296 10600
rect 23348 10588 23354 10600
rect 23477 10591 23535 10597
rect 23477 10588 23489 10591
rect 23348 10560 23489 10588
rect 23348 10548 23354 10560
rect 23477 10557 23489 10560
rect 23523 10557 23535 10591
rect 23477 10551 23535 10557
rect 13265 10455 13323 10461
rect 13265 10452 13277 10455
rect 10008 10424 13277 10452
rect 10008 10412 10014 10424
rect 13265 10421 13277 10424
rect 13311 10421 13323 10455
rect 13265 10415 13323 10421
rect 15194 10412 15200 10464
rect 15252 10412 15258 10464
rect 21358 10412 21364 10464
rect 21416 10452 21422 10464
rect 23308 10461 23336 10548
rect 25225 10523 25283 10529
rect 25225 10489 25237 10523
rect 25271 10520 25283 10523
rect 25271 10492 26234 10520
rect 25271 10489 25283 10492
rect 25225 10483 25283 10489
rect 23293 10455 23351 10461
rect 23293 10452 23305 10455
rect 21416 10424 23305 10452
rect 21416 10412 21422 10424
rect 23293 10421 23305 10424
rect 23339 10421 23351 10455
rect 26206 10452 26234 10492
rect 33134 10452 33140 10464
rect 26206 10424 33140 10452
rect 23293 10415 23351 10421
rect 33134 10412 33140 10424
rect 33192 10412 33198 10464
rect 1104 10362 35248 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 35248 10362
rect 1104 10288 35248 10310
rect 5626 10208 5632 10260
rect 5684 10248 5690 10260
rect 5684 10220 6914 10248
rect 5684 10208 5690 10220
rect 6886 10044 6914 10220
rect 14458 10208 14464 10260
rect 14516 10208 14522 10260
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 32950 10248 32956 10260
rect 15252 10220 32956 10248
rect 15252 10208 15258 10220
rect 32950 10208 32956 10220
rect 33008 10208 33014 10260
rect 14369 10047 14427 10053
rect 14369 10044 14381 10047
rect 6886 10016 14381 10044
rect 14369 10013 14381 10016
rect 14415 10044 14427 10047
rect 14829 10047 14887 10053
rect 14829 10044 14841 10047
rect 14415 10016 14841 10044
rect 14415 10013 14427 10016
rect 14369 10007 14427 10013
rect 14829 10013 14841 10016
rect 14875 10044 14887 10047
rect 23382 10044 23388 10056
rect 14875 10016 23388 10044
rect 14875 10013 14887 10016
rect 14829 10007 14887 10013
rect 23382 10004 23388 10016
rect 23440 10004 23446 10056
rect 33134 10004 33140 10056
rect 33192 10004 33198 10056
rect 34330 9936 34336 9988
rect 34388 9936 34394 9988
rect 1104 9818 35236 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 35236 9818
rect 1104 9744 35236 9766
rect 1104 9274 35248 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 35248 9274
rect 1104 9200 35248 9222
rect 1581 9163 1639 9169
rect 1581 9129 1593 9163
rect 1627 9160 1639 9163
rect 4798 9160 4804 9172
rect 1627 9132 4804 9160
rect 1627 9129 1639 9132
rect 1581 9123 1639 9129
rect 4798 9120 4804 9132
rect 4856 9120 4862 9172
rect 6178 9120 6184 9172
rect 6236 9160 6242 9172
rect 6273 9163 6331 9169
rect 6273 9160 6285 9163
rect 6236 9132 6285 9160
rect 6236 9120 6242 9132
rect 6273 9129 6285 9132
rect 6319 9129 6331 9163
rect 6273 9123 6331 9129
rect 3973 9027 4031 9033
rect 3973 8993 3985 9027
rect 4019 9024 4031 9027
rect 6196 9024 6224 9120
rect 4019 8996 6224 9024
rect 4019 8993 4031 8996
rect 3973 8987 4031 8993
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 4249 8891 4307 8897
rect 4249 8857 4261 8891
rect 4295 8888 4307 8891
rect 4522 8888 4528 8900
rect 4295 8860 4528 8888
rect 4295 8857 4307 8860
rect 4249 8851 4307 8857
rect 4522 8848 4528 8860
rect 4580 8848 4586 8900
rect 4982 8848 4988 8900
rect 5040 8848 5046 8900
rect 5920 8820 5948 8996
rect 5997 8891 6055 8897
rect 5997 8857 6009 8891
rect 6043 8888 6055 8891
rect 10042 8888 10048 8900
rect 6043 8860 10048 8888
rect 6043 8857 6055 8860
rect 5997 8851 6055 8857
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 9950 8820 9956 8832
rect 5920 8792 9956 8820
rect 9950 8780 9956 8792
rect 10008 8780 10014 8832
rect 1104 8730 35236 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 35236 8730
rect 1104 8656 35236 8678
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 5040 8588 5089 8616
rect 5040 8576 5046 8588
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 5537 8619 5595 8625
rect 5537 8585 5549 8619
rect 5583 8616 5595 8619
rect 5626 8616 5632 8628
rect 5583 8588 5632 8616
rect 5583 8585 5595 8588
rect 5537 8579 5595 8585
rect 4985 8483 5043 8489
rect 4985 8449 4997 8483
rect 5031 8480 5043 8483
rect 5552 8480 5580 8579
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5031 8452 5580 8480
rect 5031 8449 5043 8452
rect 4985 8443 5043 8449
rect 1104 8186 35248 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 35248 8186
rect 1104 8112 35248 8134
rect 32950 8032 32956 8084
rect 33008 8032 33014 8084
rect 32968 7868 32996 8032
rect 33137 7871 33195 7877
rect 33137 7868 33149 7871
rect 32968 7840 33149 7868
rect 33137 7837 33149 7840
rect 33183 7837 33195 7871
rect 33137 7831 33195 7837
rect 34333 7803 34391 7809
rect 34333 7769 34345 7803
rect 34379 7800 34391 7803
rect 34882 7800 34888 7812
rect 34379 7772 34888 7800
rect 34379 7769 34391 7772
rect 34333 7763 34391 7769
rect 34882 7760 34888 7772
rect 34940 7760 34946 7812
rect 1104 7642 35236 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 35236 7642
rect 1104 7568 35236 7590
rect 1104 7098 35248 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 35248 7098
rect 1104 7024 35248 7046
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 992 6752 1409 6780
rect 992 6740 998 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 1397 6743 1455 6749
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 4890 6644 4896 6656
rect 1627 6616 4896 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 4890 6604 4896 6616
rect 4948 6604 4954 6656
rect 1104 6554 35236 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 35236 6554
rect 1104 6480 35236 6502
rect 1104 6010 35248 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 35248 6010
rect 1104 5936 35248 5958
rect 21634 5720 21640 5772
rect 21692 5720 21698 5772
rect 21358 5692 21364 5704
rect 21192 5664 21364 5692
rect 20806 5516 20812 5568
rect 20864 5556 20870 5568
rect 21192 5565 21220 5664
rect 21358 5652 21364 5664
rect 21416 5652 21422 5704
rect 23198 5652 23204 5704
rect 23256 5692 23262 5704
rect 23385 5695 23443 5701
rect 23385 5692 23397 5695
rect 23256 5664 23397 5692
rect 23256 5652 23262 5664
rect 23385 5661 23397 5664
rect 23431 5692 23443 5695
rect 23661 5695 23719 5701
rect 23661 5692 23673 5695
rect 23431 5664 23673 5692
rect 23431 5661 23443 5664
rect 23385 5655 23443 5661
rect 23661 5661 23673 5664
rect 23707 5661 23719 5695
rect 33137 5695 33195 5701
rect 33137 5692 33149 5695
rect 23661 5655 23719 5661
rect 26206 5664 33149 5692
rect 23293 5627 23351 5633
rect 23293 5624 23305 5627
rect 22862 5596 23305 5624
rect 23293 5593 23305 5596
rect 23339 5593 23351 5627
rect 26206 5624 26234 5664
rect 33137 5661 33149 5664
rect 33183 5661 33195 5695
rect 33137 5655 33195 5661
rect 23293 5587 23351 5593
rect 23584 5596 26234 5624
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 20864 5528 21189 5556
rect 20864 5516 20870 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 21177 5519 21235 5525
rect 23109 5559 23167 5565
rect 23109 5525 23121 5559
rect 23155 5556 23167 5559
rect 23584 5556 23612 5596
rect 34330 5584 34336 5636
rect 34388 5584 34394 5636
rect 23155 5528 23612 5556
rect 23155 5525 23167 5528
rect 23109 5519 23167 5525
rect 1104 5466 35236 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 35236 5466
rect 1104 5392 35236 5414
rect 1104 4922 35248 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 35248 4922
rect 1104 4848 35248 4870
rect 1581 4811 1639 4817
rect 1581 4777 1593 4811
rect 1627 4808 1639 4811
rect 4614 4808 4620 4820
rect 1627 4780 4620 4808
rect 1627 4777 1639 4780
rect 1581 4771 1639 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 934 4564 940 4616
rect 992 4604 998 4616
rect 1397 4607 1455 4613
rect 1397 4604 1409 4607
rect 992 4576 1409 4604
rect 992 4564 998 4576
rect 1397 4573 1409 4576
rect 1443 4573 1455 4607
rect 1397 4567 1455 4573
rect 1104 4378 35236 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 35236 4378
rect 1104 4304 35236 4326
rect 1104 3834 35248 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 35248 3834
rect 1104 3760 35248 3782
rect 20714 3680 20720 3732
rect 20772 3680 20778 3732
rect 20732 3584 20760 3680
rect 21085 3587 21143 3593
rect 21085 3584 21097 3587
rect 20732 3556 21097 3584
rect 21085 3553 21097 3556
rect 21131 3553 21143 3587
rect 21085 3547 21143 3553
rect 20806 3516 20812 3528
rect 20456 3488 20812 3516
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 20456 3389 20484 3488
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 23198 3516 23204 3528
rect 22879 3488 23204 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 33137 3519 33195 3525
rect 33137 3516 33149 3519
rect 26206 3488 33149 3516
rect 22741 3451 22799 3457
rect 22741 3448 22753 3451
rect 22310 3420 22753 3448
rect 22741 3417 22753 3420
rect 22787 3417 22799 3451
rect 26206 3448 26234 3488
rect 33137 3485 33149 3488
rect 33183 3485 33195 3519
rect 33137 3479 33195 3485
rect 22741 3411 22799 3417
rect 23032 3420 26234 3448
rect 34333 3451 34391 3457
rect 20441 3383 20499 3389
rect 20441 3380 20453 3383
rect 10008 3352 20453 3380
rect 10008 3340 10014 3352
rect 20441 3349 20453 3352
rect 20487 3349 20499 3383
rect 20441 3343 20499 3349
rect 22557 3383 22615 3389
rect 22557 3349 22569 3383
rect 22603 3380 22615 3383
rect 23032 3380 23060 3420
rect 34333 3417 34345 3451
rect 34379 3448 34391 3451
rect 34882 3448 34888 3460
rect 34379 3420 34888 3448
rect 34379 3417 34391 3420
rect 34333 3411 34391 3417
rect 34882 3408 34888 3420
rect 34940 3408 34946 3460
rect 22603 3352 23060 3380
rect 22603 3349 22615 3352
rect 22557 3343 22615 3349
rect 23198 3340 23204 3392
rect 23256 3340 23262 3392
rect 1104 3290 35236 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 35236 3290
rect 1104 3216 35236 3238
rect 20714 3136 20720 3188
rect 20772 3136 20778 3188
rect 1104 2746 35248 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 35248 2746
rect 1104 2672 35248 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 4706 2632 4712 2644
rect 1627 2604 4712 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 9950 2456 9956 2508
rect 10008 2456 10014 2508
rect 23198 2456 23204 2508
rect 23256 2496 23262 2508
rect 27801 2499 27859 2505
rect 27801 2496 27813 2499
rect 23256 2468 27813 2496
rect 23256 2456 23262 2468
rect 27801 2465 27813 2468
rect 27847 2465 27859 2499
rect 27801 2459 27859 2465
rect 934 2388 940 2440
rect 992 2428 998 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 992 2400 1409 2428
rect 992 2388 998 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 27338 2388 27344 2440
rect 27396 2388 27402 2440
rect 1104 2202 35236 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 35236 2202
rect 1104 2128 35236 2150
<< via1 >>
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 940 36116 992 36168
rect 25596 36116 25648 36168
rect 34336 36091 34388 36100
rect 34336 36057 34345 36091
rect 34345 36057 34379 36091
rect 34379 36057 34388 36091
rect 34336 36048 34388 36057
rect 4620 35980 4672 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 940 35028 992 35080
rect 3884 34892 3936 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 23664 33940 23716 33992
rect 34888 33872 34940 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 940 32852 992 32904
rect 4712 32716 4764 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 33140 31807 33192 31816
rect 33140 31773 33149 31807
rect 33149 31773 33183 31807
rect 33183 31773 33192 31807
rect 33140 31764 33192 31773
rect 34336 31739 34388 31748
rect 34336 31705 34345 31739
rect 34345 31705 34379 31739
rect 34379 31705 34388 31739
rect 34336 31696 34388 31705
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1400 30719 1452 30728
rect 1400 30685 1409 30719
rect 1409 30685 1443 30719
rect 1443 30685 1452 30719
rect 1400 30676 1452 30685
rect 4804 30540 4856 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 33324 29588 33376 29640
rect 34888 29520 34940 29572
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 940 28500 992 28552
rect 1584 28407 1636 28416
rect 1584 28373 1593 28407
rect 1593 28373 1627 28407
rect 1627 28373 1636 28407
rect 1584 28364 1636 28373
rect 23572 28364 23624 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 23572 28160 23624 28212
rect 23664 28203 23716 28212
rect 23664 28169 23673 28203
rect 23673 28169 23707 28203
rect 23707 28169 23716 28203
rect 23664 28160 23716 28169
rect 25596 28203 25648 28212
rect 25596 28169 25605 28203
rect 25605 28169 25639 28203
rect 25639 28169 25648 28203
rect 25596 28160 25648 28169
rect 6000 28024 6052 28076
rect 22928 28092 22980 28144
rect 24860 28092 24912 28144
rect 23848 28067 23900 28076
rect 23848 28033 23857 28067
rect 23857 28033 23891 28067
rect 23891 28033 23900 28067
rect 23848 28024 23900 28033
rect 22192 27999 22244 28008
rect 22192 27965 22201 27999
rect 22201 27965 22235 27999
rect 22235 27965 22244 27999
rect 22192 27956 22244 27965
rect 5908 27820 5960 27872
rect 22652 27820 22704 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 1584 27616 1636 27668
rect 11980 27548 12032 27600
rect 12440 27523 12492 27532
rect 12440 27489 12449 27523
rect 12449 27489 12483 27523
rect 12483 27489 12492 27523
rect 12440 27480 12492 27489
rect 22192 27616 22244 27668
rect 22652 27659 22704 27668
rect 22652 27625 22661 27659
rect 22661 27625 22695 27659
rect 22695 27625 22704 27659
rect 22652 27616 22704 27625
rect 22928 27616 22980 27668
rect 23848 27659 23900 27668
rect 23848 27625 23857 27659
rect 23857 27625 23891 27659
rect 23891 27625 23900 27659
rect 23848 27616 23900 27625
rect 4068 27412 4120 27464
rect 4712 27319 4764 27328
rect 4712 27285 4721 27319
rect 4721 27285 4755 27319
rect 4755 27285 4764 27319
rect 4712 27276 4764 27285
rect 12532 27455 12584 27464
rect 12532 27421 12541 27455
rect 12541 27421 12575 27455
rect 12575 27421 12584 27455
rect 12532 27412 12584 27421
rect 12992 27455 13044 27464
rect 12992 27421 13001 27455
rect 13001 27421 13035 27455
rect 13035 27421 13044 27455
rect 12992 27412 13044 27421
rect 14924 27480 14976 27532
rect 18972 27480 19024 27532
rect 5908 27344 5960 27396
rect 7012 27344 7064 27396
rect 6000 27276 6052 27328
rect 6552 27276 6604 27328
rect 11888 27276 11940 27328
rect 13084 27276 13136 27328
rect 14464 27344 14516 27396
rect 14832 27455 14884 27464
rect 14832 27421 14841 27455
rect 14841 27421 14875 27455
rect 14875 27421 14884 27455
rect 14832 27412 14884 27421
rect 18144 27412 18196 27464
rect 19248 27412 19300 27464
rect 22376 27548 22428 27600
rect 24124 27480 24176 27532
rect 21824 27455 21876 27464
rect 21824 27421 21833 27455
rect 21833 27421 21867 27455
rect 21867 27421 21876 27455
rect 21824 27412 21876 27421
rect 22192 27455 22244 27464
rect 22192 27421 22201 27455
rect 22201 27421 22235 27455
rect 22235 27421 22244 27455
rect 22192 27412 22244 27421
rect 22376 27455 22428 27464
rect 22376 27421 22385 27455
rect 22385 27421 22419 27455
rect 22419 27421 22428 27455
rect 22376 27412 22428 27421
rect 22008 27344 22060 27396
rect 33232 27455 33284 27464
rect 33232 27421 33241 27455
rect 33241 27421 33275 27455
rect 33275 27421 33284 27455
rect 33232 27412 33284 27421
rect 24676 27387 24728 27396
rect 24676 27353 24685 27387
rect 24685 27353 24719 27387
rect 24719 27353 24728 27387
rect 24676 27344 24728 27353
rect 25412 27344 25464 27396
rect 34888 27344 34940 27396
rect 14556 27276 14608 27328
rect 17132 27276 17184 27328
rect 17684 27276 17736 27328
rect 18512 27276 18564 27328
rect 19156 27276 19208 27328
rect 22192 27276 22244 27328
rect 22284 27276 22336 27328
rect 24032 27276 24084 27328
rect 24860 27276 24912 27328
rect 33140 27276 33192 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 12532 27072 12584 27124
rect 4068 27004 4120 27056
rect 4712 27004 4764 27056
rect 12992 27072 13044 27124
rect 14464 27072 14516 27124
rect 14832 27072 14884 27124
rect 11888 26979 11940 26988
rect 11888 26945 11897 26979
rect 11897 26945 11931 26979
rect 11931 26945 11940 26979
rect 11888 26936 11940 26945
rect 4804 26868 4856 26920
rect 5908 26911 5960 26920
rect 5908 26877 5917 26911
rect 5917 26877 5951 26911
rect 5951 26877 5960 26911
rect 5908 26868 5960 26877
rect 11980 26868 12032 26920
rect 12992 26979 13044 26988
rect 12992 26945 13001 26979
rect 13001 26945 13035 26979
rect 13035 26945 13044 26979
rect 12992 26936 13044 26945
rect 6552 26775 6604 26784
rect 6552 26741 6561 26775
rect 6561 26741 6595 26775
rect 6595 26741 6604 26775
rect 6552 26732 6604 26741
rect 13176 26979 13228 26988
rect 13176 26945 13185 26979
rect 13185 26945 13219 26979
rect 13219 26945 13228 26979
rect 13176 26936 13228 26945
rect 14188 26936 14240 26988
rect 16028 27004 16080 27056
rect 16764 27004 16816 27056
rect 14924 26936 14976 26988
rect 14556 26868 14608 26920
rect 15568 26979 15620 26988
rect 15568 26945 15577 26979
rect 15577 26945 15611 26979
rect 15611 26945 15620 26979
rect 15568 26936 15620 26945
rect 15936 26979 15988 26988
rect 15936 26945 15945 26979
rect 15945 26945 15979 26979
rect 15979 26945 15988 26979
rect 15936 26936 15988 26945
rect 17776 27072 17828 27124
rect 17592 27004 17644 27056
rect 19156 27115 19208 27124
rect 19156 27081 19165 27115
rect 19165 27081 19199 27115
rect 19199 27081 19208 27115
rect 19156 27072 19208 27081
rect 19248 27115 19300 27124
rect 19248 27081 19257 27115
rect 19257 27081 19291 27115
rect 19291 27081 19300 27115
rect 19248 27072 19300 27081
rect 20168 27072 20220 27124
rect 18512 26936 18564 26988
rect 18696 26979 18748 26988
rect 18696 26945 18705 26979
rect 18705 26945 18739 26979
rect 18739 26945 18748 26979
rect 18696 26936 18748 26945
rect 18972 26979 19024 26988
rect 18972 26945 18981 26979
rect 18981 26945 19015 26979
rect 19015 26945 19024 26979
rect 18972 26936 19024 26945
rect 15844 26911 15896 26920
rect 15844 26877 15853 26911
rect 15853 26877 15887 26911
rect 15887 26877 15896 26911
rect 15844 26868 15896 26877
rect 17684 26868 17736 26920
rect 12992 26732 13044 26784
rect 16120 26800 16172 26852
rect 16764 26732 16816 26784
rect 17040 26843 17092 26852
rect 17040 26809 17049 26843
rect 17049 26809 17083 26843
rect 17083 26809 17092 26843
rect 17040 26800 17092 26809
rect 18052 26843 18104 26852
rect 18052 26809 18061 26843
rect 18061 26809 18095 26843
rect 18095 26809 18104 26843
rect 18052 26800 18104 26809
rect 18144 26800 18196 26852
rect 19248 26732 19300 26784
rect 19984 26800 20036 26852
rect 25412 27072 25464 27124
rect 22008 26979 22060 26988
rect 22008 26945 22017 26979
rect 22017 26945 22051 26979
rect 22051 26945 22060 26979
rect 22008 26936 22060 26945
rect 22192 26936 22244 26988
rect 24032 26936 24084 26988
rect 21824 26868 21876 26920
rect 22284 26868 22336 26920
rect 24676 26868 24728 26920
rect 22100 26732 22152 26784
rect 22376 26732 22428 26784
rect 25228 26775 25280 26784
rect 25228 26741 25237 26775
rect 25237 26741 25271 26775
rect 25271 26741 25280 26775
rect 25228 26732 25280 26741
rect 25964 26775 26016 26784
rect 25964 26741 25973 26775
rect 25973 26741 26007 26775
rect 26007 26741 26016 26775
rect 25964 26732 26016 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6000 26571 6052 26580
rect 6000 26537 6009 26571
rect 6009 26537 6043 26571
rect 6043 26537 6052 26571
rect 6000 26528 6052 26537
rect 12440 26528 12492 26580
rect 13176 26528 13228 26580
rect 14188 26571 14240 26580
rect 14188 26537 14197 26571
rect 14197 26537 14231 26571
rect 14231 26537 14240 26571
rect 14188 26528 14240 26537
rect 18696 26528 18748 26580
rect 24124 26571 24176 26580
rect 24124 26537 24133 26571
rect 24133 26537 24167 26571
rect 24167 26537 24176 26571
rect 24124 26528 24176 26537
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 5448 26324 5500 26376
rect 11704 26367 11756 26376
rect 11704 26333 11713 26367
rect 11713 26333 11747 26367
rect 11747 26333 11756 26367
rect 11704 26324 11756 26333
rect 4620 26256 4672 26308
rect 5540 26256 5592 26308
rect 12256 26324 12308 26376
rect 15108 26460 15160 26512
rect 15568 26460 15620 26512
rect 14188 26367 14240 26376
rect 14188 26333 14197 26367
rect 14197 26333 14231 26367
rect 14231 26333 14240 26367
rect 14188 26324 14240 26333
rect 12808 26256 12860 26308
rect 15200 26256 15252 26308
rect 5632 26231 5684 26240
rect 5632 26197 5641 26231
rect 5641 26197 5675 26231
rect 5675 26197 5684 26231
rect 5632 26188 5684 26197
rect 11796 26188 11848 26240
rect 15384 26188 15436 26240
rect 16028 26367 16080 26376
rect 16028 26333 16037 26367
rect 16037 26333 16071 26367
rect 16071 26333 16080 26367
rect 16028 26324 16080 26333
rect 17040 26460 17092 26512
rect 17132 26460 17184 26512
rect 18052 26460 18104 26512
rect 23020 26460 23072 26512
rect 33324 26392 33376 26444
rect 22836 26324 22888 26376
rect 23112 26324 23164 26376
rect 16120 26256 16172 26308
rect 16764 26256 16816 26308
rect 17592 26256 17644 26308
rect 17776 26256 17828 26308
rect 19248 26256 19300 26308
rect 23480 26256 23532 26308
rect 24676 26299 24728 26308
rect 24676 26265 24685 26299
rect 24685 26265 24719 26299
rect 24719 26265 24728 26299
rect 24676 26256 24728 26265
rect 25228 26256 25280 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 4528 25959 4580 25968
rect 4528 25925 4537 25959
rect 4537 25925 4571 25959
rect 4571 25925 4580 25959
rect 4528 25916 4580 25925
rect 5540 25916 5592 25968
rect 10692 25891 10744 25900
rect 10692 25857 10701 25891
rect 10701 25857 10735 25891
rect 10735 25857 10744 25891
rect 10692 25848 10744 25857
rect 10784 25891 10836 25900
rect 10784 25857 10793 25891
rect 10793 25857 10827 25891
rect 10827 25857 10836 25891
rect 10784 25848 10836 25857
rect 11704 25916 11756 25968
rect 14188 25984 14240 26036
rect 15936 25984 15988 26036
rect 17776 25984 17828 26036
rect 22192 26027 22244 26036
rect 22192 25993 22201 26027
rect 22201 25993 22235 26027
rect 22235 25993 22244 26027
rect 22192 25984 22244 25993
rect 23480 25984 23532 26036
rect 24676 25984 24728 26036
rect 11796 25891 11848 25900
rect 11796 25857 11805 25891
rect 11805 25857 11839 25891
rect 11839 25857 11848 25891
rect 11796 25848 11848 25857
rect 12808 25848 12860 25900
rect 15200 25916 15252 25968
rect 4068 25780 4120 25832
rect 12256 25780 12308 25832
rect 6920 25712 6972 25764
rect 15108 25848 15160 25900
rect 15568 25891 15620 25900
rect 15568 25857 15577 25891
rect 15577 25857 15611 25891
rect 15611 25857 15620 25891
rect 15568 25848 15620 25857
rect 15660 25891 15712 25900
rect 15660 25857 15669 25891
rect 15669 25857 15703 25891
rect 15703 25857 15712 25891
rect 15660 25848 15712 25857
rect 16396 25848 16448 25900
rect 22100 25916 22152 25968
rect 18420 25848 18472 25900
rect 19984 25848 20036 25900
rect 6092 25644 6144 25696
rect 6552 25687 6604 25696
rect 6552 25653 6561 25687
rect 6561 25653 6595 25687
rect 6595 25653 6604 25687
rect 6552 25644 6604 25653
rect 6644 25644 6696 25696
rect 10140 25644 10192 25696
rect 11704 25644 11756 25696
rect 12164 25644 12216 25696
rect 13820 25712 13872 25764
rect 16028 25780 16080 25832
rect 17132 25780 17184 25832
rect 20996 25823 21048 25832
rect 20996 25789 21005 25823
rect 21005 25789 21039 25823
rect 21039 25789 21048 25823
rect 20996 25780 21048 25789
rect 15384 25644 15436 25696
rect 18236 25644 18288 25696
rect 20444 25644 20496 25696
rect 22100 25687 22152 25696
rect 22100 25653 22109 25687
rect 22109 25653 22143 25687
rect 22143 25653 22152 25687
rect 22100 25644 22152 25653
rect 22836 25891 22888 25900
rect 22836 25857 22845 25891
rect 22845 25857 22879 25891
rect 22879 25857 22888 25891
rect 22836 25848 22888 25857
rect 24124 25891 24176 25900
rect 24124 25857 24133 25891
rect 24133 25857 24167 25891
rect 24167 25857 24176 25891
rect 24124 25848 24176 25857
rect 23112 25780 23164 25832
rect 24400 25823 24452 25832
rect 24400 25789 24409 25823
rect 24409 25789 24443 25823
rect 24443 25789 24452 25823
rect 24400 25780 24452 25789
rect 22836 25644 22888 25696
rect 23020 25687 23072 25696
rect 23020 25653 23029 25687
rect 23029 25653 23063 25687
rect 23063 25653 23072 25687
rect 23020 25644 23072 25653
rect 25504 25644 25556 25696
rect 25964 25848 26016 25900
rect 33232 25780 33284 25832
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 4896 25304 4948 25356
rect 4068 25236 4120 25288
rect 5632 25440 5684 25492
rect 8024 25483 8076 25492
rect 8024 25449 8033 25483
rect 8033 25449 8067 25483
rect 8067 25449 8076 25483
rect 8024 25440 8076 25449
rect 10140 25483 10192 25492
rect 10140 25449 10149 25483
rect 10149 25449 10183 25483
rect 10183 25449 10192 25483
rect 10140 25440 10192 25449
rect 9956 25304 10008 25356
rect 10692 25440 10744 25492
rect 10784 25440 10836 25492
rect 11796 25483 11848 25492
rect 11796 25449 11805 25483
rect 11805 25449 11839 25483
rect 11839 25449 11848 25483
rect 11796 25440 11848 25449
rect 12624 25483 12676 25492
rect 12624 25449 12633 25483
rect 12633 25449 12667 25483
rect 12667 25449 12676 25483
rect 12624 25440 12676 25449
rect 12992 25440 13044 25492
rect 15844 25440 15896 25492
rect 20168 25483 20220 25492
rect 20168 25449 20177 25483
rect 20177 25449 20211 25483
rect 20211 25449 20220 25483
rect 20168 25440 20220 25449
rect 12532 25372 12584 25424
rect 11704 25347 11756 25356
rect 11704 25313 11713 25347
rect 11713 25313 11747 25347
rect 11747 25313 11756 25347
rect 11704 25304 11756 25313
rect 12164 25347 12216 25356
rect 12164 25313 12173 25347
rect 12173 25313 12207 25347
rect 12207 25313 12216 25347
rect 12164 25304 12216 25313
rect 6920 25236 6972 25288
rect 7012 25236 7064 25288
rect 7288 25279 7340 25288
rect 7288 25245 7297 25279
rect 7297 25245 7331 25279
rect 7331 25245 7340 25279
rect 7288 25236 7340 25245
rect 7380 25279 7432 25288
rect 7380 25245 7389 25279
rect 7389 25245 7423 25279
rect 7423 25245 7432 25279
rect 7380 25236 7432 25245
rect 7840 25279 7892 25288
rect 7840 25245 7849 25279
rect 7849 25245 7883 25279
rect 7883 25245 7892 25279
rect 7840 25236 7892 25245
rect 6184 25211 6236 25220
rect 6184 25177 6193 25211
rect 6193 25177 6227 25211
rect 6227 25177 6236 25211
rect 6184 25168 6236 25177
rect 7932 25168 7984 25220
rect 10140 25168 10192 25220
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 6092 25100 6144 25152
rect 7472 25100 7524 25152
rect 7656 25143 7708 25152
rect 7656 25109 7665 25143
rect 7665 25109 7699 25143
rect 7699 25109 7708 25143
rect 7656 25100 7708 25109
rect 8208 25100 8260 25152
rect 11152 25168 11204 25220
rect 11796 25236 11848 25288
rect 11612 25211 11664 25220
rect 11612 25177 11621 25211
rect 11621 25177 11655 25211
rect 11655 25177 11664 25211
rect 11612 25168 11664 25177
rect 12532 25279 12584 25288
rect 12532 25245 12541 25279
rect 12541 25245 12575 25279
rect 12575 25245 12584 25279
rect 12532 25236 12584 25245
rect 15384 25236 15436 25288
rect 15660 25372 15712 25424
rect 16396 25372 16448 25424
rect 18420 25372 18472 25424
rect 18604 25415 18656 25424
rect 18604 25381 18613 25415
rect 18613 25381 18647 25415
rect 18647 25381 18656 25415
rect 18604 25372 18656 25381
rect 20444 25440 20496 25492
rect 20996 25440 21048 25492
rect 24400 25440 24452 25492
rect 11888 25100 11940 25152
rect 12072 25100 12124 25152
rect 13176 25100 13228 25152
rect 15108 25143 15160 25152
rect 15108 25109 15117 25143
rect 15117 25109 15151 25143
rect 15151 25109 15160 25143
rect 15108 25100 15160 25109
rect 15476 25100 15528 25152
rect 16212 25279 16264 25288
rect 16212 25245 16221 25279
rect 16221 25245 16255 25279
rect 16255 25245 16264 25279
rect 16212 25236 16264 25245
rect 17592 25168 17644 25220
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 20904 25304 20956 25356
rect 23020 25372 23072 25424
rect 19340 25236 19392 25288
rect 20352 25279 20404 25288
rect 20352 25245 20361 25279
rect 20361 25245 20395 25279
rect 20395 25245 20404 25279
rect 20352 25236 20404 25245
rect 19432 25168 19484 25220
rect 19984 25168 20036 25220
rect 20536 25236 20588 25288
rect 20812 25279 20864 25288
rect 20812 25245 20821 25279
rect 20821 25245 20855 25279
rect 20855 25245 20864 25279
rect 20812 25236 20864 25245
rect 20996 25236 21048 25288
rect 20812 25100 20864 25152
rect 23112 25236 23164 25288
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 33140 25279 33192 25288
rect 33140 25245 33149 25279
rect 33149 25245 33183 25279
rect 33183 25245 33192 25279
rect 33140 25236 33192 25245
rect 34336 25211 34388 25220
rect 34336 25177 34345 25211
rect 34345 25177 34379 25211
rect 34379 25177 34388 25211
rect 34336 25168 34388 25177
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 7012 24896 7064 24948
rect 7288 24896 7340 24948
rect 7932 24896 7984 24948
rect 11152 24939 11204 24948
rect 11152 24905 11161 24939
rect 11161 24905 11195 24939
rect 11195 24905 11204 24939
rect 11152 24896 11204 24905
rect 11704 24896 11756 24948
rect 12072 24939 12124 24948
rect 12072 24905 12081 24939
rect 12081 24905 12115 24939
rect 12115 24905 12124 24939
rect 12072 24896 12124 24905
rect 12624 24896 12676 24948
rect 13544 24896 13596 24948
rect 7840 24828 7892 24880
rect 9956 24828 10008 24880
rect 5448 24760 5500 24812
rect 6920 24803 6972 24812
rect 6920 24769 6929 24803
rect 6929 24769 6963 24803
rect 6963 24769 6972 24803
rect 6920 24760 6972 24769
rect 7472 24803 7524 24812
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 9220 24803 9272 24812
rect 9220 24769 9229 24803
rect 9229 24769 9263 24803
rect 9263 24769 9272 24803
rect 9220 24760 9272 24769
rect 10784 24760 10836 24812
rect 13176 24828 13228 24880
rect 10508 24692 10560 24744
rect 11612 24692 11664 24744
rect 13360 24760 13412 24812
rect 15108 24896 15160 24948
rect 15384 24896 15436 24948
rect 19340 24896 19392 24948
rect 20996 24939 21048 24948
rect 20996 24905 21005 24939
rect 21005 24905 21039 24939
rect 21039 24905 21048 24939
rect 20996 24896 21048 24905
rect 14556 24803 14608 24812
rect 13820 24692 13872 24744
rect 14556 24769 14565 24803
rect 14565 24769 14599 24803
rect 14599 24769 14608 24803
rect 14556 24760 14608 24769
rect 14096 24735 14148 24744
rect 14096 24701 14105 24735
rect 14105 24701 14139 24735
rect 14139 24701 14148 24735
rect 14096 24692 14148 24701
rect 11336 24624 11388 24676
rect 13360 24624 13412 24676
rect 13728 24667 13780 24676
rect 13728 24633 13737 24667
rect 13737 24633 13771 24667
rect 13771 24633 13780 24667
rect 13728 24624 13780 24633
rect 5172 24556 5224 24608
rect 6092 24599 6144 24608
rect 6092 24565 6101 24599
rect 6101 24565 6135 24599
rect 6135 24565 6144 24599
rect 6092 24556 6144 24565
rect 14096 24556 14148 24608
rect 15016 24760 15068 24812
rect 15476 24803 15528 24812
rect 15476 24769 15485 24803
rect 15485 24769 15519 24803
rect 15519 24769 15528 24803
rect 15476 24760 15528 24769
rect 15660 24803 15712 24812
rect 15660 24769 15673 24803
rect 15673 24769 15712 24803
rect 15660 24760 15712 24769
rect 16212 24803 16264 24812
rect 16212 24769 16221 24803
rect 16221 24769 16255 24803
rect 16255 24769 16264 24803
rect 16212 24760 16264 24769
rect 19432 24828 19484 24880
rect 19340 24760 19392 24812
rect 16120 24692 16172 24744
rect 19800 24692 19852 24744
rect 19984 24624 20036 24676
rect 20904 24735 20956 24744
rect 20904 24701 20913 24735
rect 20913 24701 20947 24735
rect 20947 24701 20956 24735
rect 20904 24692 20956 24701
rect 16120 24599 16172 24608
rect 16120 24565 16129 24599
rect 16129 24565 16163 24599
rect 16163 24565 16172 24599
rect 16120 24556 16172 24565
rect 18512 24556 18564 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8852 24352 8904 24404
rect 940 24148 992 24200
rect 3608 24148 3660 24200
rect 4068 24148 4120 24200
rect 8024 24284 8076 24336
rect 11796 24352 11848 24404
rect 11888 24395 11940 24404
rect 11888 24361 11897 24395
rect 11897 24361 11931 24395
rect 11931 24361 11940 24395
rect 11888 24352 11940 24361
rect 11980 24352 12032 24404
rect 12440 24352 12492 24404
rect 12716 24352 12768 24404
rect 12808 24352 12860 24404
rect 13728 24352 13780 24404
rect 9220 24259 9272 24268
rect 9220 24225 9229 24259
rect 9229 24225 9263 24259
rect 9263 24225 9272 24259
rect 9220 24216 9272 24225
rect 5172 24080 5224 24132
rect 8024 24191 8076 24200
rect 8024 24157 8033 24191
rect 8033 24157 8067 24191
rect 8067 24157 8076 24191
rect 8024 24148 8076 24157
rect 8484 24148 8536 24200
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 11428 24191 11480 24200
rect 11428 24157 11437 24191
rect 11437 24157 11471 24191
rect 11471 24157 11480 24191
rect 11428 24148 11480 24157
rect 12256 24284 12308 24336
rect 15108 24352 15160 24404
rect 16120 24352 16172 24404
rect 17592 24395 17644 24404
rect 17592 24361 17601 24395
rect 17601 24361 17635 24395
rect 17635 24361 17644 24395
rect 17592 24352 17644 24361
rect 18512 24395 18564 24404
rect 18512 24361 18521 24395
rect 18521 24361 18555 24395
rect 18555 24361 18564 24395
rect 18512 24352 18564 24361
rect 18604 24395 18656 24404
rect 18604 24361 18613 24395
rect 18613 24361 18647 24395
rect 18647 24361 18656 24395
rect 18604 24352 18656 24361
rect 24124 24395 24176 24404
rect 24124 24361 24133 24395
rect 24133 24361 24167 24395
rect 24167 24361 24176 24395
rect 24124 24352 24176 24361
rect 7288 24080 7340 24132
rect 9680 24080 9732 24132
rect 10508 24080 10560 24132
rect 11980 24148 12032 24200
rect 7104 24012 7156 24064
rect 7380 24012 7432 24064
rect 9496 24055 9548 24064
rect 9496 24021 9505 24055
rect 9505 24021 9539 24055
rect 9539 24021 9548 24055
rect 9496 24012 9548 24021
rect 11888 24080 11940 24132
rect 12348 24216 12400 24268
rect 15660 24327 15712 24336
rect 15660 24293 15669 24327
rect 15669 24293 15703 24327
rect 15703 24293 15712 24327
rect 15660 24284 15712 24293
rect 12624 24191 12676 24200
rect 12624 24157 12633 24191
rect 12633 24157 12667 24191
rect 12667 24157 12676 24191
rect 12624 24148 12676 24157
rect 16764 24216 16816 24268
rect 13084 24148 13136 24200
rect 12716 24123 12768 24132
rect 12716 24089 12725 24123
rect 12725 24089 12759 24123
rect 12759 24089 12768 24123
rect 13268 24191 13320 24200
rect 13268 24157 13277 24191
rect 13277 24157 13311 24191
rect 13311 24157 13320 24191
rect 13268 24148 13320 24157
rect 12716 24080 12768 24089
rect 12808 24012 12860 24064
rect 13544 24148 13596 24200
rect 14924 24148 14976 24200
rect 15200 24191 15252 24200
rect 15200 24157 15209 24191
rect 15209 24157 15243 24191
rect 15243 24157 15252 24191
rect 15200 24148 15252 24157
rect 14096 24123 14148 24132
rect 14096 24089 14105 24123
rect 14105 24089 14139 24123
rect 14139 24089 14148 24123
rect 14096 24080 14148 24089
rect 16856 24148 16908 24200
rect 24676 24123 24728 24132
rect 24676 24089 24685 24123
rect 24685 24089 24719 24123
rect 24719 24089 24728 24123
rect 24676 24080 24728 24089
rect 24952 24080 25004 24132
rect 14004 24012 14056 24064
rect 14464 24055 14516 24064
rect 14464 24021 14473 24055
rect 14473 24021 14507 24055
rect 14507 24021 14516 24055
rect 14464 24012 14516 24021
rect 18144 24012 18196 24064
rect 33140 24012 33192 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 9220 23808 9272 23860
rect 12716 23808 12768 23860
rect 4988 23740 5040 23792
rect 6184 23672 6236 23724
rect 6920 23740 6972 23792
rect 7288 23740 7340 23792
rect 6828 23672 6880 23724
rect 7656 23715 7708 23724
rect 7656 23681 7665 23715
rect 7665 23681 7699 23715
rect 7699 23681 7708 23715
rect 7656 23672 7708 23681
rect 8024 23715 8076 23724
rect 8024 23681 8033 23715
rect 8033 23681 8067 23715
rect 8067 23681 8076 23715
rect 8024 23672 8076 23681
rect 3608 23604 3660 23656
rect 4620 23604 4672 23656
rect 6000 23647 6052 23656
rect 6000 23613 6009 23647
rect 6009 23613 6043 23647
rect 6043 23613 6052 23647
rect 6000 23604 6052 23613
rect 8208 23604 8260 23656
rect 9772 23672 9824 23724
rect 10416 23672 10468 23724
rect 11428 23672 11480 23724
rect 12072 23672 12124 23724
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 10508 23536 10560 23588
rect 11980 23536 12032 23588
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 13728 23808 13780 23860
rect 14004 23808 14056 23860
rect 14464 23808 14516 23860
rect 20812 23808 20864 23860
rect 23664 23808 23716 23860
rect 24676 23808 24728 23860
rect 24952 23851 25004 23860
rect 24952 23817 24961 23851
rect 24961 23817 24995 23851
rect 24995 23817 25004 23851
rect 24952 23808 25004 23817
rect 23112 23783 23164 23792
rect 23112 23749 23121 23783
rect 23121 23749 23155 23783
rect 23155 23749 23164 23783
rect 23112 23740 23164 23749
rect 20628 23715 20680 23724
rect 20628 23681 20637 23715
rect 20637 23681 20671 23715
rect 20671 23681 20680 23715
rect 20628 23672 20680 23681
rect 21088 23715 21140 23724
rect 21088 23681 21097 23715
rect 21097 23681 21131 23715
rect 21131 23681 21140 23715
rect 21088 23672 21140 23681
rect 14096 23604 14148 23656
rect 20444 23647 20496 23656
rect 20444 23613 20453 23647
rect 20453 23613 20487 23647
rect 20487 23613 20496 23647
rect 20444 23604 20496 23613
rect 21456 23604 21508 23656
rect 21916 23647 21968 23656
rect 21916 23613 21925 23647
rect 21925 23613 21959 23647
rect 21959 23613 21968 23647
rect 21916 23604 21968 23613
rect 13268 23536 13320 23588
rect 13544 23536 13596 23588
rect 21180 23536 21232 23588
rect 23020 23715 23072 23724
rect 23020 23681 23029 23715
rect 23029 23681 23063 23715
rect 23063 23681 23072 23715
rect 23020 23672 23072 23681
rect 23388 23672 23440 23724
rect 11888 23468 11940 23520
rect 23020 23468 23072 23520
rect 25504 23468 25556 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4988 23264 5040 23316
rect 5448 23264 5500 23316
rect 7104 23307 7156 23316
rect 7104 23273 7113 23307
rect 7113 23273 7147 23307
rect 7147 23273 7156 23307
rect 7104 23264 7156 23273
rect 8208 23264 8260 23316
rect 13084 23307 13136 23316
rect 13084 23273 13093 23307
rect 13093 23273 13127 23307
rect 13127 23273 13136 23307
rect 13084 23264 13136 23273
rect 15844 23264 15896 23316
rect 16856 23264 16908 23316
rect 20444 23264 20496 23316
rect 21916 23264 21968 23316
rect 23020 23264 23072 23316
rect 12624 23196 12676 23248
rect 6828 23171 6880 23180
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 6920 23103 6972 23112
rect 6920 23069 6929 23103
rect 6929 23069 6963 23103
rect 6963 23069 6972 23103
rect 6920 23060 6972 23069
rect 7932 23103 7984 23112
rect 7932 23069 7941 23103
rect 7941 23069 7975 23103
rect 7975 23069 7984 23103
rect 7932 23060 7984 23069
rect 9772 23103 9824 23112
rect 9772 23069 9781 23103
rect 9781 23069 9815 23103
rect 9815 23069 9824 23103
rect 9772 23060 9824 23069
rect 10416 23103 10468 23112
rect 10416 23069 10425 23103
rect 10425 23069 10459 23103
rect 10459 23069 10468 23103
rect 10416 23060 10468 23069
rect 12072 23103 12124 23112
rect 12072 23069 12081 23103
rect 12081 23069 12115 23103
rect 12115 23069 12124 23103
rect 12072 23060 12124 23069
rect 12256 23060 12308 23112
rect 12808 23128 12860 23180
rect 13360 23103 13412 23112
rect 13360 23069 13369 23103
rect 13369 23069 13403 23103
rect 13403 23069 13412 23103
rect 13360 23060 13412 23069
rect 5632 22967 5684 22976
rect 5632 22933 5641 22967
rect 5641 22933 5675 22967
rect 5675 22933 5684 22967
rect 6092 22967 6144 22976
rect 5632 22924 5684 22933
rect 6092 22933 6101 22967
rect 6101 22933 6135 22967
rect 6135 22933 6144 22967
rect 6092 22924 6144 22933
rect 8300 22967 8352 22976
rect 8300 22933 8309 22967
rect 8309 22933 8343 22967
rect 8343 22933 8352 22967
rect 8300 22924 8352 22933
rect 8576 22924 8628 22976
rect 12716 23035 12768 23044
rect 12716 23001 12725 23035
rect 12725 23001 12759 23035
rect 12759 23001 12768 23035
rect 12716 22992 12768 23001
rect 12808 22992 12860 23044
rect 15292 23171 15344 23180
rect 15292 23137 15301 23171
rect 15301 23137 15335 23171
rect 15335 23137 15344 23171
rect 15292 23128 15344 23137
rect 16672 23171 16724 23180
rect 16672 23137 16681 23171
rect 16681 23137 16715 23171
rect 16715 23137 16724 23171
rect 16672 23128 16724 23137
rect 19432 23128 19484 23180
rect 13268 22967 13320 22976
rect 13268 22933 13277 22967
rect 13277 22933 13311 22967
rect 13311 22933 13320 22967
rect 13268 22924 13320 22933
rect 14832 22924 14884 22976
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 19984 23060 20036 23112
rect 20444 23060 20496 23112
rect 21088 23196 21140 23248
rect 21180 23171 21232 23180
rect 21180 23137 21189 23171
rect 21189 23137 21223 23171
rect 21223 23137 21232 23171
rect 21180 23128 21232 23137
rect 22100 23060 22152 23112
rect 22652 23060 22704 23112
rect 33140 23103 33192 23112
rect 33140 23069 33149 23103
rect 33149 23069 33183 23103
rect 33183 23069 33192 23103
rect 33140 23060 33192 23069
rect 15844 22924 15896 22976
rect 17132 22967 17184 22976
rect 17132 22933 17141 22967
rect 17141 22933 17175 22967
rect 17175 22933 17184 22967
rect 17132 22924 17184 22933
rect 20628 23035 20680 23044
rect 20628 23001 20637 23035
rect 20637 23001 20671 23035
rect 20671 23001 20680 23035
rect 20628 22992 20680 23001
rect 34888 22992 34940 23044
rect 20720 22924 20772 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 5448 22720 5500 22772
rect 3884 22695 3936 22704
rect 3884 22661 3893 22695
rect 3893 22661 3927 22695
rect 3927 22661 3936 22695
rect 3884 22652 3936 22661
rect 9496 22720 9548 22772
rect 8852 22652 8904 22704
rect 6828 22584 6880 22636
rect 6920 22584 6972 22636
rect 7932 22627 7984 22636
rect 7932 22593 7941 22627
rect 7941 22593 7975 22627
rect 7975 22593 7984 22627
rect 7932 22584 7984 22593
rect 8576 22627 8628 22636
rect 8576 22593 8585 22627
rect 8585 22593 8619 22627
rect 8619 22593 8628 22627
rect 8576 22584 8628 22593
rect 8760 22584 8812 22636
rect 12072 22652 12124 22704
rect 12716 22720 12768 22772
rect 15016 22720 15068 22772
rect 16028 22720 16080 22772
rect 17132 22720 17184 22772
rect 19340 22763 19392 22772
rect 19340 22729 19349 22763
rect 19349 22729 19383 22763
rect 19383 22729 19392 22763
rect 19340 22720 19392 22729
rect 19432 22720 19484 22772
rect 13360 22584 13412 22636
rect 14556 22584 14608 22636
rect 14648 22627 14700 22636
rect 14648 22593 14657 22627
rect 14657 22593 14691 22627
rect 14691 22593 14700 22627
rect 14648 22584 14700 22593
rect 3608 22559 3660 22568
rect 3608 22525 3617 22559
rect 3617 22525 3651 22559
rect 3651 22525 3660 22559
rect 3608 22516 3660 22525
rect 6276 22516 6328 22568
rect 8300 22448 8352 22500
rect 9588 22516 9640 22568
rect 11980 22516 12032 22568
rect 14464 22559 14516 22568
rect 14464 22525 14473 22559
rect 14473 22525 14507 22559
rect 14507 22525 14516 22559
rect 14464 22516 14516 22525
rect 9680 22448 9732 22500
rect 10232 22448 10284 22500
rect 12716 22448 12768 22500
rect 14832 22516 14884 22568
rect 15384 22627 15436 22636
rect 15384 22593 15393 22627
rect 15393 22593 15427 22627
rect 15427 22593 15436 22627
rect 15384 22584 15436 22593
rect 15476 22584 15528 22636
rect 15108 22559 15160 22568
rect 15108 22525 15117 22559
rect 15117 22525 15151 22559
rect 15151 22525 15160 22559
rect 15108 22516 15160 22525
rect 15844 22559 15896 22568
rect 15844 22525 15853 22559
rect 15853 22525 15887 22559
rect 15887 22525 15896 22559
rect 15844 22516 15896 22525
rect 17224 22516 17276 22568
rect 18328 22516 18380 22568
rect 18788 22559 18840 22568
rect 18788 22525 18797 22559
rect 18797 22525 18831 22559
rect 18831 22525 18840 22559
rect 18788 22516 18840 22525
rect 19984 22584 20036 22636
rect 22560 22584 22612 22636
rect 23020 22720 23072 22772
rect 23388 22763 23440 22772
rect 23388 22729 23397 22763
rect 23397 22729 23431 22763
rect 23431 22729 23440 22763
rect 23388 22720 23440 22729
rect 22928 22627 22980 22636
rect 22928 22593 22937 22627
rect 22937 22593 22971 22627
rect 22971 22593 22980 22627
rect 22928 22584 22980 22593
rect 23204 22627 23256 22636
rect 23204 22593 23213 22627
rect 23213 22593 23247 22627
rect 23247 22593 23256 22627
rect 23204 22584 23256 22593
rect 24124 22720 24176 22772
rect 33140 22720 33192 22772
rect 25504 22584 25556 22636
rect 24216 22559 24268 22568
rect 24216 22525 24225 22559
rect 24225 22525 24259 22559
rect 24259 22525 24268 22559
rect 24216 22516 24268 22525
rect 10324 22380 10376 22432
rect 14556 22380 14608 22432
rect 15108 22380 15160 22432
rect 15200 22380 15252 22432
rect 18236 22423 18288 22432
rect 18236 22389 18245 22423
rect 18245 22389 18279 22423
rect 18279 22389 18288 22423
rect 18236 22380 18288 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 5816 22219 5868 22228
rect 5816 22185 5825 22219
rect 5825 22185 5859 22219
rect 5859 22185 5868 22219
rect 5816 22176 5868 22185
rect 6000 22176 6052 22228
rect 6920 22176 6972 22228
rect 8116 22176 8168 22228
rect 9404 22176 9456 22228
rect 10324 22219 10376 22228
rect 10324 22185 10333 22219
rect 10333 22185 10367 22219
rect 10367 22185 10376 22219
rect 10324 22176 10376 22185
rect 10416 22176 10468 22228
rect 940 21972 992 22024
rect 6644 22108 6696 22160
rect 7748 22108 7800 22160
rect 8208 22108 8260 22160
rect 8576 22108 8628 22160
rect 5908 21972 5960 22024
rect 6000 22015 6052 22024
rect 6000 21981 6009 22015
rect 6009 21981 6043 22015
rect 6043 21981 6052 22015
rect 6000 21972 6052 21981
rect 6184 21972 6236 22024
rect 8116 22015 8168 22024
rect 8116 21981 8125 22015
rect 8125 21981 8159 22015
rect 8159 21981 8168 22015
rect 8116 21972 8168 21981
rect 8392 21972 8444 22024
rect 10232 22083 10284 22092
rect 10232 22049 10241 22083
rect 10241 22049 10275 22083
rect 10275 22049 10284 22083
rect 10232 22040 10284 22049
rect 10876 22151 10928 22160
rect 10876 22117 10885 22151
rect 10885 22117 10919 22151
rect 10919 22117 10928 22151
rect 10876 22108 10928 22117
rect 14832 22176 14884 22228
rect 15292 22176 15344 22228
rect 18144 22176 18196 22228
rect 19984 22176 20036 22228
rect 21456 22219 21508 22228
rect 21456 22185 21465 22219
rect 21465 22185 21499 22219
rect 21499 22185 21508 22219
rect 21456 22176 21508 22185
rect 24216 22176 24268 22228
rect 12624 22108 12676 22160
rect 13268 22108 13320 22160
rect 20168 22108 20220 22160
rect 21088 22151 21140 22160
rect 21088 22117 21097 22151
rect 21097 22117 21131 22151
rect 21131 22117 21140 22151
rect 21088 22108 21140 22117
rect 22928 22108 22980 22160
rect 9864 22015 9916 22024
rect 9864 21981 9873 22015
rect 9873 21981 9907 22015
rect 9907 21981 9916 22015
rect 9864 21972 9916 21981
rect 10600 21972 10652 22024
rect 1584 21879 1636 21888
rect 1584 21845 1593 21879
rect 1593 21845 1627 21879
rect 1627 21845 1636 21879
rect 1584 21836 1636 21845
rect 5356 21879 5408 21888
rect 5356 21845 5365 21879
rect 5365 21845 5399 21879
rect 5399 21845 5408 21879
rect 5356 21836 5408 21845
rect 7932 21836 7984 21888
rect 10048 21836 10100 21888
rect 10784 21836 10836 21888
rect 11244 21972 11296 22024
rect 12532 21972 12584 22024
rect 13084 22040 13136 22092
rect 13544 22015 13596 22024
rect 13544 21981 13553 22015
rect 13553 21981 13587 22015
rect 13587 21981 13596 22015
rect 13544 21972 13596 21981
rect 21732 22083 21784 22092
rect 21732 22049 21741 22083
rect 21741 22049 21775 22083
rect 21775 22049 21784 22083
rect 21732 22040 21784 22049
rect 14464 21972 14516 22024
rect 14740 22015 14792 22024
rect 14740 21981 14749 22015
rect 14749 21981 14783 22015
rect 14783 21981 14792 22015
rect 14740 21972 14792 21981
rect 14924 22015 14976 22024
rect 14924 21981 14933 22015
rect 14933 21981 14967 22015
rect 14967 21981 14976 22015
rect 14924 21972 14976 21981
rect 15016 22015 15068 22024
rect 15016 21981 15025 22015
rect 15025 21981 15059 22015
rect 15059 21981 15068 22015
rect 15016 21972 15068 21981
rect 15108 22015 15160 22024
rect 15108 21981 15117 22015
rect 15117 21981 15151 22015
rect 15151 21981 15160 22015
rect 15108 21972 15160 21981
rect 15476 21972 15528 22024
rect 16396 22015 16448 22024
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16396 21972 16448 21981
rect 18236 22015 18288 22024
rect 18236 21981 18245 22015
rect 18245 21981 18279 22015
rect 18279 21981 18288 22015
rect 18236 21972 18288 21981
rect 18328 21972 18380 22024
rect 18880 21972 18932 22024
rect 14556 21904 14608 21956
rect 14648 21904 14700 21956
rect 11336 21836 11388 21888
rect 12808 21879 12860 21888
rect 12808 21845 12817 21879
rect 12817 21845 12851 21879
rect 12851 21845 12860 21879
rect 12808 21836 12860 21845
rect 12900 21836 12952 21888
rect 13268 21836 13320 21888
rect 13820 21836 13872 21888
rect 15936 21836 15988 21888
rect 16212 21836 16264 21888
rect 17408 21836 17460 21888
rect 19984 21879 20036 21888
rect 19984 21845 19993 21879
rect 19993 21845 20027 21879
rect 20027 21845 20036 21879
rect 19984 21836 20036 21845
rect 20168 22015 20220 22024
rect 20168 21981 20177 22015
rect 20177 21981 20211 22015
rect 20211 21981 20220 22015
rect 20168 21972 20220 21981
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 20536 21836 20588 21888
rect 20996 21836 21048 21888
rect 23204 21972 23256 22024
rect 22468 21836 22520 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 1584 21632 1636 21684
rect 6000 21632 6052 21684
rect 4804 21564 4856 21616
rect 8668 21632 8720 21684
rect 3608 21428 3660 21480
rect 5632 21496 5684 21548
rect 6644 21539 6696 21548
rect 6644 21505 6678 21539
rect 6678 21505 6696 21539
rect 6644 21496 6696 21505
rect 5816 21471 5868 21480
rect 5816 21437 5825 21471
rect 5825 21437 5859 21471
rect 5859 21437 5868 21471
rect 6920 21539 6972 21548
rect 6920 21505 6929 21539
rect 6929 21505 6963 21539
rect 6963 21505 6972 21539
rect 6920 21496 6972 21505
rect 7932 21539 7984 21548
rect 7932 21505 7941 21539
rect 7941 21505 7975 21539
rect 7975 21505 7984 21539
rect 7932 21496 7984 21505
rect 9864 21632 9916 21684
rect 10324 21632 10376 21684
rect 9680 21564 9732 21616
rect 5816 21428 5868 21437
rect 9956 21539 10008 21548
rect 9956 21505 9965 21539
rect 9965 21505 9999 21539
rect 9999 21505 10008 21539
rect 9956 21496 10008 21505
rect 10784 21564 10836 21616
rect 12532 21632 12584 21684
rect 12992 21564 13044 21616
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 9772 21403 9824 21412
rect 9772 21369 9781 21403
rect 9781 21369 9815 21403
rect 9815 21369 9824 21403
rect 9772 21360 9824 21369
rect 9864 21403 9916 21412
rect 9864 21369 9873 21403
rect 9873 21369 9907 21403
rect 9907 21369 9916 21403
rect 9864 21360 9916 21369
rect 10416 21471 10468 21480
rect 10416 21437 10425 21471
rect 10425 21437 10459 21471
rect 10459 21437 10468 21471
rect 10416 21428 10468 21437
rect 10876 21428 10928 21480
rect 11244 21496 11296 21548
rect 8392 21292 8444 21344
rect 10140 21292 10192 21344
rect 11612 21428 11664 21480
rect 12808 21496 12860 21548
rect 13820 21564 13872 21616
rect 12900 21471 12952 21480
rect 12900 21437 12909 21471
rect 12909 21437 12943 21471
rect 12943 21437 12952 21471
rect 12900 21428 12952 21437
rect 13268 21360 13320 21412
rect 13820 21471 13872 21480
rect 13820 21437 13829 21471
rect 13829 21437 13863 21471
rect 13863 21437 13872 21471
rect 13820 21428 13872 21437
rect 14556 21632 14608 21684
rect 16212 21632 16264 21684
rect 16396 21632 16448 21684
rect 16672 21632 16724 21684
rect 17408 21675 17460 21684
rect 17408 21641 17417 21675
rect 17417 21641 17451 21675
rect 17451 21641 17460 21675
rect 17408 21632 17460 21641
rect 20996 21675 21048 21684
rect 20996 21641 21005 21675
rect 21005 21641 21039 21675
rect 21039 21641 21048 21675
rect 20996 21632 21048 21641
rect 21088 21632 21140 21684
rect 21732 21632 21784 21684
rect 23204 21632 23256 21684
rect 14188 21496 14240 21548
rect 15384 21539 15436 21548
rect 15384 21505 15393 21539
rect 15393 21505 15427 21539
rect 15427 21505 15436 21539
rect 15384 21496 15436 21505
rect 15568 21539 15620 21548
rect 15568 21505 15577 21539
rect 15577 21505 15611 21539
rect 15611 21505 15620 21539
rect 15568 21496 15620 21505
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 17592 21564 17644 21616
rect 16856 21496 16908 21548
rect 22468 21607 22520 21616
rect 22468 21573 22477 21607
rect 22477 21573 22511 21607
rect 22511 21573 22520 21607
rect 22468 21564 22520 21573
rect 22560 21564 22612 21616
rect 14372 21471 14424 21480
rect 14372 21437 14381 21471
rect 14381 21437 14415 21471
rect 14415 21437 14424 21471
rect 14372 21428 14424 21437
rect 15660 21428 15712 21480
rect 17592 21428 17644 21480
rect 20720 21496 20772 21548
rect 17408 21360 17460 21412
rect 20996 21496 21048 21548
rect 23296 21539 23348 21548
rect 23296 21505 23305 21539
rect 23305 21505 23339 21539
rect 23339 21505 23348 21539
rect 23296 21496 23348 21505
rect 21272 21428 21324 21480
rect 13728 21292 13780 21344
rect 13912 21292 13964 21344
rect 18144 21292 18196 21344
rect 18236 21335 18288 21344
rect 18236 21301 18245 21335
rect 18245 21301 18279 21335
rect 18279 21301 18288 21335
rect 18236 21292 18288 21301
rect 22836 21335 22888 21344
rect 22836 21301 22845 21335
rect 22845 21301 22879 21335
rect 22879 21301 22888 21335
rect 22836 21292 22888 21301
rect 23204 21292 23256 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4804 21088 4856 21140
rect 5448 21088 5500 21140
rect 6184 21020 6236 21072
rect 6552 21063 6604 21072
rect 6552 21029 6561 21063
rect 6561 21029 6595 21063
rect 6595 21029 6604 21063
rect 6552 21020 6604 21029
rect 9312 21020 9364 21072
rect 10232 21020 10284 21072
rect 12992 21088 13044 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 13268 21088 13320 21140
rect 13544 21131 13596 21140
rect 13544 21097 13553 21131
rect 13553 21097 13587 21131
rect 13587 21097 13596 21131
rect 13544 21088 13596 21097
rect 13912 21088 13964 21140
rect 14372 21088 14424 21140
rect 14556 21131 14608 21140
rect 14556 21097 14565 21131
rect 14565 21097 14599 21131
rect 14599 21097 14608 21131
rect 14556 21088 14608 21097
rect 15016 21088 15068 21140
rect 15568 21131 15620 21140
rect 15568 21097 15577 21131
rect 15577 21097 15611 21131
rect 15611 21097 15620 21131
rect 15568 21088 15620 21097
rect 16856 21088 16908 21140
rect 18236 21088 18288 21140
rect 19984 21088 20036 21140
rect 20536 21131 20588 21140
rect 20536 21097 20545 21131
rect 20545 21097 20579 21131
rect 20579 21097 20588 21131
rect 20536 21088 20588 21097
rect 22836 21088 22888 21140
rect 24124 21131 24176 21140
rect 24124 21097 24133 21131
rect 24133 21097 24167 21131
rect 24167 21097 24176 21131
rect 24124 21088 24176 21097
rect 11336 21020 11388 21072
rect 5356 20952 5408 21004
rect 8944 20995 8996 21004
rect 8944 20961 8953 20995
rect 8953 20961 8987 20995
rect 8987 20961 8996 20995
rect 8944 20952 8996 20961
rect 9496 20952 9548 21004
rect 6276 20927 6328 20936
rect 6276 20893 6285 20927
rect 6285 20893 6319 20927
rect 6319 20893 6328 20927
rect 6276 20884 6328 20893
rect 6736 20884 6788 20936
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 9772 20884 9824 20936
rect 6000 20816 6052 20868
rect 8668 20816 8720 20868
rect 9496 20748 9548 20800
rect 9956 20884 10008 20936
rect 10140 20884 10192 20936
rect 10876 20952 10928 21004
rect 10968 20952 11020 21004
rect 13268 20884 13320 20936
rect 13544 20884 13596 20936
rect 14188 20927 14240 20936
rect 9956 20791 10008 20800
rect 9956 20757 9965 20791
rect 9965 20757 9999 20791
rect 9999 20757 10008 20791
rect 9956 20748 10008 20757
rect 10324 20748 10376 20800
rect 11244 20816 11296 20868
rect 14188 20893 14197 20927
rect 14197 20893 14231 20927
rect 14231 20893 14240 20927
rect 14188 20884 14240 20893
rect 14924 20995 14976 21004
rect 14924 20961 14933 20995
rect 14933 20961 14967 20995
rect 14967 20961 14976 20995
rect 14924 20952 14976 20961
rect 15384 20995 15436 21004
rect 15384 20961 15393 20995
rect 15393 20961 15427 20995
rect 15427 20961 15436 20995
rect 15384 20952 15436 20961
rect 16028 20995 16080 21004
rect 16028 20961 16037 20995
rect 16037 20961 16071 20995
rect 16071 20961 16080 20995
rect 16028 20952 16080 20961
rect 15660 20884 15712 20936
rect 17684 20884 17736 20936
rect 13728 20859 13780 20868
rect 13728 20825 13755 20859
rect 13755 20825 13780 20859
rect 13728 20816 13780 20825
rect 18144 20884 18196 20936
rect 19432 20884 19484 20936
rect 19984 20952 20036 21004
rect 20076 20927 20128 20936
rect 20076 20893 20085 20927
rect 20085 20893 20119 20927
rect 20119 20893 20128 20927
rect 20076 20884 20128 20893
rect 13360 20748 13412 20800
rect 14004 20748 14056 20800
rect 19248 20816 19300 20868
rect 17960 20748 18012 20800
rect 19156 20748 19208 20800
rect 24124 20884 24176 20936
rect 25136 20816 25188 20868
rect 23204 20748 23256 20800
rect 34336 20859 34388 20868
rect 34336 20825 34345 20859
rect 34345 20825 34379 20859
rect 34379 20825 34388 20859
rect 34336 20816 34388 20825
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 9312 20544 9364 20596
rect 9680 20544 9732 20596
rect 9772 20544 9824 20596
rect 8668 20476 8720 20528
rect 8944 20476 8996 20528
rect 7104 20408 7156 20460
rect 7288 20451 7340 20460
rect 7288 20417 7297 20451
rect 7297 20417 7331 20451
rect 7331 20417 7340 20451
rect 7288 20408 7340 20417
rect 10416 20544 10468 20596
rect 10508 20544 10560 20596
rect 9772 20451 9824 20460
rect 9772 20417 9781 20451
rect 9781 20417 9815 20451
rect 9815 20417 9824 20451
rect 9772 20408 9824 20417
rect 9496 20340 9548 20392
rect 9680 20340 9732 20392
rect 10232 20340 10284 20392
rect 12348 20544 12400 20596
rect 14924 20544 14976 20596
rect 18236 20544 18288 20596
rect 18880 20587 18932 20596
rect 18880 20553 18889 20587
rect 18889 20553 18923 20587
rect 18923 20553 18932 20587
rect 18880 20544 18932 20553
rect 19432 20544 19484 20596
rect 19984 20544 20036 20596
rect 25136 20544 25188 20596
rect 25412 20587 25464 20596
rect 25412 20553 25421 20587
rect 25421 20553 25455 20587
rect 25455 20553 25464 20587
rect 25412 20544 25464 20553
rect 10784 20476 10836 20528
rect 12900 20476 12952 20528
rect 15108 20476 15160 20528
rect 11704 20408 11756 20460
rect 12808 20408 12860 20460
rect 11612 20340 11664 20392
rect 10876 20315 10928 20324
rect 10876 20281 10885 20315
rect 10885 20281 10919 20315
rect 10919 20281 10928 20315
rect 10876 20272 10928 20281
rect 9128 20204 9180 20256
rect 12256 20272 12308 20324
rect 15660 20408 15712 20460
rect 16028 20408 16080 20460
rect 19156 20476 19208 20528
rect 17684 20383 17736 20392
rect 17684 20349 17693 20383
rect 17693 20349 17727 20383
rect 17727 20349 17736 20383
rect 17684 20340 17736 20349
rect 17960 20340 18012 20392
rect 18144 20383 18196 20392
rect 18144 20349 18153 20383
rect 18153 20349 18187 20383
rect 18187 20349 18196 20383
rect 18144 20340 18196 20349
rect 12164 20204 12216 20256
rect 18236 20272 18288 20324
rect 19248 20340 19300 20392
rect 19524 20408 19576 20460
rect 19984 20408 20036 20460
rect 13360 20204 13412 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 6276 20000 6328 20052
rect 9312 20000 9364 20052
rect 9772 20043 9824 20052
rect 9772 20009 9781 20043
rect 9781 20009 9815 20043
rect 9815 20009 9824 20043
rect 9772 20000 9824 20009
rect 10324 20000 10376 20052
rect 5816 19907 5868 19916
rect 5816 19873 5825 19907
rect 5825 19873 5859 19907
rect 5859 19873 5868 19907
rect 5816 19864 5868 19873
rect 940 19796 992 19848
rect 6000 19796 6052 19848
rect 6092 19839 6144 19848
rect 6092 19805 6101 19839
rect 6101 19805 6135 19839
rect 6135 19805 6144 19839
rect 6092 19796 6144 19805
rect 6276 19839 6328 19848
rect 6276 19805 6285 19839
rect 6285 19805 6319 19839
rect 6319 19805 6328 19839
rect 6276 19796 6328 19805
rect 7104 19839 7156 19848
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 7288 19796 7340 19848
rect 8944 19796 8996 19848
rect 9220 19796 9272 19848
rect 10600 19932 10652 19984
rect 11612 20043 11664 20052
rect 11612 20009 11621 20043
rect 11621 20009 11655 20043
rect 11655 20009 11664 20043
rect 11612 20000 11664 20009
rect 10232 19864 10284 19916
rect 11796 19932 11848 19984
rect 12716 20000 12768 20052
rect 12532 19975 12584 19984
rect 12532 19941 12541 19975
rect 12541 19941 12575 19975
rect 12575 19941 12584 19975
rect 12532 19932 12584 19941
rect 13268 19932 13320 19984
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 11152 19839 11204 19848
rect 11152 19805 11161 19839
rect 11161 19805 11195 19839
rect 11195 19805 11204 19839
rect 11152 19796 11204 19805
rect 12348 19864 12400 19916
rect 12808 19864 12860 19916
rect 11980 19839 12032 19848
rect 11980 19805 11989 19839
rect 11989 19805 12023 19839
rect 12023 19805 12032 19839
rect 11980 19796 12032 19805
rect 12164 19839 12216 19848
rect 12164 19805 12173 19839
rect 12173 19805 12207 19839
rect 12207 19805 12216 19839
rect 12164 19796 12216 19805
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 16948 19975 17000 19984
rect 16948 19941 16957 19975
rect 16957 19941 16991 19975
rect 16991 19941 17000 19975
rect 16948 19932 17000 19941
rect 13636 19907 13688 19916
rect 13636 19873 13645 19907
rect 13645 19873 13679 19907
rect 13679 19873 13688 19907
rect 13636 19864 13688 19873
rect 12624 19796 12676 19805
rect 4620 19660 4672 19712
rect 8116 19660 8168 19712
rect 9128 19660 9180 19712
rect 12072 19728 12124 19780
rect 14096 19796 14148 19848
rect 18052 19796 18104 19848
rect 11060 19660 11112 19712
rect 11244 19660 11296 19712
rect 11612 19660 11664 19712
rect 12348 19660 12400 19712
rect 16672 19728 16724 19780
rect 18236 19728 18288 19780
rect 18972 19728 19024 19780
rect 13544 19660 13596 19712
rect 17040 19703 17092 19712
rect 17040 19669 17049 19703
rect 17049 19669 17083 19703
rect 17083 19669 17092 19703
rect 17040 19660 17092 19669
rect 19432 19660 19484 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 6276 19456 6328 19508
rect 8116 19456 8168 19508
rect 11704 19456 11756 19508
rect 5816 19388 5868 19440
rect 3608 19320 3660 19372
rect 5908 19320 5960 19372
rect 9680 19388 9732 19440
rect 10876 19388 10928 19440
rect 8024 19363 8076 19372
rect 8024 19329 8033 19363
rect 8033 19329 8067 19363
rect 8067 19329 8076 19363
rect 8024 19320 8076 19329
rect 9496 19295 9548 19346
rect 10600 19320 10652 19372
rect 11060 19363 11112 19372
rect 11060 19329 11069 19363
rect 11069 19329 11103 19363
rect 11103 19329 11112 19363
rect 11060 19320 11112 19329
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 11704 19320 11756 19372
rect 12256 19456 12308 19508
rect 9496 19294 9505 19295
rect 9505 19294 9539 19295
rect 9539 19294 9548 19295
rect 12256 19363 12308 19372
rect 12256 19329 12265 19363
rect 12265 19329 12299 19363
rect 12299 19329 12308 19363
rect 12256 19320 12308 19329
rect 12348 19320 12400 19372
rect 12624 19388 12676 19440
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 13544 19363 13596 19372
rect 13544 19329 13553 19363
rect 13553 19329 13587 19363
rect 13587 19329 13596 19363
rect 13544 19320 13596 19329
rect 17040 19456 17092 19508
rect 17960 19456 18012 19508
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 15384 19320 15436 19372
rect 16580 19320 16632 19372
rect 17592 19388 17644 19440
rect 6092 19184 6144 19236
rect 6460 19184 6512 19236
rect 8024 19184 8076 19236
rect 12532 19184 12584 19236
rect 17132 19252 17184 19304
rect 18236 19320 18288 19372
rect 18512 19320 18564 19372
rect 19432 19320 19484 19372
rect 19708 19320 19760 19372
rect 18972 19295 19024 19304
rect 13268 19227 13320 19236
rect 13268 19193 13277 19227
rect 13277 19193 13311 19227
rect 13311 19193 13320 19227
rect 13268 19184 13320 19193
rect 13544 19184 13596 19236
rect 16764 19227 16816 19236
rect 16764 19193 16773 19227
rect 16773 19193 16807 19227
rect 16807 19193 16816 19227
rect 16764 19184 16816 19193
rect 16948 19184 17000 19236
rect 18972 19261 18981 19295
rect 18981 19261 19015 19295
rect 19015 19261 19024 19295
rect 18972 19252 19024 19261
rect 6000 19116 6052 19168
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13452 19116 13504 19125
rect 17776 19116 17828 19168
rect 19340 19159 19392 19168
rect 19340 19125 19349 19159
rect 19349 19125 19383 19159
rect 19383 19125 19392 19159
rect 19340 19116 19392 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 8024 18955 8076 18964
rect 8024 18921 8033 18955
rect 8033 18921 8067 18955
rect 8067 18921 8076 18955
rect 8024 18912 8076 18921
rect 8392 18955 8444 18964
rect 8392 18921 8401 18955
rect 8401 18921 8435 18955
rect 8435 18921 8444 18955
rect 8392 18912 8444 18921
rect 17132 18912 17184 18964
rect 17224 18955 17276 18964
rect 17224 18921 17233 18955
rect 17233 18921 17267 18955
rect 17267 18921 17276 18955
rect 17224 18912 17276 18921
rect 17684 18955 17736 18964
rect 17684 18921 17693 18955
rect 17693 18921 17727 18955
rect 17727 18921 17736 18955
rect 17684 18912 17736 18921
rect 19340 18912 19392 18964
rect 5264 18844 5316 18896
rect 6000 18844 6052 18896
rect 3608 18776 3660 18828
rect 4804 18776 4856 18828
rect 6460 18776 6512 18828
rect 5816 18708 5868 18760
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 8116 18819 8168 18828
rect 8116 18785 8125 18819
rect 8125 18785 8159 18819
rect 8159 18785 8168 18819
rect 8116 18776 8168 18785
rect 14740 18776 14792 18828
rect 16948 18819 17000 18828
rect 16948 18785 16957 18819
rect 16957 18785 16991 18819
rect 16991 18785 17000 18819
rect 16948 18776 17000 18785
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 4896 18640 4948 18692
rect 7012 18640 7064 18692
rect 7748 18683 7800 18692
rect 7748 18649 7757 18683
rect 7757 18649 7791 18683
rect 7791 18649 7800 18683
rect 7748 18640 7800 18649
rect 7564 18572 7616 18624
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 16672 18708 16724 18760
rect 17592 18844 17644 18896
rect 20996 18887 21048 18896
rect 20996 18853 21005 18887
rect 21005 18853 21039 18887
rect 21039 18853 21048 18887
rect 20996 18844 21048 18853
rect 20720 18776 20772 18828
rect 17868 18751 17920 18760
rect 17868 18717 17877 18751
rect 17877 18717 17911 18751
rect 17911 18717 17920 18751
rect 17868 18708 17920 18717
rect 19340 18708 19392 18760
rect 19708 18751 19760 18760
rect 19708 18717 19717 18751
rect 19717 18717 19751 18751
rect 19751 18717 19760 18751
rect 19708 18708 19760 18717
rect 20812 18708 20864 18760
rect 33140 18751 33192 18760
rect 33140 18717 33149 18751
rect 33149 18717 33183 18751
rect 33183 18717 33192 18751
rect 33140 18708 33192 18717
rect 10324 18572 10376 18624
rect 12624 18572 12676 18624
rect 12992 18572 13044 18624
rect 13636 18572 13688 18624
rect 14464 18572 14516 18624
rect 14556 18572 14608 18624
rect 17776 18683 17828 18692
rect 17776 18649 17785 18683
rect 17785 18649 17819 18683
rect 17819 18649 17828 18683
rect 17776 18640 17828 18649
rect 34888 18640 34940 18692
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 4896 18368 4948 18420
rect 5448 18411 5500 18420
rect 5448 18377 5457 18411
rect 5457 18377 5491 18411
rect 5491 18377 5500 18411
rect 5448 18368 5500 18377
rect 5908 18368 5960 18420
rect 7748 18368 7800 18420
rect 9404 18368 9456 18420
rect 12992 18368 13044 18420
rect 7012 18232 7064 18284
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 9036 18207 9088 18216
rect 9036 18173 9045 18207
rect 9045 18173 9079 18207
rect 9079 18173 9088 18207
rect 9036 18164 9088 18173
rect 10968 18232 11020 18284
rect 9864 18164 9916 18216
rect 10692 18207 10744 18216
rect 10692 18173 10701 18207
rect 10701 18173 10735 18207
rect 10735 18173 10744 18207
rect 10692 18164 10744 18173
rect 12624 18275 12676 18284
rect 12624 18241 12633 18275
rect 12633 18241 12667 18275
rect 12667 18241 12676 18275
rect 12624 18232 12676 18241
rect 13268 18232 13320 18284
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 14556 18368 14608 18420
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 16580 18368 16632 18420
rect 17868 18411 17920 18420
rect 17868 18377 17877 18411
rect 17877 18377 17911 18411
rect 17911 18377 17920 18411
rect 17868 18368 17920 18377
rect 9772 18096 9824 18148
rect 12624 18096 12676 18148
rect 14464 18232 14516 18284
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 15108 18232 15160 18284
rect 14280 18096 14332 18148
rect 14556 18096 14608 18148
rect 15568 18275 15620 18284
rect 15568 18241 15577 18275
rect 15577 18241 15611 18275
rect 15611 18241 15620 18275
rect 15568 18232 15620 18241
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 13820 18028 13872 18080
rect 18512 18096 18564 18148
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 5908 17824 5960 17876
rect 10692 17824 10744 17876
rect 10968 17867 11020 17876
rect 10968 17833 10977 17867
rect 10977 17833 11011 17867
rect 11011 17833 11020 17867
rect 10968 17824 11020 17833
rect 15292 17824 15344 17876
rect 19340 17824 19392 17876
rect 20076 17867 20128 17876
rect 20076 17833 20085 17867
rect 20085 17833 20119 17867
rect 20119 17833 20128 17867
rect 20076 17824 20128 17833
rect 20812 17867 20864 17876
rect 20812 17833 20821 17867
rect 20821 17833 20855 17867
rect 20855 17833 20864 17867
rect 20812 17824 20864 17833
rect 23204 17867 23256 17876
rect 23204 17833 23213 17867
rect 23213 17833 23247 17867
rect 23247 17833 23256 17867
rect 23204 17824 23256 17833
rect 24124 17867 24176 17876
rect 24124 17833 24133 17867
rect 24133 17833 24167 17867
rect 24167 17833 24176 17867
rect 24124 17824 24176 17833
rect 3608 17688 3660 17740
rect 10324 17799 10376 17808
rect 10324 17765 10333 17799
rect 10333 17765 10367 17799
rect 10367 17765 10376 17799
rect 10324 17756 10376 17765
rect 940 17620 992 17672
rect 7012 17663 7064 17672
rect 7012 17629 7021 17663
rect 7021 17629 7055 17663
rect 7055 17629 7064 17663
rect 7012 17620 7064 17629
rect 7748 17663 7800 17672
rect 4896 17552 4948 17604
rect 7748 17629 7757 17663
rect 7757 17629 7791 17663
rect 7791 17629 7800 17663
rect 7748 17620 7800 17629
rect 9220 17620 9272 17672
rect 8944 17595 8996 17604
rect 8944 17561 8953 17595
rect 8953 17561 8987 17595
rect 8987 17561 8996 17595
rect 8944 17552 8996 17561
rect 9772 17620 9824 17672
rect 9036 17484 9088 17536
rect 9312 17527 9364 17536
rect 9312 17493 9321 17527
rect 9321 17493 9355 17527
rect 9355 17493 9364 17527
rect 9312 17484 9364 17493
rect 9404 17484 9456 17536
rect 9588 17484 9640 17536
rect 10232 17552 10284 17604
rect 10784 17688 10836 17740
rect 13176 17756 13228 17808
rect 16672 17756 16724 17808
rect 20444 17756 20496 17808
rect 20996 17756 21048 17808
rect 11612 17663 11664 17672
rect 11612 17629 11621 17663
rect 11621 17629 11655 17663
rect 11655 17629 11664 17663
rect 15200 17688 15252 17740
rect 11612 17620 11664 17629
rect 10692 17484 10744 17536
rect 11336 17484 11388 17536
rect 11428 17527 11480 17536
rect 11428 17493 11437 17527
rect 11437 17493 11471 17527
rect 11471 17493 11480 17527
rect 14464 17620 14516 17672
rect 14648 17663 14700 17672
rect 14648 17629 14657 17663
rect 14657 17629 14691 17663
rect 14691 17629 14700 17663
rect 14648 17620 14700 17629
rect 14740 17620 14792 17672
rect 12532 17595 12584 17604
rect 12532 17561 12541 17595
rect 12541 17561 12575 17595
rect 12575 17561 12584 17595
rect 12532 17552 12584 17561
rect 14556 17552 14608 17604
rect 15568 17620 15620 17672
rect 15660 17620 15712 17672
rect 18052 17620 18104 17672
rect 11428 17484 11480 17493
rect 12256 17484 12308 17536
rect 12440 17484 12492 17536
rect 14832 17484 14884 17536
rect 15200 17552 15252 17604
rect 18880 17663 18932 17672
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 22008 17688 22060 17740
rect 20444 17663 20496 17672
rect 20444 17629 20453 17663
rect 20453 17629 20487 17663
rect 20487 17629 20496 17663
rect 20444 17620 20496 17629
rect 20628 17663 20680 17672
rect 20628 17629 20644 17663
rect 20644 17629 20680 17663
rect 20628 17620 20680 17629
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 20904 17620 20956 17672
rect 18052 17484 18104 17536
rect 18604 17484 18656 17536
rect 20168 17484 20220 17536
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 23296 17552 23348 17604
rect 24124 17620 24176 17672
rect 25136 17552 25188 17604
rect 21180 17484 21232 17536
rect 23112 17484 23164 17536
rect 33140 17484 33192 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4896 17280 4948 17332
rect 5448 17323 5500 17332
rect 5448 17289 5457 17323
rect 5457 17289 5491 17323
rect 5491 17289 5500 17323
rect 5448 17280 5500 17289
rect 5908 17280 5960 17332
rect 9036 17280 9088 17332
rect 4712 17144 4764 17196
rect 8944 17212 8996 17264
rect 9588 17280 9640 17332
rect 11428 17280 11480 17332
rect 13176 17280 13228 17332
rect 13452 17280 13504 17332
rect 14832 17323 14884 17332
rect 14832 17289 14841 17323
rect 14841 17289 14875 17323
rect 14875 17289 14884 17323
rect 14832 17280 14884 17289
rect 15200 17280 15252 17332
rect 8760 17187 8812 17196
rect 8760 17153 8769 17187
rect 8769 17153 8803 17187
rect 8803 17153 8812 17187
rect 8760 17144 8812 17153
rect 8852 17187 8904 17196
rect 8852 17153 8861 17187
rect 8861 17153 8895 17187
rect 8895 17153 8904 17187
rect 8852 17144 8904 17153
rect 9036 17187 9088 17196
rect 9036 17153 9045 17187
rect 9045 17153 9079 17187
rect 9079 17153 9088 17187
rect 9036 17144 9088 17153
rect 9404 17144 9456 17196
rect 12256 17255 12308 17264
rect 12256 17221 12265 17255
rect 12265 17221 12299 17255
rect 12299 17221 12308 17255
rect 12256 17212 12308 17221
rect 12532 17212 12584 17264
rect 8668 17076 8720 17128
rect 9312 17076 9364 17128
rect 9864 17187 9916 17196
rect 9864 17153 9873 17187
rect 9873 17153 9907 17187
rect 9907 17153 9916 17187
rect 9864 17144 9916 17153
rect 13084 17144 13136 17196
rect 9680 17076 9732 17128
rect 12256 17076 12308 17128
rect 12440 17076 12492 17128
rect 9220 17008 9272 17060
rect 10692 17008 10744 17060
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 8576 16983 8628 16992
rect 8576 16949 8622 16983
rect 8622 16949 8628 16983
rect 8576 16940 8628 16949
rect 10600 16940 10652 16992
rect 13268 17076 13320 17128
rect 14924 17144 14976 17196
rect 15108 17144 15160 17196
rect 18880 17212 18932 17264
rect 22008 17323 22060 17332
rect 22008 17289 22017 17323
rect 22017 17289 22051 17323
rect 22051 17289 22060 17323
rect 22008 17280 22060 17289
rect 23296 17280 23348 17332
rect 25136 17280 25188 17332
rect 17960 17187 18012 17196
rect 17960 17153 17969 17187
rect 17969 17153 18003 17187
rect 18003 17153 18012 17187
rect 17960 17144 18012 17153
rect 18604 17187 18656 17196
rect 18604 17153 18613 17187
rect 18613 17153 18647 17187
rect 18647 17153 18656 17187
rect 18604 17144 18656 17153
rect 18052 17119 18104 17128
rect 18052 17085 18061 17119
rect 18061 17085 18095 17119
rect 18095 17085 18104 17119
rect 18052 17076 18104 17085
rect 14556 17051 14608 17060
rect 14556 17017 14565 17051
rect 14565 17017 14599 17051
rect 14599 17017 14608 17051
rect 14556 17008 14608 17017
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 20904 17144 20956 17196
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 21180 17212 21232 17264
rect 25412 17280 25464 17332
rect 20628 17076 20680 17128
rect 13452 16940 13504 16992
rect 13728 16983 13780 16992
rect 13728 16949 13737 16983
rect 13737 16949 13771 16983
rect 13771 16949 13780 16983
rect 13728 16940 13780 16949
rect 15660 16940 15712 16992
rect 19340 16940 19392 16992
rect 21180 16940 21232 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 8760 16736 8812 16788
rect 8484 16668 8536 16720
rect 10232 16736 10284 16788
rect 10784 16736 10836 16788
rect 12716 16736 12768 16788
rect 12808 16736 12860 16788
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 13728 16779 13780 16788
rect 13728 16745 13737 16779
rect 13737 16745 13771 16779
rect 13771 16745 13780 16779
rect 13728 16736 13780 16745
rect 3608 16600 3660 16652
rect 4620 16600 4672 16652
rect 8576 16600 8628 16652
rect 9496 16600 9548 16652
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 6828 16575 6880 16584
rect 6828 16541 6837 16575
rect 6837 16541 6871 16575
rect 6871 16541 6880 16575
rect 6828 16532 6880 16541
rect 9956 16643 10008 16652
rect 9956 16609 9965 16643
rect 9965 16609 9999 16643
rect 9999 16609 10008 16643
rect 9956 16600 10008 16609
rect 10232 16600 10284 16652
rect 4620 16464 4672 16516
rect 8944 16464 8996 16516
rect 9496 16464 9548 16516
rect 10324 16507 10376 16516
rect 10324 16473 10351 16507
rect 10351 16473 10376 16507
rect 10324 16464 10376 16473
rect 9404 16396 9456 16448
rect 10508 16507 10560 16516
rect 10508 16473 10517 16507
rect 10517 16473 10551 16507
rect 10551 16473 10560 16507
rect 10508 16464 10560 16473
rect 12256 16532 12308 16584
rect 14648 16736 14700 16788
rect 15660 16779 15712 16788
rect 15660 16745 15669 16779
rect 15669 16745 15703 16779
rect 15703 16745 15712 16779
rect 15660 16736 15712 16745
rect 20812 16736 20864 16788
rect 21180 16779 21232 16788
rect 21180 16745 21189 16779
rect 21189 16745 21223 16779
rect 21223 16745 21232 16779
rect 21180 16736 21232 16745
rect 15476 16668 15528 16720
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 12624 16575 12676 16584
rect 12624 16541 12633 16575
rect 12633 16541 12667 16575
rect 12667 16541 12676 16575
rect 12624 16532 12676 16541
rect 12900 16532 12952 16584
rect 13360 16532 13412 16584
rect 13728 16532 13780 16584
rect 12532 16464 12584 16516
rect 13176 16464 13228 16516
rect 10784 16396 10836 16448
rect 13360 16396 13412 16448
rect 14188 16532 14240 16584
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 14832 16532 14884 16584
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15108 16532 15160 16541
rect 16396 16600 16448 16652
rect 19248 16668 19300 16720
rect 15476 16464 15528 16516
rect 16304 16532 16356 16584
rect 19340 16600 19392 16652
rect 18788 16575 18840 16584
rect 18788 16541 18797 16575
rect 18797 16541 18831 16575
rect 18831 16541 18840 16575
rect 18788 16532 18840 16541
rect 19432 16532 19484 16584
rect 20628 16532 20680 16584
rect 14648 16439 14700 16448
rect 14648 16405 14657 16439
rect 14657 16405 14691 16439
rect 14691 16405 14700 16439
rect 14648 16396 14700 16405
rect 20168 16464 20220 16516
rect 20904 16532 20956 16584
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 33140 16575 33192 16584
rect 33140 16541 33149 16575
rect 33149 16541 33183 16575
rect 33183 16541 33192 16575
rect 33140 16532 33192 16541
rect 21272 16464 21324 16516
rect 34888 16464 34940 16516
rect 19984 16396 20036 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4620 16192 4672 16244
rect 4712 16192 4764 16244
rect 6368 16192 6420 16244
rect 5264 16099 5316 16108
rect 5264 16065 5273 16099
rect 5273 16065 5307 16099
rect 5307 16065 5316 16099
rect 5264 16056 5316 16065
rect 6460 16056 6512 16108
rect 6828 16099 6880 16108
rect 6828 16065 6837 16099
rect 6837 16065 6871 16099
rect 6871 16065 6880 16099
rect 6828 16056 6880 16065
rect 8484 16124 8536 16176
rect 8576 16167 8628 16176
rect 8576 16133 8585 16167
rect 8585 16133 8619 16167
rect 8619 16133 8628 16167
rect 8576 16124 8628 16133
rect 9036 16124 9088 16176
rect 9496 16124 9548 16176
rect 11244 16056 11296 16108
rect 7932 15988 7984 16040
rect 8392 15988 8444 16040
rect 6552 15920 6604 15972
rect 6644 15920 6696 15972
rect 10048 15988 10100 16040
rect 10416 15988 10468 16040
rect 12164 16056 12216 16108
rect 12716 16056 12768 16108
rect 12992 16056 13044 16108
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 14832 16192 14884 16244
rect 15384 16192 15436 16244
rect 16580 16192 16632 16244
rect 18788 16192 18840 16244
rect 19984 16192 20036 16244
rect 20260 16192 20312 16244
rect 19248 16124 19300 16176
rect 21088 16192 21140 16244
rect 12256 16031 12308 16040
rect 12256 15997 12265 16031
rect 12265 15997 12299 16031
rect 12299 15997 12308 16031
rect 12256 15988 12308 15997
rect 20076 16099 20128 16108
rect 20076 16065 20085 16099
rect 20085 16065 20119 16099
rect 20119 16065 20128 16099
rect 20076 16056 20128 16065
rect 20260 16056 20312 16108
rect 20444 16099 20496 16108
rect 20444 16065 20453 16099
rect 20453 16065 20487 16099
rect 20487 16065 20496 16099
rect 20444 16056 20496 16065
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 23112 16235 23164 16244
rect 23112 16201 23121 16235
rect 23121 16201 23155 16235
rect 23155 16201 23164 16235
rect 23112 16192 23164 16201
rect 23296 16192 23348 16244
rect 33140 16192 33192 16244
rect 22008 16099 22060 16108
rect 22008 16065 22017 16099
rect 22017 16065 22051 16099
rect 22051 16065 22060 16099
rect 22008 16056 22060 16065
rect 22468 16099 22520 16108
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 22836 16056 22888 16108
rect 25412 16056 25464 16108
rect 26056 16056 26108 16108
rect 10232 15963 10284 15972
rect 10232 15929 10241 15963
rect 10241 15929 10275 15963
rect 10275 15929 10284 15963
rect 10232 15920 10284 15929
rect 12992 15963 13044 15972
rect 12992 15929 13001 15963
rect 13001 15929 13035 15963
rect 13035 15929 13044 15963
rect 12992 15920 13044 15929
rect 6736 15852 6788 15904
rect 9956 15852 10008 15904
rect 11612 15852 11664 15904
rect 12072 15895 12124 15904
rect 12072 15861 12081 15895
rect 12081 15861 12115 15895
rect 12115 15861 12124 15895
rect 12072 15852 12124 15861
rect 12348 15852 12400 15904
rect 13268 15895 13320 15904
rect 13268 15861 13277 15895
rect 13277 15861 13311 15895
rect 13311 15861 13320 15895
rect 13268 15852 13320 15861
rect 16488 15920 16540 15972
rect 20904 15920 20956 15972
rect 24124 15988 24176 16040
rect 15660 15852 15712 15904
rect 16304 15852 16356 15904
rect 16764 15895 16816 15904
rect 16764 15861 16773 15895
rect 16773 15861 16807 15895
rect 16807 15861 16816 15895
rect 16764 15852 16816 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 6184 15691 6236 15700
rect 6184 15657 6193 15691
rect 6193 15657 6227 15691
rect 6227 15657 6236 15691
rect 6184 15648 6236 15657
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 4344 15308 4396 15360
rect 6828 15648 6880 15700
rect 7196 15648 7248 15700
rect 8852 15648 8904 15700
rect 10324 15648 10376 15700
rect 11612 15648 11664 15700
rect 13176 15648 13228 15700
rect 15292 15691 15344 15700
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 6460 15580 6512 15632
rect 6644 15623 6696 15632
rect 6644 15589 6653 15623
rect 6653 15589 6687 15623
rect 6687 15589 6696 15623
rect 6644 15580 6696 15589
rect 6920 15580 6972 15632
rect 6552 15487 6604 15496
rect 6552 15453 6558 15487
rect 6558 15453 6604 15487
rect 6552 15444 6604 15453
rect 10692 15580 10744 15632
rect 12072 15580 12124 15632
rect 12716 15580 12768 15632
rect 12992 15580 13044 15632
rect 13360 15580 13412 15632
rect 16580 15648 16632 15700
rect 16764 15648 16816 15700
rect 22008 15648 22060 15700
rect 22468 15648 22520 15700
rect 24124 15648 24176 15700
rect 16396 15580 16448 15632
rect 16488 15580 16540 15632
rect 7288 15444 7340 15496
rect 7932 15487 7984 15496
rect 7196 15376 7248 15428
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 8208 15487 8260 15496
rect 8208 15453 8217 15487
rect 8217 15453 8251 15487
rect 8251 15453 8260 15487
rect 8208 15444 8260 15453
rect 8392 15444 8444 15496
rect 10232 15512 10284 15564
rect 9680 15487 9732 15496
rect 9680 15453 9689 15487
rect 9689 15453 9723 15487
rect 9723 15453 9732 15487
rect 9680 15444 9732 15453
rect 9772 15487 9824 15496
rect 9772 15453 9781 15487
rect 9781 15453 9815 15487
rect 9815 15453 9824 15487
rect 9772 15444 9824 15453
rect 10048 15444 10100 15496
rect 10416 15487 10468 15496
rect 10416 15453 10425 15487
rect 10425 15453 10459 15487
rect 10459 15453 10468 15487
rect 10416 15444 10468 15453
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 10784 15444 10836 15453
rect 11244 15444 11296 15496
rect 13268 15512 13320 15564
rect 10784 15308 10836 15360
rect 12348 15444 12400 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 12992 15444 13044 15496
rect 13820 15512 13872 15564
rect 15108 15512 15160 15564
rect 13544 15444 13596 15496
rect 13728 15376 13780 15428
rect 15384 15487 15436 15496
rect 15384 15453 15393 15487
rect 15393 15453 15427 15487
rect 15427 15453 15436 15487
rect 15384 15444 15436 15453
rect 15660 15487 15712 15496
rect 15660 15453 15669 15487
rect 15669 15453 15703 15487
rect 15703 15453 15712 15487
rect 15660 15444 15712 15453
rect 20444 15512 20496 15564
rect 20720 15512 20772 15564
rect 20536 15444 20588 15496
rect 12808 15308 12860 15360
rect 13084 15308 13136 15360
rect 16580 15308 16632 15360
rect 16764 15351 16816 15360
rect 16764 15317 16773 15351
rect 16773 15317 16807 15351
rect 16807 15317 16816 15351
rect 16764 15308 16816 15317
rect 19984 15308 20036 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 6736 15104 6788 15156
rect 9496 15104 9548 15156
rect 4344 15079 4396 15088
rect 4344 15045 4353 15079
rect 4353 15045 4387 15079
rect 4387 15045 4396 15079
rect 4344 15036 4396 15045
rect 5080 15036 5132 15088
rect 3608 14968 3660 15020
rect 4068 15011 4120 15020
rect 4068 14977 4077 15011
rect 4077 14977 4111 15011
rect 4111 14977 4120 15011
rect 4068 14968 4120 14977
rect 6920 15036 6972 15088
rect 8944 15036 8996 15088
rect 9680 15079 9732 15088
rect 9680 15045 9689 15079
rect 9689 15045 9723 15079
rect 9723 15045 9732 15079
rect 9680 15036 9732 15045
rect 9772 15036 9824 15088
rect 10416 15079 10468 15088
rect 10416 15045 10425 15079
rect 10425 15045 10459 15079
rect 10459 15045 10468 15079
rect 10416 15036 10468 15045
rect 12532 15104 12584 15156
rect 13820 15104 13872 15156
rect 16580 15104 16632 15156
rect 16672 15104 16724 15156
rect 19340 15104 19392 15156
rect 19432 15104 19484 15156
rect 11244 15079 11296 15088
rect 11244 15045 11253 15079
rect 11253 15045 11287 15079
rect 11287 15045 11296 15079
rect 11244 15036 11296 15045
rect 7196 14968 7248 15020
rect 7656 14943 7708 14952
rect 6828 14832 6880 14884
rect 6552 14764 6604 14816
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 7472 14832 7524 14884
rect 8668 14968 8720 15020
rect 10692 14968 10744 15020
rect 8208 14900 8260 14952
rect 9772 14900 9824 14952
rect 10968 14968 11020 15020
rect 12164 14968 12216 15020
rect 12716 14968 12768 15020
rect 14924 14968 14976 15020
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 19248 15036 19300 15088
rect 13452 14900 13504 14952
rect 15292 14900 15344 14952
rect 16764 14900 16816 14952
rect 18052 14900 18104 14952
rect 18972 14943 19024 14952
rect 18972 14909 18981 14943
rect 18981 14909 19015 14943
rect 19015 14909 19024 14943
rect 18972 14900 19024 14909
rect 20076 14900 20128 14952
rect 10876 14832 10928 14884
rect 11428 14832 11480 14884
rect 11980 14832 12032 14884
rect 12900 14832 12952 14884
rect 20352 14832 20404 14884
rect 20996 14832 21048 14884
rect 10600 14764 10652 14816
rect 13544 14764 13596 14816
rect 15660 14764 15712 14816
rect 18236 14807 18288 14816
rect 18236 14773 18245 14807
rect 18245 14773 18279 14807
rect 18279 14773 18288 14807
rect 18236 14764 18288 14773
rect 19340 14764 19392 14816
rect 20444 14764 20496 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 4712 14560 4764 14612
rect 5080 14560 5132 14612
rect 5264 14560 5316 14612
rect 6092 14560 6144 14612
rect 6828 14603 6880 14612
rect 6828 14569 6837 14603
rect 6837 14569 6871 14603
rect 6871 14569 6880 14603
rect 6828 14560 6880 14569
rect 10048 14603 10100 14612
rect 10048 14569 10057 14603
rect 10057 14569 10091 14603
rect 10091 14569 10100 14603
rect 10048 14560 10100 14569
rect 10968 14560 11020 14612
rect 11796 14560 11848 14612
rect 12348 14560 12400 14612
rect 13084 14560 13136 14612
rect 14556 14560 14608 14612
rect 18052 14560 18104 14612
rect 18236 14560 18288 14612
rect 19340 14560 19392 14612
rect 19984 14603 20036 14612
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 5908 14492 5960 14544
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 6736 14356 6788 14408
rect 7196 14356 7248 14408
rect 8484 14356 8536 14408
rect 10232 14356 10284 14408
rect 7840 14288 7892 14340
rect 10140 14288 10192 14340
rect 10968 14356 11020 14408
rect 11060 14356 11112 14408
rect 11244 14356 11296 14408
rect 12072 14467 12124 14476
rect 12072 14433 12081 14467
rect 12081 14433 12115 14467
rect 12115 14433 12124 14467
rect 12072 14424 12124 14433
rect 14464 14492 14516 14544
rect 10692 14331 10744 14340
rect 10692 14297 10701 14331
rect 10701 14297 10735 14331
rect 10735 14297 10744 14331
rect 10692 14288 10744 14297
rect 10784 14331 10836 14340
rect 10784 14297 10793 14331
rect 10793 14297 10827 14331
rect 10827 14297 10836 14331
rect 10784 14288 10836 14297
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 11704 14356 11756 14408
rect 11980 14399 12032 14408
rect 11980 14365 11989 14399
rect 11989 14365 12023 14399
rect 12023 14365 12032 14399
rect 11980 14356 12032 14365
rect 12164 14356 12216 14408
rect 12348 14399 12400 14408
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 12716 14424 12768 14476
rect 13452 14467 13504 14476
rect 13452 14433 13461 14467
rect 13461 14433 13495 14467
rect 13495 14433 13504 14467
rect 13452 14424 13504 14433
rect 13544 14424 13596 14476
rect 12532 14356 12584 14408
rect 12900 14356 12952 14408
rect 13636 14399 13688 14408
rect 13636 14365 13645 14399
rect 13645 14365 13679 14399
rect 13679 14365 13688 14399
rect 13636 14356 13688 14365
rect 13728 14356 13780 14408
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 16396 14492 16448 14544
rect 15292 14399 15344 14408
rect 5448 14263 5500 14272
rect 5448 14229 5457 14263
rect 5457 14229 5491 14263
rect 5491 14229 5500 14263
rect 5448 14220 5500 14229
rect 11520 14220 11572 14272
rect 12256 14220 12308 14272
rect 12808 14288 12860 14340
rect 13360 14331 13412 14340
rect 13360 14297 13369 14331
rect 13369 14297 13403 14331
rect 13403 14297 13412 14331
rect 13360 14288 13412 14297
rect 13820 14288 13872 14340
rect 12532 14263 12584 14272
rect 12532 14229 12541 14263
rect 12541 14229 12575 14263
rect 12575 14229 12584 14263
rect 12532 14220 12584 14229
rect 13176 14263 13228 14272
rect 13176 14229 13185 14263
rect 13185 14229 13219 14263
rect 13219 14229 13228 14263
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16120 14356 16172 14408
rect 20720 14535 20772 14544
rect 20720 14501 20729 14535
rect 20729 14501 20763 14535
rect 20763 14501 20772 14535
rect 20720 14492 20772 14501
rect 19432 14424 19484 14476
rect 20812 14424 20864 14476
rect 19340 14356 19392 14408
rect 18788 14288 18840 14340
rect 20260 14356 20312 14408
rect 20352 14356 20404 14408
rect 20996 14399 21048 14408
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 22468 14560 22520 14612
rect 22836 14560 22888 14612
rect 22560 14424 22612 14476
rect 13176 14220 13228 14229
rect 15752 14263 15804 14272
rect 15752 14229 15761 14263
rect 15761 14229 15795 14263
rect 15795 14229 15804 14263
rect 15752 14220 15804 14229
rect 17040 14220 17092 14272
rect 18880 14220 18932 14272
rect 19984 14220 20036 14272
rect 20812 14331 20864 14340
rect 20812 14297 20840 14331
rect 20840 14297 20864 14331
rect 20812 14288 20864 14297
rect 20720 14220 20772 14272
rect 22468 14399 22520 14408
rect 22468 14365 22477 14399
rect 22477 14365 22511 14399
rect 22511 14365 22520 14399
rect 22468 14356 22520 14365
rect 33140 14399 33192 14408
rect 33140 14365 33149 14399
rect 33149 14365 33183 14399
rect 33183 14365 33192 14399
rect 33140 14356 33192 14365
rect 34888 14288 34940 14340
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 5908 14016 5960 14068
rect 6368 14016 6420 14068
rect 8944 14016 8996 14068
rect 10140 14016 10192 14068
rect 6092 13991 6144 14000
rect 6092 13957 6101 13991
rect 6101 13957 6135 13991
rect 6135 13957 6144 13991
rect 6092 13948 6144 13957
rect 4068 13923 4120 13932
rect 4068 13889 4077 13923
rect 4077 13889 4111 13923
rect 4111 13889 4120 13923
rect 4068 13880 4120 13889
rect 5448 13880 5500 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 7656 13880 7708 13932
rect 8668 13787 8720 13796
rect 8668 13753 8677 13787
rect 8677 13753 8711 13787
rect 8711 13753 8720 13787
rect 8668 13744 8720 13753
rect 10232 13880 10284 13932
rect 12256 14016 12308 14068
rect 13452 14016 13504 14068
rect 13084 13948 13136 14000
rect 11060 13923 11112 13932
rect 11060 13889 11069 13923
rect 11069 13889 11103 13923
rect 11103 13889 11112 13923
rect 11060 13880 11112 13889
rect 13176 13923 13228 13932
rect 13176 13889 13185 13923
rect 13185 13889 13219 13923
rect 13219 13889 13228 13923
rect 13176 13880 13228 13889
rect 13452 13923 13504 13932
rect 13452 13889 13461 13923
rect 13461 13889 13495 13923
rect 13495 13889 13504 13923
rect 13452 13880 13504 13889
rect 14556 13991 14608 14000
rect 14556 13957 14565 13991
rect 14565 13957 14599 13991
rect 14599 13957 14608 13991
rect 14556 13948 14608 13957
rect 15292 14016 15344 14068
rect 15752 14016 15804 14068
rect 18880 14059 18932 14068
rect 18880 14025 18889 14059
rect 18889 14025 18923 14059
rect 18923 14025 18932 14059
rect 18880 14016 18932 14025
rect 18972 14016 19024 14068
rect 20260 14059 20312 14068
rect 20260 14025 20269 14059
rect 20269 14025 20303 14059
rect 20303 14025 20312 14059
rect 20260 14016 20312 14025
rect 20444 14016 20496 14068
rect 13728 13880 13780 13932
rect 14096 13880 14148 13932
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 14372 13923 14424 13932
rect 14372 13889 14381 13923
rect 14381 13889 14415 13923
rect 14415 13889 14424 13923
rect 14372 13880 14424 13889
rect 11704 13744 11756 13796
rect 12716 13744 12768 13796
rect 13360 13744 13412 13796
rect 4712 13676 4764 13728
rect 10692 13719 10744 13728
rect 10692 13685 10701 13719
rect 10701 13685 10735 13719
rect 10735 13685 10744 13719
rect 10692 13676 10744 13685
rect 11980 13676 12032 13728
rect 12348 13719 12400 13728
rect 12348 13685 12357 13719
rect 12357 13685 12391 13719
rect 12391 13685 12400 13719
rect 12348 13676 12400 13685
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 13912 13719 13964 13728
rect 13912 13685 13921 13719
rect 13921 13685 13955 13719
rect 13955 13685 13964 13719
rect 13912 13676 13964 13685
rect 14096 13744 14148 13796
rect 15108 13880 15160 13932
rect 15660 13923 15712 13932
rect 15660 13889 15669 13923
rect 15669 13889 15703 13923
rect 15703 13889 15712 13923
rect 15660 13880 15712 13889
rect 17960 13880 18012 13932
rect 18052 13812 18104 13864
rect 18880 13880 18932 13932
rect 19248 13948 19300 14000
rect 19616 13880 19668 13932
rect 21272 14016 21324 14068
rect 22468 14016 22520 14068
rect 24124 14016 24176 14068
rect 33140 14016 33192 14068
rect 19432 13812 19484 13864
rect 14924 13719 14976 13728
rect 14924 13685 14933 13719
rect 14933 13685 14967 13719
rect 14967 13685 14976 13719
rect 14924 13676 14976 13685
rect 16304 13676 16356 13728
rect 19340 13676 19392 13728
rect 21732 13744 21784 13796
rect 22560 13880 22612 13932
rect 26056 13991 26108 14000
rect 26056 13957 26065 13991
rect 26065 13957 26099 13991
rect 26099 13957 26108 13991
rect 26056 13948 26108 13957
rect 23480 13812 23532 13864
rect 24124 13812 24176 13864
rect 25044 13812 25096 13864
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 6368 13515 6420 13524
rect 6368 13481 6377 13515
rect 6377 13481 6411 13515
rect 6411 13481 6420 13515
rect 6368 13472 6420 13481
rect 8392 13515 8444 13524
rect 8392 13481 8401 13515
rect 8401 13481 8435 13515
rect 8435 13481 8444 13515
rect 8392 13472 8444 13481
rect 12072 13472 12124 13524
rect 12624 13472 12676 13524
rect 12716 13515 12768 13524
rect 12716 13481 12725 13515
rect 12725 13481 12759 13515
rect 12759 13481 12768 13515
rect 12716 13472 12768 13481
rect 12808 13472 12860 13524
rect 17960 13472 18012 13524
rect 19340 13472 19392 13524
rect 19432 13472 19484 13524
rect 4068 13379 4120 13388
rect 4068 13345 4077 13379
rect 4077 13345 4111 13379
rect 4111 13345 4120 13379
rect 4068 13336 4120 13345
rect 12348 13404 12400 13456
rect 13728 13404 13780 13456
rect 11796 13336 11848 13388
rect 940 13268 992 13320
rect 7104 13268 7156 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 7840 13268 7892 13320
rect 10692 13268 10744 13320
rect 11980 13311 12032 13320
rect 11980 13277 11989 13311
rect 11989 13277 12023 13311
rect 12023 13277 12032 13311
rect 11980 13268 12032 13277
rect 5080 13200 5132 13252
rect 11704 13200 11756 13252
rect 12624 13336 12676 13388
rect 12808 13336 12860 13388
rect 12992 13268 13044 13320
rect 14096 13311 14148 13320
rect 14096 13277 14105 13311
rect 14105 13277 14139 13311
rect 14139 13277 14148 13311
rect 14096 13268 14148 13277
rect 18880 13404 18932 13456
rect 17040 13268 17092 13320
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 11520 13132 11572 13184
rect 13544 13132 13596 13184
rect 19984 13515 20036 13524
rect 19984 13481 19993 13515
rect 19993 13481 20027 13515
rect 20027 13481 20036 13515
rect 19984 13472 20036 13481
rect 22560 13472 22612 13524
rect 22652 13515 22704 13524
rect 22652 13481 22661 13515
rect 22661 13481 22695 13515
rect 22695 13481 22704 13515
rect 22652 13472 22704 13481
rect 19616 13268 19668 13320
rect 21456 13268 21508 13320
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 22192 13311 22244 13320
rect 22192 13277 22201 13311
rect 22201 13277 22235 13311
rect 22235 13277 22244 13311
rect 22192 13268 22244 13277
rect 22468 13200 22520 13252
rect 14004 13132 14056 13184
rect 16028 13132 16080 13184
rect 17868 13132 17920 13184
rect 18604 13132 18656 13184
rect 22100 13132 22152 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 5080 12928 5132 12980
rect 5540 12971 5592 12980
rect 5540 12937 5549 12971
rect 5549 12937 5583 12971
rect 5583 12937 5592 12971
rect 5540 12928 5592 12937
rect 10784 12860 10836 12912
rect 7288 12835 7340 12844
rect 7288 12801 7297 12835
rect 7297 12801 7331 12835
rect 7331 12801 7340 12835
rect 7288 12792 7340 12801
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 10232 12835 10284 12844
rect 10232 12801 10241 12835
rect 10241 12801 10275 12835
rect 10275 12801 10284 12835
rect 10232 12792 10284 12801
rect 10048 12699 10100 12708
rect 10048 12665 10057 12699
rect 10057 12665 10091 12699
rect 10091 12665 10100 12699
rect 10048 12656 10100 12665
rect 10876 12767 10928 12776
rect 10876 12733 10885 12767
rect 10885 12733 10919 12767
rect 10919 12733 10928 12767
rect 10876 12724 10928 12733
rect 11980 12928 12032 12980
rect 12900 12928 12952 12980
rect 11244 12792 11296 12844
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 12808 12860 12860 12912
rect 14004 12928 14056 12980
rect 14096 12928 14148 12980
rect 11336 12724 11388 12776
rect 13912 12792 13964 12844
rect 14924 12928 14976 12980
rect 16028 12903 16080 12912
rect 16028 12869 16037 12903
rect 16037 12869 16071 12903
rect 16071 12869 16080 12903
rect 16028 12860 16080 12869
rect 14372 12792 14424 12844
rect 14556 12835 14608 12844
rect 14556 12801 14565 12835
rect 14565 12801 14599 12835
rect 14599 12801 14608 12835
rect 14556 12792 14608 12801
rect 14924 12792 14976 12844
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 17040 12928 17092 12980
rect 18052 12928 18104 12980
rect 17132 12903 17184 12912
rect 17132 12869 17141 12903
rect 17141 12869 17175 12903
rect 17175 12869 17184 12903
rect 17132 12860 17184 12869
rect 16580 12724 16632 12776
rect 16948 12835 17000 12844
rect 16948 12801 16957 12835
rect 16957 12801 16991 12835
rect 16991 12801 17000 12835
rect 16948 12792 17000 12801
rect 17040 12792 17092 12844
rect 17500 12792 17552 12844
rect 16120 12699 16172 12708
rect 16120 12665 16129 12699
rect 16129 12665 16163 12699
rect 16163 12665 16172 12699
rect 16120 12656 16172 12665
rect 17868 12724 17920 12776
rect 17960 12724 18012 12776
rect 22468 12792 22520 12844
rect 18604 12767 18656 12776
rect 18604 12733 18613 12767
rect 18613 12733 18647 12767
rect 18647 12733 18656 12767
rect 18604 12724 18656 12733
rect 22100 12724 22152 12776
rect 12164 12588 12216 12640
rect 12440 12588 12492 12640
rect 13544 12588 13596 12640
rect 13728 12588 13780 12640
rect 15752 12631 15804 12640
rect 15752 12597 15761 12631
rect 15761 12597 15795 12631
rect 15795 12597 15804 12631
rect 15752 12588 15804 12597
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 23572 12588 23624 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 6184 12384 6236 12436
rect 10876 12384 10928 12436
rect 11888 12384 11940 12436
rect 12164 12384 12216 12436
rect 3884 12248 3936 12300
rect 14924 12384 14976 12436
rect 16580 12384 16632 12436
rect 17040 12427 17092 12436
rect 17040 12393 17049 12427
rect 17049 12393 17083 12427
rect 17083 12393 17092 12427
rect 17040 12384 17092 12393
rect 17868 12427 17920 12436
rect 17868 12393 17877 12427
rect 17877 12393 17911 12427
rect 17911 12393 17920 12427
rect 17868 12384 17920 12393
rect 22468 12427 22520 12436
rect 22468 12393 22477 12427
rect 22477 12393 22511 12427
rect 22511 12393 22520 12427
rect 22468 12384 22520 12393
rect 10048 12180 10100 12232
rect 4712 12112 4764 12164
rect 5172 12112 5224 12164
rect 7196 12112 7248 12164
rect 10232 12112 10284 12164
rect 10968 12180 11020 12232
rect 11336 12180 11388 12232
rect 11520 12180 11572 12232
rect 11888 12180 11940 12232
rect 12532 12223 12584 12232
rect 12532 12189 12541 12223
rect 12541 12189 12575 12223
rect 12575 12189 12584 12223
rect 12532 12180 12584 12189
rect 13728 12248 13780 12300
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 14188 12180 14240 12232
rect 14372 12180 14424 12232
rect 21640 12316 21692 12368
rect 17132 12180 17184 12232
rect 17500 12223 17552 12232
rect 17500 12189 17509 12223
rect 17509 12189 17543 12223
rect 17543 12189 17552 12223
rect 17500 12180 17552 12189
rect 22192 12291 22244 12300
rect 22192 12257 22201 12291
rect 22201 12257 22235 12291
rect 22235 12257 22244 12291
rect 22192 12248 22244 12257
rect 16764 12112 16816 12164
rect 16856 12112 16908 12164
rect 16948 12112 17000 12164
rect 33140 12223 33192 12232
rect 33140 12189 33149 12223
rect 33149 12189 33183 12223
rect 33183 12189 33192 12223
rect 33140 12180 33192 12189
rect 34888 12112 34940 12164
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 15660 12044 15712 12096
rect 16120 12044 16172 12096
rect 17500 12044 17552 12096
rect 20720 12044 20772 12096
rect 21824 12087 21876 12096
rect 21824 12053 21833 12087
rect 21833 12053 21867 12087
rect 21867 12053 21876 12087
rect 21824 12044 21876 12053
rect 22008 12044 22060 12096
rect 24400 12044 24452 12096
rect 24952 12087 25004 12096
rect 24952 12053 24961 12087
rect 24961 12053 24995 12087
rect 24995 12053 25004 12087
rect 24952 12044 25004 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 5172 11840 5224 11892
rect 5540 11840 5592 11892
rect 11612 11840 11664 11892
rect 11888 11840 11940 11892
rect 12164 11840 12216 11892
rect 12440 11840 12492 11892
rect 15660 11883 15712 11892
rect 15660 11849 15669 11883
rect 15669 11849 15703 11883
rect 15703 11849 15712 11883
rect 15660 11840 15712 11849
rect 15752 11840 15804 11892
rect 16120 11840 16172 11892
rect 16764 11840 16816 11892
rect 14188 11772 14240 11824
rect 11888 11679 11940 11688
rect 11888 11645 11897 11679
rect 11897 11645 11931 11679
rect 11931 11645 11940 11679
rect 11888 11636 11940 11645
rect 14372 11704 14424 11756
rect 16856 11772 16908 11824
rect 23572 11772 23624 11824
rect 24400 11772 24452 11824
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 16672 11704 16724 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 22008 11679 22060 11688
rect 22008 11645 22017 11679
rect 22017 11645 22051 11679
rect 22051 11645 22060 11679
rect 22008 11636 22060 11645
rect 21824 11568 21876 11620
rect 23296 11636 23348 11688
rect 12624 11543 12676 11552
rect 12624 11509 12633 11543
rect 12633 11509 12667 11543
rect 12667 11509 12676 11543
rect 12624 11500 12676 11509
rect 14464 11500 14516 11552
rect 20720 11500 20772 11552
rect 23296 11543 23348 11552
rect 23296 11509 23305 11543
rect 23305 11509 23339 11543
rect 23339 11509 23348 11543
rect 23296 11500 23348 11509
rect 23480 11500 23532 11552
rect 33140 11840 33192 11892
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 6184 11296 6236 11348
rect 12164 11296 12216 11348
rect 12624 11296 12676 11348
rect 7288 11160 7340 11212
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 3884 11092 3936 11144
rect 5540 11024 5592 11076
rect 12348 11024 12400 11076
rect 20720 11024 20772 11076
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 23388 10956 23440 11008
rect 24952 11135 25004 11144
rect 24952 11101 24961 11135
rect 24961 11101 24995 11135
rect 24995 11101 25004 11135
rect 24952 11092 25004 11101
rect 24860 11024 24912 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 5540 10752 5592 10804
rect 5632 10795 5684 10804
rect 5632 10761 5641 10795
rect 5641 10761 5675 10795
rect 5675 10761 5684 10795
rect 5632 10752 5684 10761
rect 12624 10684 12676 10736
rect 14464 10684 14516 10736
rect 23480 10684 23532 10736
rect 24860 10616 24912 10668
rect 9956 10412 10008 10464
rect 23296 10548 23348 10600
rect 15200 10455 15252 10464
rect 15200 10421 15209 10455
rect 15209 10421 15243 10455
rect 15243 10421 15252 10455
rect 15200 10412 15252 10421
rect 21364 10412 21416 10464
rect 33140 10412 33192 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 5632 10208 5684 10260
rect 14464 10251 14516 10260
rect 14464 10217 14473 10251
rect 14473 10217 14507 10251
rect 14507 10217 14516 10251
rect 14464 10208 14516 10217
rect 15200 10208 15252 10260
rect 32956 10208 33008 10260
rect 23388 10004 23440 10056
rect 33140 10047 33192 10056
rect 33140 10013 33149 10047
rect 33149 10013 33183 10047
rect 33183 10013 33192 10047
rect 33140 10004 33192 10013
rect 34336 9979 34388 9988
rect 34336 9945 34345 9979
rect 34345 9945 34379 9979
rect 34379 9945 34388 9979
rect 34336 9936 34388 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 4804 9120 4856 9172
rect 6184 9120 6236 9172
rect 940 8916 992 8968
rect 4528 8848 4580 8900
rect 4988 8848 5040 8900
rect 10048 8848 10100 8900
rect 9956 8780 10008 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4988 8576 5040 8628
rect 5632 8576 5684 8628
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 32956 8075 33008 8084
rect 32956 8041 32965 8075
rect 32965 8041 32999 8075
rect 32999 8041 33008 8075
rect 32956 8032 33008 8041
rect 34888 7760 34940 7812
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 940 6740 992 6792
rect 4896 6604 4948 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 21640 5763 21692 5772
rect 21640 5729 21649 5763
rect 21649 5729 21683 5763
rect 21683 5729 21692 5763
rect 21640 5720 21692 5729
rect 21364 5695 21416 5704
rect 20812 5516 20864 5568
rect 21364 5661 21373 5695
rect 21373 5661 21407 5695
rect 21407 5661 21416 5695
rect 21364 5652 21416 5661
rect 23204 5652 23256 5704
rect 34336 5627 34388 5636
rect 34336 5593 34345 5627
rect 34345 5593 34379 5627
rect 34379 5593 34388 5627
rect 34336 5584 34388 5593
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 4620 4768 4672 4820
rect 940 4564 992 4616
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 20720 3680 20772 3732
rect 20812 3519 20864 3528
rect 9956 3340 10008 3392
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 23204 3476 23256 3528
rect 34888 3408 34940 3460
rect 23204 3383 23256 3392
rect 23204 3349 23213 3383
rect 23213 3349 23247 3383
rect 23247 3349 23256 3383
rect 23204 3340 23256 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 20720 3179 20772 3188
rect 20720 3145 20729 3179
rect 20729 3145 20763 3179
rect 20763 3145 20772 3179
rect 20720 3136 20772 3145
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4712 2592 4764 2644
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 9956 2456 10008 2465
rect 23204 2456 23256 2508
rect 940 2388 992 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 27344 2431 27396 2440
rect 27344 2397 27353 2431
rect 27353 2397 27387 2431
rect 27387 2397 27396 2431
rect 27344 2388 27396 2397
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 952 36174 980 36751
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 940 36168 992 36174
rect 940 36110 992 36116
rect 25596 36168 25648 36174
rect 25596 36110 25648 36116
rect 4620 36032 4672 36038
rect 4620 35974 4672 35980
rect 4632 35894 4660 35974
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 4632 35866 4936 35894
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 940 35080 992 35086
rect 940 35022 992 35028
rect 952 34649 980 35022
rect 3884 34944 3936 34950
rect 3884 34886 3936 34892
rect 938 34640 994 34649
rect 938 34575 994 34584
rect 940 32904 992 32910
rect 940 32846 992 32852
rect 952 32473 980 32846
rect 938 32464 994 32473
rect 938 32399 994 32408
rect 1400 30728 1452 30734
rect 1400 30670 1452 30676
rect 1412 30297 1440 30670
rect 1398 30288 1454 30297
rect 1398 30223 1454 30232
rect 940 28552 992 28558
rect 940 28494 992 28500
rect 952 28121 980 28494
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 938 28112 994 28121
rect 938 28047 994 28056
rect 1596 27674 1624 28358
rect 1584 27668 1636 27674
rect 1584 27610 1636 27616
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 26217 1440 26318
rect 1398 26208 1454 26217
rect 1398 26143 1454 26152
rect 940 24200 992 24206
rect 940 24142 992 24148
rect 3608 24200 3660 24206
rect 3608 24142 3660 24148
rect 952 23769 980 24142
rect 938 23760 994 23769
rect 938 23695 994 23704
rect 3620 23662 3648 24142
rect 3608 23656 3660 23662
rect 3608 23598 3660 23604
rect 3620 22574 3648 23598
rect 3896 22710 3924 34886
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4712 32768 4764 32774
rect 4712 32710 4764 32716
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4724 31754 4752 32710
rect 4632 31726 4752 31754
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 27464 4120 27470
rect 4068 27406 4120 27412
rect 4080 27062 4108 27406
rect 4068 27056 4120 27062
rect 4068 26998 4120 27004
rect 4080 25838 4108 26998
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26568 4660 31726
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4712 27328 4764 27334
rect 4712 27270 4764 27276
rect 4724 27062 4752 27270
rect 4712 27056 4764 27062
rect 4712 26998 4764 27004
rect 4816 26926 4844 30534
rect 4804 26920 4856 26926
rect 4804 26862 4856 26868
rect 4540 26540 4660 26568
rect 4540 25974 4568 26540
rect 4620 26308 4672 26314
rect 4620 26250 4672 26256
rect 4528 25968 4580 25974
rect 4528 25910 4580 25916
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 4080 25294 4108 25774
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4080 24206 4108 25230
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 4632 23662 4660 26250
rect 4908 25362 4936 35866
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 23664 33992 23716 33998
rect 23664 33934 23716 33940
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 23572 28416 23624 28422
rect 23572 28358 23624 28364
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 23584 28218 23612 28358
rect 23676 28218 23704 33934
rect 25608 28218 25636 36110
rect 34336 36100 34388 36106
rect 34336 36042 34388 36048
rect 34348 35737 34376 36042
rect 34334 35728 34390 35737
rect 34334 35663 34390 35672
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34888 33924 34940 33930
rect 34888 33866 34940 33872
rect 34900 33561 34928 33866
rect 34886 33552 34942 33561
rect 34886 33487 34942 33496
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 33140 31816 33192 31822
rect 33140 31758 33192 31764
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 25596 28212 25648 28218
rect 25596 28154 25648 28160
rect 22928 28144 22980 28150
rect 22928 28086 22980 28092
rect 24860 28144 24912 28150
rect 24860 28086 24912 28092
rect 6000 28076 6052 28082
rect 6000 28018 6052 28024
rect 5908 27872 5960 27878
rect 5908 27814 5960 27820
rect 5920 27402 5948 27814
rect 5908 27396 5960 27402
rect 5908 27338 5960 27344
rect 6012 27334 6040 28018
rect 22192 28008 22244 28014
rect 22192 27950 22244 27956
rect 22204 27674 22232 27950
rect 22652 27872 22704 27878
rect 22652 27814 22704 27820
rect 22664 27674 22692 27814
rect 22940 27674 22968 28086
rect 23848 28076 23900 28082
rect 23848 28018 23900 28024
rect 23860 27674 23888 28018
rect 22192 27668 22244 27674
rect 22192 27610 22244 27616
rect 22652 27668 22704 27674
rect 22652 27610 22704 27616
rect 22928 27668 22980 27674
rect 22928 27610 22980 27616
rect 23848 27668 23900 27674
rect 23848 27610 23900 27616
rect 11980 27600 12032 27606
rect 11980 27542 12032 27548
rect 22376 27600 22428 27606
rect 22376 27542 22428 27548
rect 7012 27396 7064 27402
rect 7012 27338 7064 27344
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 6552 27328 6604 27334
rect 6552 27270 6604 27276
rect 5908 26920 5960 26926
rect 5908 26862 5960 26868
rect 5448 26376 5500 26382
rect 5448 26318 5500 26324
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 5460 24818 5488 26318
rect 5540 26308 5592 26314
rect 5540 26250 5592 26256
rect 5552 25974 5580 26250
rect 5632 26240 5684 26246
rect 5632 26182 5684 26188
rect 5540 25968 5592 25974
rect 5540 25910 5592 25916
rect 5644 25498 5672 26182
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 5448 24812 5500 24818
rect 5448 24754 5500 24760
rect 5172 24608 5224 24614
rect 5172 24550 5224 24556
rect 5184 24138 5212 24550
rect 5172 24132 5224 24138
rect 5172 24074 5224 24080
rect 4988 23792 5040 23798
rect 4988 23734 5040 23740
rect 4620 23656 4672 23662
rect 4620 23598 4672 23604
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 5000 23322 5028 23734
rect 5460 23322 5488 24754
rect 4988 23316 5040 23322
rect 4988 23258 5040 23264
rect 5448 23316 5500 23322
rect 5448 23258 5500 23264
rect 5460 22778 5488 23258
rect 5632 22976 5684 22982
rect 5632 22918 5684 22924
rect 5448 22772 5500 22778
rect 5448 22714 5500 22720
rect 3884 22704 3936 22710
rect 3884 22646 3936 22652
rect 3608 22568 3660 22574
rect 3608 22510 3660 22516
rect 940 22024 992 22030
rect 940 21966 992 21972
rect 952 21593 980 21966
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 1596 21690 1624 21830
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 3620 21486 3648 22510
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 4804 21616 4856 21622
rect 4804 21558 4856 21564
rect 3608 21480 3660 21486
rect 3608 21422 3660 21428
rect 940 19848 992 19854
rect 940 19790 992 19796
rect 952 19417 980 19790
rect 938 19408 994 19417
rect 3620 19378 3648 21422
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4816 21146 4844 21558
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 5368 21010 5396 21830
rect 5460 21146 5488 22714
rect 5644 21554 5672 22918
rect 5816 22228 5868 22234
rect 5816 22170 5868 22176
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 5828 21486 5856 22170
rect 5920 22094 5948 26862
rect 6012 26586 6040 27270
rect 6564 26790 6592 27270
rect 6552 26784 6604 26790
rect 6552 26726 6604 26732
rect 6000 26580 6052 26586
rect 6000 26522 6052 26528
rect 6564 25702 6592 26726
rect 6920 25764 6972 25770
rect 6920 25706 6972 25712
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 6552 25696 6604 25702
rect 6552 25638 6604 25644
rect 6644 25696 6696 25702
rect 6644 25638 6696 25644
rect 6104 25158 6132 25638
rect 6656 25514 6684 25638
rect 6564 25486 6684 25514
rect 6184 25220 6236 25226
rect 6184 25162 6236 25168
rect 6092 25152 6144 25158
rect 6092 25094 6144 25100
rect 6104 24614 6132 25094
rect 6092 24608 6144 24614
rect 6092 24550 6144 24556
rect 6000 23656 6052 23662
rect 6000 23598 6052 23604
rect 6012 22234 6040 23598
rect 6104 22982 6132 24550
rect 6196 23730 6224 25162
rect 6184 23724 6236 23730
rect 6184 23666 6236 23672
rect 6092 22976 6144 22982
rect 6092 22918 6144 22924
rect 6276 22568 6328 22574
rect 6276 22510 6328 22516
rect 6000 22228 6052 22234
rect 6000 22170 6052 22176
rect 5920 22066 6224 22094
rect 5920 22030 5948 22066
rect 6196 22030 6224 22066
rect 5908 22024 5960 22030
rect 5908 21966 5960 21972
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6012 21690 6040 21966
rect 6000 21684 6052 21690
rect 6000 21626 6052 21632
rect 5816 21480 5868 21486
rect 5816 21422 5868 21428
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 938 19343 994 19352
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3620 18834 3648 19314
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3620 17746 3648 18770
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 3608 17740 3660 17746
rect 3608 17682 3660 17688
rect 940 17672 992 17678
rect 940 17614 992 17620
rect 952 17241 980 17614
rect 938 17232 994 17241
rect 938 17167 994 17176
rect 3620 16658 3648 17682
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4632 16658 4660 19654
rect 5264 18896 5316 18902
rect 5264 18838 5316 18844
rect 4804 18828 4856 18834
rect 4804 18770 4856 18776
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 3608 16652 3660 16658
rect 3608 16594 3660 16600
rect 4620 16652 4672 16658
rect 4620 16594 4672 16600
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15201 1440 15438
rect 1398 15192 1454 15201
rect 1398 15127 1454 15136
rect 3620 15026 3648 16594
rect 4620 16516 4672 16522
rect 4620 16458 4672 16464
rect 4632 16250 4660 16458
rect 4724 16250 4752 17138
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4356 15094 4384 15302
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4080 13938 4108 14962
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 14618 4752 16186
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 4080 13394 4108 13874
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 952 12889 980 13262
rect 938 12880 994 12889
rect 938 12815 994 12824
rect 4080 12434 4108 13330
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3896 12406 4108 12434
rect 3896 12306 3924 12406
rect 4724 12322 4752 13670
rect 3884 12300 3936 12306
rect 3884 12242 3936 12248
rect 4632 12294 4752 12322
rect 3896 11150 3924 12242
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 3884 11144 3936 11150
rect 3884 11086 3936 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 940 8968 992 8974
rect 940 8910 992 8916
rect 952 8537 980 8910
rect 4528 8900 4580 8906
rect 4528 8842 4580 8848
rect 938 8528 994 8537
rect 938 8463 994 8472
rect 4540 8378 4568 8842
rect 4632 8650 4660 12294
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4724 8786 4752 12106
rect 4816 9178 4844 18770
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4908 18426 4936 18634
rect 4896 18420 4948 18426
rect 4896 18362 4948 18368
rect 4896 17604 4948 17610
rect 4896 17546 4948 17552
rect 4908 17338 4936 17546
rect 4896 17332 4948 17338
rect 4896 17274 4948 17280
rect 5276 16114 5304 18838
rect 5460 18426 5488 21082
rect 6184 21072 6236 21078
rect 6184 21014 6236 21020
rect 6000 20868 6052 20874
rect 6000 20810 6052 20816
rect 5816 19916 5868 19922
rect 5816 19858 5868 19864
rect 5828 19446 5856 19858
rect 6012 19854 6040 20810
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 6092 19848 6144 19854
rect 6092 19790 6144 19796
rect 5816 19440 5868 19446
rect 5816 19382 5868 19388
rect 5828 18766 5856 19382
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5920 18426 5948 19314
rect 6012 19174 6040 19790
rect 6104 19242 6132 19790
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 18902 6040 19110
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5460 17338 5488 18362
rect 5920 17882 5948 18362
rect 5908 17876 5960 17882
rect 5908 17818 5960 17824
rect 5920 17338 5948 17818
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5092 14618 5120 15030
rect 5276 14618 5304 16050
rect 5080 14612 5132 14618
rect 5080 14554 5132 14560
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5920 14550 5948 17274
rect 6196 15706 6224 21014
rect 6288 20942 6316 22510
rect 6564 21078 6592 25486
rect 6932 25294 6960 25706
rect 7024 25294 7052 27338
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11900 26994 11928 27270
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11992 26926 12020 27542
rect 12440 27532 12492 27538
rect 12440 27474 12492 27480
rect 14924 27532 14976 27538
rect 14924 27474 14976 27480
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11716 25974 11744 26318
rect 11796 26240 11848 26246
rect 11796 26182 11848 26188
rect 11704 25968 11756 25974
rect 11704 25910 11756 25916
rect 11808 25906 11836 26182
rect 10692 25900 10744 25906
rect 10692 25842 10744 25848
rect 10784 25900 10836 25906
rect 10784 25842 10836 25848
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10152 25498 10180 25638
rect 10704 25498 10732 25842
rect 10796 25498 10824 25842
rect 11704 25696 11756 25702
rect 11704 25638 11756 25644
rect 8024 25492 8076 25498
rect 8024 25434 8076 25440
rect 10140 25492 10192 25498
rect 10140 25434 10192 25440
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 7012 25288 7064 25294
rect 7012 25230 7064 25236
rect 7288 25288 7340 25294
rect 7288 25230 7340 25236
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7840 25288 7892 25294
rect 7840 25230 7892 25236
rect 6932 24818 6960 25230
rect 7024 24954 7052 25230
rect 7300 24954 7328 25230
rect 7012 24948 7064 24954
rect 7012 24890 7064 24896
rect 7288 24948 7340 24954
rect 7288 24890 7340 24896
rect 6920 24812 6972 24818
rect 6920 24754 6972 24760
rect 7300 24138 7328 24890
rect 7288 24132 7340 24138
rect 7288 24074 7340 24080
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6920 23792 6972 23798
rect 6920 23734 6972 23740
rect 6828 23724 6880 23730
rect 6828 23666 6880 23672
rect 6840 23186 6868 23666
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6840 22642 6868 23122
rect 6932 23118 6960 23734
rect 7116 23322 7144 24006
rect 7300 23798 7328 24074
rect 7392 24070 7420 25230
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7656 25152 7708 25158
rect 7656 25094 7708 25100
rect 7484 24818 7512 25094
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7288 23792 7340 23798
rect 7288 23734 7340 23740
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 6920 23112 6972 23118
rect 6972 23060 7144 23066
rect 6920 23054 7144 23060
rect 6932 23038 7144 23054
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6920 22636 6972 22642
rect 6920 22578 6972 22584
rect 6644 22160 6696 22166
rect 6644 22102 6696 22108
rect 6656 21554 6684 22102
rect 6840 22094 6868 22578
rect 6932 22234 6960 22578
rect 6920 22228 6972 22234
rect 6920 22170 6972 22176
rect 6748 22066 6868 22094
rect 6644 21548 6696 21554
rect 6644 21490 6696 21496
rect 6552 21072 6604 21078
rect 6552 21014 6604 21020
rect 6748 20942 6776 22066
rect 6932 21554 6960 22170
rect 6920 21548 6972 21554
rect 6920 21490 6972 21496
rect 6276 20936 6328 20942
rect 6276 20878 6328 20884
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6288 20058 6316 20878
rect 7116 20618 7144 23038
rect 7300 20618 7328 23734
rect 7668 23730 7696 25094
rect 7852 24886 7880 25230
rect 7932 25220 7984 25226
rect 7932 25162 7984 25168
rect 7944 24954 7972 25162
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 7840 24880 7892 24886
rect 7840 24822 7892 24828
rect 8036 24342 8064 25434
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 8208 25152 8260 25158
rect 8128 25100 8208 25106
rect 8128 25094 8260 25100
rect 8128 25078 8248 25094
rect 8024 24336 8076 24342
rect 8024 24278 8076 24284
rect 8036 24206 8064 24278
rect 8024 24200 8076 24206
rect 8024 24142 8076 24148
rect 8036 23730 8064 24142
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 8024 23724 8076 23730
rect 8024 23666 8076 23672
rect 8128 23202 8156 25078
rect 9968 24886 9996 25298
rect 10152 25226 10180 25434
rect 11716 25362 11744 25638
rect 11808 25498 11836 25842
rect 11796 25492 11848 25498
rect 11796 25434 11848 25440
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10140 25220 10192 25226
rect 10140 25162 10192 25168
rect 9956 24880 10008 24886
rect 9956 24822 10008 24828
rect 10796 24818 10824 25230
rect 11152 25220 11204 25226
rect 11152 25162 11204 25168
rect 11612 25220 11664 25226
rect 11612 25162 11664 25168
rect 11164 24954 11192 25162
rect 11152 24948 11204 24954
rect 11152 24890 11204 24896
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 10784 24812 10836 24818
rect 10784 24754 10836 24760
rect 8496 24206 8524 24754
rect 8852 24404 8904 24410
rect 8852 24346 8904 24352
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 8220 23322 8248 23598
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8128 23174 8248 23202
rect 7932 23112 7984 23118
rect 7932 23054 7984 23060
rect 7944 22642 7972 23054
rect 7932 22636 7984 22642
rect 7760 22596 7932 22624
rect 7760 22166 7788 22596
rect 7932 22578 7984 22584
rect 8116 22228 8168 22234
rect 8116 22170 8168 22176
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 8128 22030 8156 22170
rect 8220 22166 8248 23174
rect 8300 22976 8352 22982
rect 8300 22918 8352 22924
rect 8576 22976 8628 22982
rect 8576 22918 8628 22924
rect 8312 22506 8340 22918
rect 8588 22642 8616 22918
rect 8864 22710 8892 24346
rect 9232 24274 9260 24754
rect 11624 24750 11652 25162
rect 11716 24954 11744 25298
rect 11796 25288 11848 25294
rect 11796 25230 11848 25236
rect 11704 24948 11756 24954
rect 11704 24890 11756 24896
rect 10508 24744 10560 24750
rect 10508 24686 10560 24692
rect 11612 24744 11664 24750
rect 11612 24686 11664 24692
rect 9220 24268 9272 24274
rect 9220 24210 9272 24216
rect 9232 23866 9260 24210
rect 10520 24138 10548 24686
rect 11336 24676 11388 24682
rect 11336 24618 11388 24624
rect 11348 24206 11376 24618
rect 11808 24410 11836 25230
rect 11888 25152 11940 25158
rect 11888 25094 11940 25100
rect 11900 24410 11928 25094
rect 11992 24410 12020 26862
rect 12452 26586 12480 27474
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 12544 27130 12572 27406
rect 13004 27130 13032 27406
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 12532 27124 12584 27130
rect 12532 27066 12584 27072
rect 12992 27124 13044 27130
rect 12992 27066 13044 27072
rect 12992 26988 13044 26994
rect 13096 26976 13124 27270
rect 14476 27130 14504 27338
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14464 27124 14516 27130
rect 14464 27066 14516 27072
rect 13044 26948 13124 26976
rect 13176 26988 13228 26994
rect 12992 26930 13044 26936
rect 13176 26930 13228 26936
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 13004 26790 13032 26930
rect 12992 26784 13044 26790
rect 12992 26726 13044 26732
rect 12440 26580 12492 26586
rect 12440 26522 12492 26528
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12268 25838 12296 26318
rect 12808 26308 12860 26314
rect 12808 26250 12860 26256
rect 12820 25906 12848 26250
rect 12808 25900 12860 25906
rect 12808 25842 12860 25848
rect 12256 25832 12308 25838
rect 12256 25774 12308 25780
rect 12164 25696 12216 25702
rect 12164 25638 12216 25644
rect 12176 25362 12204 25638
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 12532 25424 12584 25430
rect 12532 25366 12584 25372
rect 12164 25356 12216 25362
rect 12164 25298 12216 25304
rect 12544 25294 12572 25366
rect 12532 25288 12584 25294
rect 12532 25230 12584 25236
rect 12072 25152 12124 25158
rect 12072 25094 12124 25100
rect 12084 24954 12112 25094
rect 12072 24948 12124 24954
rect 12072 24890 12124 24896
rect 11796 24404 11848 24410
rect 11796 24346 11848 24352
rect 11888 24404 11940 24410
rect 11888 24346 11940 24352
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12256 24336 12308 24342
rect 12256 24278 12308 24284
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 11428 24200 11480 24206
rect 11428 24142 11480 24148
rect 11980 24200 12032 24206
rect 12032 24160 12112 24188
rect 11980 24142 12032 24148
rect 9680 24132 9732 24138
rect 9680 24074 9732 24080
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9508 22778 9536 24006
rect 9496 22772 9548 22778
rect 9496 22714 9548 22720
rect 8852 22704 8904 22710
rect 8852 22646 8904 22652
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8760 22636 8812 22642
rect 8760 22578 8812 22584
rect 8300 22500 8352 22506
rect 8300 22442 8352 22448
rect 8588 22166 8616 22578
rect 8772 22522 8800 22578
rect 8680 22494 8800 22522
rect 8208 22160 8260 22166
rect 8208 22102 8260 22108
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 8116 22024 8168 22030
rect 8116 21966 8168 21972
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21554 7972 21830
rect 7932 21548 7984 21554
rect 7932 21490 7984 21496
rect 6932 20590 7144 20618
rect 7208 20590 7328 20618
rect 6276 20052 6328 20058
rect 6276 19994 6328 20000
rect 6276 19848 6328 19854
rect 6276 19790 6328 19796
rect 6288 19514 6316 19790
rect 6276 19508 6328 19514
rect 6276 19450 6328 19456
rect 6460 19236 6512 19242
rect 6460 19178 6512 19184
rect 6472 18834 6500 19178
rect 6460 18828 6512 18834
rect 6460 18770 6512 18776
rect 6932 16674 6960 20590
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 19854 7144 20402
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7116 18766 7144 19790
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 7024 18290 7052 18634
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 7024 17678 7052 18226
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 6748 16646 6960 16674
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6380 16250 6408 16526
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6472 15638 6500 16050
rect 6552 15972 6604 15978
rect 6552 15914 6604 15920
rect 6644 15972 6696 15978
rect 6644 15914 6696 15920
rect 6460 15632 6512 15638
rect 6460 15574 6512 15580
rect 6564 15502 6592 15914
rect 6656 15638 6684 15914
rect 6748 15910 6776 16646
rect 6828 16584 6880 16590
rect 6828 16526 6880 16532
rect 6840 16114 6868 16526
rect 6828 16108 6880 16114
rect 6828 16050 6880 16056
rect 6736 15904 6788 15910
rect 6736 15846 6788 15852
rect 6644 15632 6696 15638
rect 6644 15574 6696 15580
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6564 14822 6592 15438
rect 6748 15162 6776 15846
rect 6840 15706 6868 16050
rect 6828 15700 6880 15706
rect 6828 15642 6880 15648
rect 6920 15632 6972 15638
rect 6920 15574 6972 15580
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 5908 14544 5960 14550
rect 5908 14486 5960 14492
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5460 13938 5488 14214
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 5092 12986 5120 13194
rect 5552 12986 5580 14350
rect 5920 14074 5948 14486
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6104 14006 6132 14554
rect 6748 14414 6776 15098
rect 6932 15094 6960 15574
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 6840 14618 6868 14826
rect 6828 14612 6880 14618
rect 6828 14554 6880 14560
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6380 13530 6408 14010
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5184 11898 5212 12106
rect 5552 11898 5580 12922
rect 6184 12436 6236 12442
rect 6380 12434 6408 13466
rect 7116 13326 7144 18702
rect 7208 15706 7236 20590
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19854 7328 20402
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8128 19514 8156 19654
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8036 19242 8064 19314
rect 8024 19236 8076 19242
rect 8024 19178 8076 19184
rect 8036 18970 8064 19178
rect 8024 18964 8076 18970
rect 8024 18906 8076 18912
rect 8128 18834 8156 19450
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7576 18630 7604 18702
rect 7748 18692 7800 18698
rect 7748 18634 7800 18640
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7760 18426 7788 18634
rect 7748 18420 7800 18426
rect 7748 18362 7800 18368
rect 7760 17678 7788 18362
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7944 15502 7972 15982
rect 8220 15502 8248 22102
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8404 21350 8432 21966
rect 8680 21690 8708 22494
rect 8864 22094 8892 22646
rect 9404 22228 9456 22234
rect 9404 22170 9456 22176
rect 8772 22066 8892 22094
rect 8668 21684 8720 21690
rect 8588 21644 8668 21672
rect 8392 21344 8444 21350
rect 8392 21286 8444 21292
rect 8404 18970 8432 21286
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8588 17105 8616 21644
rect 8668 21626 8720 21632
rect 8668 20868 8720 20874
rect 8668 20810 8720 20816
rect 8680 20534 8708 20810
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8772 17202 8800 22066
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 8944 21004 8996 21010
rect 8944 20946 8996 20952
rect 8956 20534 8984 20946
rect 9324 20942 9352 21014
rect 9416 20942 9444 22170
rect 9508 21010 9536 22714
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9496 21004 9548 21010
rect 9496 20946 9548 20952
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9324 20602 9352 20878
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8956 19854 8984 20470
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8944 19848 8996 19854
rect 8944 19790 8996 19796
rect 9140 19718 9168 20198
rect 9324 20058 9352 20538
rect 9312 20052 9364 20058
rect 9312 19994 9364 20000
rect 9310 19952 9366 19961
rect 9310 19887 9366 19896
rect 9220 19848 9272 19854
rect 9324 19836 9352 19887
rect 9272 19808 9352 19836
rect 9220 19790 9272 19796
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17610 8984 18226
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8956 17270 8984 17546
rect 9048 17542 9076 18158
rect 9232 17678 9260 19790
rect 9416 18426 9444 20878
rect 9496 20800 9548 20806
rect 9494 20768 9496 20777
rect 9548 20768 9550 20777
rect 9494 20703 9550 20712
rect 9496 20392 9548 20398
rect 9496 20334 9548 20340
rect 9508 19352 9536 20334
rect 9496 19346 9548 19352
rect 9496 19288 9548 19294
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9220 17672 9272 17678
rect 9600 17626 9628 22510
rect 9692 22506 9720 24074
rect 11440 23730 11468 24142
rect 11888 24132 11940 24138
rect 11888 24074 11940 24080
rect 11900 24018 11928 24074
rect 11900 23990 12020 24018
rect 9772 23724 9824 23730
rect 9772 23666 9824 23672
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 11428 23724 11480 23730
rect 11428 23666 11480 23672
rect 9784 23118 9812 23666
rect 10428 23118 10456 23666
rect 11992 23594 12020 23990
rect 12084 23730 12112 24160
rect 12072 23724 12124 23730
rect 12072 23666 12124 23672
rect 10508 23588 10560 23594
rect 10508 23530 10560 23536
rect 11980 23588 12032 23594
rect 11980 23530 12032 23536
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 10416 23112 10468 23118
rect 10416 23054 10468 23060
rect 9680 22500 9732 22506
rect 9680 22442 9732 22448
rect 10232 22500 10284 22506
rect 10232 22442 10284 22448
rect 10244 22098 10272 22442
rect 10324 22432 10376 22438
rect 10324 22374 10376 22380
rect 10336 22234 10364 22374
rect 10428 22234 10456 23054
rect 10324 22228 10376 22234
rect 10324 22170 10376 22176
rect 10416 22228 10468 22234
rect 10416 22170 10468 22176
rect 10232 22092 10284 22098
rect 10232 22034 10284 22040
rect 9864 22024 9916 22030
rect 9864 21966 9916 21972
rect 9876 21690 9904 21966
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9680 21616 9732 21622
rect 9680 21558 9732 21564
rect 9692 20602 9720 21558
rect 9956 21548 10008 21554
rect 9956 21490 10008 21496
rect 9862 21448 9918 21457
rect 9772 21412 9824 21418
rect 9862 21383 9864 21392
rect 9772 21354 9824 21360
rect 9916 21383 9918 21392
rect 9864 21354 9916 21360
rect 9784 20942 9812 21354
rect 9968 20942 9996 21490
rect 10060 21486 10088 21830
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9772 20936 9824 20942
rect 9772 20878 9824 20884
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 9784 20602 9812 20878
rect 9956 20800 10008 20806
rect 10060 20788 10088 21422
rect 10140 21344 10192 21350
rect 10140 21286 10192 21292
rect 10152 20942 10180 21286
rect 10244 21078 10272 22034
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10232 21072 10284 21078
rect 10232 21014 10284 21020
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 10336 20806 10364 21626
rect 10416 21480 10468 21486
rect 10416 21422 10468 21428
rect 10008 20760 10088 20788
rect 10324 20800 10376 20806
rect 9956 20742 10008 20748
rect 10324 20742 10376 20748
rect 10230 20632 10286 20641
rect 9680 20596 9732 20602
rect 9680 20538 9732 20544
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 10152 20590 10230 20618
rect 9772 20460 9824 20466
rect 9772 20402 9824 20408
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9692 19446 9720 20334
rect 9784 20058 9812 20402
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9864 18216 9916 18222
rect 9864 18158 9916 18164
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17678 9812 18090
rect 9220 17614 9272 17620
rect 9036 17536 9088 17542
rect 9036 17478 9088 17484
rect 9048 17338 9076 17478
rect 9036 17332 9088 17338
rect 9036 17274 9088 17280
rect 8944 17264 8996 17270
rect 8944 17206 8996 17212
rect 9048 17202 9076 17274
rect 8760 17196 8812 17202
rect 8760 17138 8812 17144
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8668 17128 8720 17134
rect 8574 17096 8630 17105
rect 8668 17070 8720 17076
rect 8574 17031 8630 17040
rect 8588 16998 8616 17031
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8496 16726 8524 16934
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8588 16182 8616 16594
rect 8484 16176 8536 16182
rect 8484 16118 8536 16124
rect 8576 16176 8628 16182
rect 8576 16118 8628 16124
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8404 15502 8432 15982
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 7196 15428 7248 15434
rect 7196 15370 7248 15376
rect 7208 15026 7236 15370
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 7208 14414 7236 14962
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 6236 12406 6408 12434
rect 6184 12378 6236 12384
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5540 11892 5592 11898
rect 5540 11834 5592 11840
rect 5552 11778 5580 11834
rect 5552 11750 5672 11778
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5552 10810 5580 11018
rect 5644 10810 5672 11750
rect 6196 11354 6224 12378
rect 7208 12170 7236 14350
rect 7300 13326 7328 15438
rect 8220 14958 8248 15438
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7472 14884 7524 14890
rect 7472 14826 7524 14832
rect 7484 13938 7512 14826
rect 7668 13938 7696 14894
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 7852 13326 7880 14282
rect 8404 13530 8432 15438
rect 8496 14414 8524 16118
rect 8680 15026 8708 17070
rect 8772 16794 8800 17138
rect 8760 16788 8812 16794
rect 8760 16730 8812 16736
rect 8864 15706 8892 17138
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8852 15700 8904 15706
rect 8852 15642 8904 15648
rect 8956 15094 8984 16458
rect 9048 16182 9076 17138
rect 9232 17066 9260 17614
rect 9508 17598 9628 17626
rect 9772 17672 9824 17678
rect 9772 17614 9824 17620
rect 9312 17536 9364 17542
rect 9312 17478 9364 17484
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9324 17134 9352 17478
rect 9416 17202 9444 17478
rect 9404 17196 9456 17202
rect 9404 17138 9456 17144
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9416 16454 9444 17138
rect 9508 16658 9536 17598
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9600 17338 9628 17478
rect 9588 17332 9640 17338
rect 9588 17274 9640 17280
rect 9876 17202 9904 18158
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 9680 17128 9732 17134
rect 9600 17105 9680 17116
rect 9586 17096 9680 17105
rect 9642 17088 9680 17096
rect 9680 17070 9732 17076
rect 9586 17031 9642 17040
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9496 16516 9548 16522
rect 9600 16504 9628 17031
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9548 16476 9628 16504
rect 9496 16458 9548 16464
rect 9404 16448 9456 16454
rect 9404 16390 9456 16396
rect 9508 16182 9536 16458
rect 9036 16176 9088 16182
rect 9036 16118 9088 16124
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9508 15162 9536 16118
rect 9968 15910 9996 16594
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9956 15904 10008 15910
rect 9784 15864 9956 15892
rect 9784 15502 9812 15864
rect 9956 15846 10008 15852
rect 10060 15502 10088 15982
rect 9680 15496 9732 15502
rect 9680 15438 9732 15444
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9692 15094 9720 15438
rect 9784 15094 9812 15438
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8680 13802 8708 14962
rect 8956 14074 8984 15030
rect 9784 14958 9812 15030
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 10060 14618 10088 15438
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10152 14346 10180 20590
rect 10230 20567 10286 20576
rect 10232 20392 10284 20398
rect 10232 20334 10284 20340
rect 10244 19922 10272 20334
rect 10336 20058 10364 20742
rect 10428 20602 10456 21422
rect 10520 20602 10548 23530
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 10876 22160 10928 22166
rect 10928 22108 11008 22114
rect 10876 22102 11008 22108
rect 10888 22086 11008 22102
rect 10600 22024 10652 22030
rect 10600 21966 10652 21972
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10508 20596 10560 20602
rect 10508 20538 10560 20544
rect 10612 20516 10640 21966
rect 10784 21888 10836 21894
rect 10784 21830 10836 21836
rect 10796 21622 10824 21830
rect 10784 21616 10836 21622
rect 10784 21558 10836 21564
rect 10876 21480 10928 21486
rect 10876 21422 10928 21428
rect 10888 21010 10916 21422
rect 10980 21010 11008 22086
rect 11244 22024 11296 22030
rect 11244 21966 11296 21972
rect 11256 21554 11284 21966
rect 11336 21888 11388 21894
rect 11336 21830 11388 21836
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 10876 21004 10928 21010
rect 10876 20946 10928 20952
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 11256 20874 11284 21490
rect 11348 21078 11376 21830
rect 11612 21480 11664 21486
rect 11610 21448 11612 21457
rect 11664 21448 11666 21457
rect 11610 21383 11666 21392
rect 11336 21072 11388 21078
rect 11336 21014 11388 21020
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 10784 20528 10836 20534
rect 10612 20488 10784 20516
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 10612 19990 10640 20488
rect 10784 20470 10836 20476
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 10600 19984 10652 19990
rect 10600 19926 10652 19932
rect 10232 19916 10284 19922
rect 10232 19858 10284 19864
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 19378 10640 19790
rect 10888 19446 10916 20266
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 10876 19440 10928 19446
rect 10876 19382 10928 19388
rect 10600 19372 10652 19378
rect 10600 19314 10652 19320
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 17814 10364 18566
rect 10692 18216 10744 18222
rect 10692 18158 10744 18164
rect 10704 17882 10732 18158
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10324 17808 10376 17814
rect 10324 17750 10376 17756
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 16794 10272 17546
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17066 10732 17478
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10600 16992 10652 16998
rect 10796 16946 10824 17682
rect 10600 16934 10652 16940
rect 10232 16788 10284 16794
rect 10232 16730 10284 16736
rect 10230 16688 10286 16697
rect 10230 16623 10232 16632
rect 10284 16623 10286 16632
rect 10232 16594 10284 16600
rect 10324 16516 10376 16522
rect 10508 16516 10560 16522
rect 10324 16458 10376 16464
rect 10428 16476 10508 16504
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10244 15570 10272 15914
rect 10336 15706 10364 16458
rect 10428 16046 10456 16476
rect 10508 16458 10560 16464
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10428 15502 10456 15982
rect 10416 15496 10468 15502
rect 10416 15438 10468 15444
rect 10428 15094 10456 15438
rect 10416 15088 10468 15094
rect 10416 15030 10468 15036
rect 10612 14822 10640 16934
rect 10704 16918 10824 16946
rect 10704 15638 10732 16918
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10796 16454 10824 16730
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10796 15502 10824 16390
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 14929 10732 14962
rect 10690 14920 10746 14929
rect 10690 14855 10746 14864
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 10140 14340 10192 14346
rect 10140 14282 10192 14288
rect 10152 14074 10180 14282
rect 8944 14068 8996 14074
rect 8944 14010 8996 14016
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10244 13938 10272 14350
rect 10612 14328 10640 14758
rect 10796 14346 10824 15302
rect 10888 14890 10916 19382
rect 11072 19378 11100 19654
rect 11164 19378 11192 19790
rect 11256 19718 11284 20810
rect 11704 20460 11756 20466
rect 11704 20402 11756 20408
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11624 20058 11652 20334
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11624 19718 11652 19994
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11612 19712 11664 19718
rect 11612 19654 11664 19660
rect 11716 19514 11744 20402
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11702 19408 11758 19417
rect 11060 19372 11112 19378
rect 11060 19314 11112 19320
rect 11152 19372 11204 19378
rect 11702 19343 11704 19352
rect 11152 19314 11204 19320
rect 11756 19343 11758 19352
rect 11704 19314 11756 19320
rect 11072 18306 11100 19314
rect 10968 18284 11020 18290
rect 11072 18278 11192 18306
rect 10968 18226 11020 18232
rect 10980 17882 11008 18226
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 11164 17626 11192 18278
rect 11612 17672 11664 17678
rect 11072 17598 11192 17626
rect 11348 17620 11612 17626
rect 11348 17614 11664 17620
rect 11348 17598 11652 17614
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10876 14884 10928 14890
rect 10876 14826 10928 14832
rect 10980 14618 11008 14962
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11072 14414 11100 17598
rect 11348 17542 11376 17598
rect 11336 17536 11388 17542
rect 11336 17478 11388 17484
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 17338 11468 17478
rect 11428 17332 11480 17338
rect 11428 17274 11480 17280
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 15502 11284 16050
rect 11624 15910 11652 17598
rect 11612 15904 11664 15910
rect 11612 15846 11664 15852
rect 11624 15706 11652 15846
rect 11612 15700 11664 15706
rect 11612 15642 11664 15648
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 11256 15094 11284 15438
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11440 14414 11468 14826
rect 11808 14618 11836 19926
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11702 14512 11758 14521
rect 11702 14447 11758 14456
rect 11716 14414 11744 14447
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 10692 14340 10744 14346
rect 10612 14300 10692 14328
rect 10692 14282 10744 14288
rect 10784 14340 10836 14346
rect 10784 14282 10836 14288
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8392 13524 8444 13530
rect 8392 13466 8444 13472
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7300 12850 7328 13262
rect 7852 12850 7880 13262
rect 10244 12850 10272 13874
rect 10692 13728 10744 13734
rect 10692 13670 10744 13676
rect 10704 13326 10732 13670
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10796 12918 10824 14282
rect 10980 14249 11008 14350
rect 10966 14240 11022 14249
rect 10966 14175 11022 14184
rect 11256 13954 11284 14350
rect 11072 13938 11284 13954
rect 11060 13932 11284 13938
rect 11112 13926 11284 13932
rect 11060 13874 11112 13880
rect 11072 13410 11100 13874
rect 10980 13382 11100 13410
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 6184 11348 6236 11354
rect 6184 11290 6236 11296
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5644 10266 5672 10746
rect 5632 10260 5684 10266
rect 5632 10202 5684 10208
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4724 8758 4936 8786
rect 4632 8622 4752 8650
rect 4540 8350 4660 8378
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 940 6792 992 6798
rect 940 6734 992 6740
rect 952 6361 980 6734
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4632 4826 4660 8350
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 940 4616 992 4622
rect 940 4558 992 4564
rect 952 4185 980 4558
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4724 2650 4752 8622
rect 4908 6662 4936 8758
rect 5000 8634 5028 8842
rect 5644 8634 5672 10202
rect 6196 9178 6224 11290
rect 7300 11218 7328 12786
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10060 12238 10088 12650
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 6184 9172 6236 9178
rect 6184 9114 6236 9120
rect 9968 8838 9996 10406
rect 10060 8906 10088 12174
rect 10244 12170 10272 12786
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 10888 12442 10916 12718
rect 10876 12436 10928 12442
rect 10876 12378 10928 12384
rect 10980 12238 11008 13382
rect 11440 13274 11468 14350
rect 11520 14272 11572 14278
rect 11520 14214 11572 14220
rect 11532 13977 11560 14214
rect 11518 13968 11574 13977
rect 11518 13903 11574 13912
rect 11716 13802 11744 14350
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11808 13394 11836 14554
rect 11796 13388 11848 13394
rect 11796 13330 11848 13336
rect 11348 13246 11468 13274
rect 11704 13252 11756 13258
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11256 12434 11284 12786
rect 11348 12782 11376 13246
rect 11704 13194 11756 13200
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11256 12406 11376 12434
rect 11348 12238 11376 12406
rect 11532 12238 11560 13126
rect 11716 12850 11744 13194
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11900 12442 11928 23462
rect 11992 22574 12020 23530
rect 12084 23118 12112 23666
rect 12268 23118 12296 24278
rect 12348 24268 12400 24274
rect 12452 24256 12480 24346
rect 12400 24228 12480 24256
rect 12348 24210 12400 24216
rect 12544 24188 12572 25230
rect 12636 24954 12664 25434
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12714 24440 12770 24449
rect 12820 24410 12848 25842
rect 13004 25498 13032 26726
rect 13188 26586 13216 26930
rect 14200 26586 14228 26930
rect 14568 26926 14596 27270
rect 14844 27130 14872 27406
rect 14832 27124 14884 27130
rect 14832 27066 14884 27072
rect 14936 26994 14964 27474
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 17132 27328 17184 27334
rect 17132 27270 17184 27276
rect 17684 27328 17736 27334
rect 17684 27270 17736 27276
rect 16028 27056 16080 27062
rect 16028 26998 16080 27004
rect 16764 27056 16816 27062
rect 16764 26998 16816 27004
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15568 26988 15620 26994
rect 15568 26930 15620 26936
rect 15936 26988 15988 26994
rect 15936 26930 15988 26936
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 14188 26580 14240 26586
rect 14188 26522 14240 26528
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14200 26042 14228 26318
rect 14188 26036 14240 26042
rect 14188 25978 14240 25984
rect 13820 25764 13872 25770
rect 13820 25706 13872 25712
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 13176 25152 13228 25158
rect 13176 25094 13228 25100
rect 13188 24886 13216 25094
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13176 24880 13228 24886
rect 13176 24822 13228 24828
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13372 24682 13400 24754
rect 13360 24676 13412 24682
rect 13360 24618 13412 24624
rect 12714 24375 12716 24384
rect 12768 24375 12770 24384
rect 12808 24404 12860 24410
rect 12716 24346 12768 24352
rect 12808 24346 12860 24352
rect 12624 24200 12676 24206
rect 12544 24160 12624 24188
rect 12624 24142 12676 24148
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 13268 24200 13320 24206
rect 13268 24142 13320 24148
rect 12636 23254 12664 24142
rect 12716 24132 12768 24138
rect 12716 24074 12768 24080
rect 12728 23866 12756 24074
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12820 23730 12848 24006
rect 13096 23730 13124 24142
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 13096 23322 13124 23666
rect 13280 23594 13308 24142
rect 13268 23588 13320 23594
rect 13268 23530 13320 23536
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12072 23112 12124 23118
rect 12072 23054 12124 23060
rect 12256 23112 12308 23118
rect 12256 23054 12308 23060
rect 12084 22710 12112 23054
rect 12072 22704 12124 22710
rect 12072 22646 12124 22652
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 11992 19854 12020 22510
rect 12636 22166 12664 23190
rect 12808 23180 12860 23186
rect 12808 23122 12860 23128
rect 12820 23050 12848 23122
rect 13372 23118 13400 24618
rect 13556 24206 13584 24890
rect 13832 24750 13860 25706
rect 14568 24818 14596 26862
rect 15580 26518 15608 26930
rect 15844 26920 15896 26926
rect 15844 26862 15896 26868
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 15568 26512 15620 26518
rect 15568 26454 15620 26460
rect 15120 25906 15148 26454
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15212 25974 15240 26250
rect 15384 26240 15436 26246
rect 15384 26182 15436 26188
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15120 24954 15148 25094
rect 15108 24948 15160 24954
rect 15108 24890 15160 24896
rect 14556 24812 14608 24818
rect 14556 24754 14608 24760
rect 15016 24812 15068 24818
rect 15016 24754 15068 24760
rect 13820 24744 13872 24750
rect 13820 24686 13872 24692
rect 14096 24744 14148 24750
rect 14096 24686 14148 24692
rect 13728 24676 13780 24682
rect 13728 24618 13780 24624
rect 13740 24410 13768 24618
rect 14108 24614 14136 24686
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 13728 24404 13780 24410
rect 13728 24346 13780 24352
rect 13544 24200 13596 24206
rect 13544 24142 13596 24148
rect 13556 23594 13584 24142
rect 13740 23866 13768 24346
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14096 24132 14148 24138
rect 14096 24074 14148 24080
rect 14004 24064 14056 24070
rect 14004 24006 14056 24012
rect 14016 23866 14044 24006
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14108 23662 14136 24074
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14476 23866 14504 24006
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14096 23656 14148 23662
rect 14096 23598 14148 23604
rect 13544 23588 13596 23594
rect 13544 23530 13596 23536
rect 13360 23112 13412 23118
rect 13360 23054 13412 23060
rect 12716 23044 12768 23050
rect 12716 22986 12768 22992
rect 12808 23044 12860 23050
rect 12808 22986 12860 22992
rect 12728 22778 12756 22986
rect 12716 22772 12768 22778
rect 12716 22714 12768 22720
rect 12820 22658 12848 22986
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 12728 22630 12848 22658
rect 12728 22506 12756 22630
rect 12716 22500 12768 22506
rect 12716 22442 12768 22448
rect 12624 22160 12676 22166
rect 12624 22102 12676 22108
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12544 21690 12572 21966
rect 12532 21684 12584 21690
rect 12532 21626 12584 21632
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12176 19854 12204 20198
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 12164 19848 12216 19854
rect 12164 19790 12216 19796
rect 12072 19780 12124 19786
rect 12072 19722 12124 19728
rect 12084 19417 12112 19722
rect 12070 19408 12126 19417
rect 11992 19352 12070 19360
rect 11992 19343 12126 19352
rect 12176 19360 12204 19790
rect 12268 19514 12296 20266
rect 12360 19922 12388 20538
rect 12532 19984 12584 19990
rect 12532 19926 12584 19932
rect 12348 19916 12400 19922
rect 12348 19858 12400 19864
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12360 19378 12388 19654
rect 12256 19372 12308 19378
rect 11992 19332 12112 19343
rect 12176 19332 12256 19360
rect 11992 14890 12020 19332
rect 12256 19314 12308 19320
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12544 19242 12572 19926
rect 12636 19854 12664 22102
rect 12728 20448 12756 22442
rect 13280 22166 13308 22918
rect 13372 22642 13400 23054
rect 14832 22976 14884 22982
rect 14832 22918 14884 22924
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 14464 22568 14516 22574
rect 14464 22510 14516 22516
rect 13268 22160 13320 22166
rect 13268 22102 13320 22108
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 12808 21888 12860 21894
rect 12808 21830 12860 21836
rect 12900 21888 12952 21894
rect 12900 21830 12952 21836
rect 12820 21554 12848 21830
rect 12808 21548 12860 21554
rect 12808 21490 12860 21496
rect 12912 21486 12940 21830
rect 12992 21616 13044 21622
rect 12992 21558 13044 21564
rect 12900 21480 12952 21486
rect 12900 21422 12952 21428
rect 13004 21146 13032 21558
rect 13096 21146 13124 22034
rect 14476 22030 14504 22510
rect 14568 22438 14596 22578
rect 14556 22432 14608 22438
rect 14556 22374 14608 22380
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 14464 22024 14516 22030
rect 14464 21966 14516 21972
rect 13268 21888 13320 21894
rect 13268 21830 13320 21836
rect 13280 21418 13308 21830
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13280 21298 13308 21354
rect 13280 21270 13400 21298
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 13268 21140 13320 21146
rect 13268 21082 13320 21088
rect 13280 20942 13308 21082
rect 13268 20936 13320 20942
rect 13268 20878 13320 20884
rect 13372 20806 13400 21270
rect 13556 21146 13584 21966
rect 14660 21962 14688 22578
rect 14844 22574 14872 22918
rect 14832 22568 14884 22574
rect 14832 22510 14884 22516
rect 14844 22234 14872 22510
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14936 22030 14964 24142
rect 15028 22778 15056 24754
rect 15106 24440 15162 24449
rect 15106 24375 15108 24384
rect 15160 24375 15162 24384
rect 15108 24346 15160 24352
rect 15016 22772 15068 22778
rect 15016 22714 15068 22720
rect 15028 22030 15056 22714
rect 15120 22574 15148 24346
rect 15212 24206 15240 25910
rect 15396 25702 15424 26182
rect 15580 25906 15608 26454
rect 15568 25900 15620 25906
rect 15568 25842 15620 25848
rect 15660 25900 15712 25906
rect 15660 25842 15712 25848
rect 15384 25696 15436 25702
rect 15384 25638 15436 25644
rect 15396 25294 15424 25638
rect 15672 25430 15700 25842
rect 15856 25498 15884 26862
rect 15948 26042 15976 26930
rect 16040 26382 16068 26998
rect 16120 26852 16172 26858
rect 16120 26794 16172 26800
rect 16028 26376 16080 26382
rect 16028 26318 16080 26324
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16040 25838 16068 26318
rect 16132 26314 16160 26794
rect 16776 26790 16804 26998
rect 17040 26852 17092 26858
rect 17040 26794 17092 26800
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16776 26314 16804 26726
rect 17052 26518 17080 26794
rect 17144 26518 17172 27270
rect 17592 27056 17644 27062
rect 17592 26998 17644 27004
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 17132 26512 17184 26518
rect 17132 26454 17184 26460
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16764 26308 16816 26314
rect 16764 26250 16816 26256
rect 16028 25832 16080 25838
rect 16028 25774 16080 25780
rect 15844 25492 15896 25498
rect 15844 25434 15896 25440
rect 15660 25424 15712 25430
rect 15660 25366 15712 25372
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15396 24954 15424 25230
rect 15476 25152 15528 25158
rect 15476 25094 15528 25100
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15488 24818 15516 25094
rect 15476 24812 15528 24818
rect 15476 24754 15528 24760
rect 15660 24812 15712 24818
rect 15660 24754 15712 24760
rect 15672 24342 15700 24754
rect 16132 24750 16160 26250
rect 16396 25900 16448 25906
rect 16396 25842 16448 25848
rect 16408 25430 16436 25842
rect 17144 25838 17172 26454
rect 17604 26314 17632 26998
rect 17696 26926 17724 27270
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17684 26920 17736 26926
rect 17684 26862 17736 26868
rect 17788 26314 17816 27066
rect 18156 26858 18184 27406
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18524 26994 18552 27270
rect 18984 26994 19012 27474
rect 22388 27470 22416 27542
rect 24124 27532 24176 27538
rect 24124 27474 24176 27480
rect 19248 27464 19300 27470
rect 19248 27406 19300 27412
rect 21824 27464 21876 27470
rect 21824 27406 21876 27412
rect 22192 27464 22244 27470
rect 22192 27406 22244 27412
rect 22376 27464 22428 27470
rect 22376 27406 22428 27412
rect 19156 27328 19208 27334
rect 19156 27270 19208 27276
rect 19168 27130 19196 27270
rect 19260 27130 19288 27406
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19156 27124 19208 27130
rect 19156 27066 19208 27072
rect 19248 27124 19300 27130
rect 19248 27066 19300 27072
rect 20168 27124 20220 27130
rect 20168 27066 20220 27072
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18696 26988 18748 26994
rect 18696 26930 18748 26936
rect 18972 26988 19024 26994
rect 18972 26930 19024 26936
rect 18052 26852 18104 26858
rect 18052 26794 18104 26800
rect 18144 26852 18196 26858
rect 18144 26794 18196 26800
rect 18064 26518 18092 26794
rect 18708 26586 18736 26930
rect 19984 26852 20036 26858
rect 19984 26794 20036 26800
rect 19248 26784 19300 26790
rect 19248 26726 19300 26732
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 18052 26512 18104 26518
rect 18052 26454 18104 26460
rect 19260 26314 19288 26726
rect 17592 26308 17644 26314
rect 17592 26250 17644 26256
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 17788 26042 17816 26250
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 17776 26036 17828 26042
rect 17776 25978 17828 25984
rect 19996 25906 20024 26794
rect 18420 25900 18472 25906
rect 18420 25842 18472 25848
rect 19984 25900 20036 25906
rect 19984 25842 20036 25848
rect 17132 25832 17184 25838
rect 17132 25774 17184 25780
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 16396 25424 16448 25430
rect 16396 25366 16448 25372
rect 18248 25294 18276 25638
rect 18432 25430 18460 25842
rect 20180 25498 20208 27066
rect 21836 26926 21864 27406
rect 22008 27396 22060 27402
rect 22008 27338 22060 27344
rect 22020 26994 22048 27338
rect 22204 27334 22232 27406
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22008 26988 22060 26994
rect 22008 26930 22060 26936
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 21824 26920 21876 26926
rect 21824 26862 21876 26868
rect 22100 26784 22152 26790
rect 22100 26726 22152 26732
rect 22112 25974 22140 26726
rect 22204 26042 22232 26930
rect 22296 26926 22324 27270
rect 22284 26920 22336 26926
rect 22284 26862 22336 26868
rect 22388 26790 22416 27406
rect 24032 27328 24084 27334
rect 24032 27270 24084 27276
rect 24044 26994 24072 27270
rect 24032 26988 24084 26994
rect 24032 26930 24084 26936
rect 22376 26784 22428 26790
rect 22376 26726 22428 26732
rect 24136 26586 24164 27474
rect 24676 27396 24728 27402
rect 24676 27338 24728 27344
rect 24688 26926 24716 27338
rect 24872 27334 24900 28086
rect 25412 27396 25464 27402
rect 25412 27338 25464 27344
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 25424 27130 25452 27338
rect 33152 27334 33180 31758
rect 34336 31748 34388 31754
rect 34336 31690 34388 31696
rect 34348 31385 34376 31690
rect 34334 31376 34390 31385
rect 34334 31311 34390 31320
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 33324 29640 33376 29646
rect 33324 29582 33376 29588
rect 33232 27464 33284 27470
rect 33232 27406 33284 27412
rect 33140 27328 33192 27334
rect 33140 27270 33192 27276
rect 25412 27124 25464 27130
rect 25412 27066 25464 27072
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25964 26784 26016 26790
rect 25964 26726 26016 26732
rect 24124 26580 24176 26586
rect 24124 26522 24176 26528
rect 23020 26512 23072 26518
rect 23020 26454 23072 26460
rect 22836 26376 22888 26382
rect 22836 26318 22888 26324
rect 22192 26036 22244 26042
rect 22192 25978 22244 25984
rect 22100 25968 22152 25974
rect 22100 25910 22152 25916
rect 20996 25832 21048 25838
rect 20996 25774 21048 25780
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20456 25498 20484 25638
rect 21008 25498 21036 25774
rect 22112 25702 22140 25910
rect 22848 25906 22876 26318
rect 22836 25900 22888 25906
rect 22836 25842 22888 25848
rect 22848 25702 22876 25842
rect 23032 25702 23060 26454
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 23124 25838 23152 26318
rect 23480 26308 23532 26314
rect 23480 26250 23532 26256
rect 23492 26042 23520 26250
rect 23480 26036 23532 26042
rect 23480 25978 23532 25984
rect 24136 25906 24164 26522
rect 25240 26314 25268 26726
rect 24676 26308 24728 26314
rect 24676 26250 24728 26256
rect 25228 26308 25280 26314
rect 25228 26250 25280 26256
rect 24688 26042 24716 26250
rect 24676 26036 24728 26042
rect 24676 25978 24728 25984
rect 25976 25906 26004 26726
rect 24124 25900 24176 25906
rect 24124 25842 24176 25848
rect 25964 25900 26016 25906
rect 25964 25842 26016 25848
rect 23112 25832 23164 25838
rect 23112 25774 23164 25780
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 23020 25696 23072 25702
rect 23020 25638 23072 25644
rect 20168 25492 20220 25498
rect 20168 25434 20220 25440
rect 20444 25492 20496 25498
rect 20996 25492 21048 25498
rect 20496 25452 20576 25480
rect 20444 25434 20496 25440
rect 18420 25424 18472 25430
rect 18420 25366 18472 25372
rect 18604 25424 18656 25430
rect 18604 25366 18656 25372
rect 16212 25288 16264 25294
rect 16212 25230 16264 25236
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 16224 24818 16252 25230
rect 17592 25220 17644 25226
rect 17592 25162 17644 25168
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16120 24744 16172 24750
rect 16120 24686 16172 24692
rect 16120 24608 16172 24614
rect 16120 24550 16172 24556
rect 16132 24410 16160 24550
rect 17604 24410 17632 25162
rect 18512 24608 18564 24614
rect 18512 24550 18564 24556
rect 18524 24410 18552 24550
rect 18616 24410 18644 25366
rect 20548 25294 20576 25452
rect 20996 25434 21048 25440
rect 20904 25356 20956 25362
rect 20904 25298 20956 25304
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 20536 25288 20588 25294
rect 20812 25288 20864 25294
rect 20536 25230 20588 25236
rect 20732 25248 20812 25276
rect 19352 24954 19380 25230
rect 19432 25220 19484 25226
rect 19432 25162 19484 25168
rect 19984 25220 20036 25226
rect 19984 25162 20036 25168
rect 19340 24948 19392 24954
rect 19340 24890 19392 24896
rect 19444 24886 19472 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19432 24880 19484 24886
rect 19484 24828 19840 24834
rect 19432 24822 19840 24828
rect 19340 24812 19392 24818
rect 19444 24806 19840 24822
rect 19340 24754 19392 24760
rect 16120 24404 16172 24410
rect 16120 24346 16172 24352
rect 17592 24404 17644 24410
rect 17592 24346 17644 24352
rect 18512 24404 18564 24410
rect 18512 24346 18564 24352
rect 18604 24404 18656 24410
rect 18604 24346 18656 24352
rect 15660 24336 15712 24342
rect 15660 24278 15712 24284
rect 16764 24268 16816 24274
rect 16764 24210 16816 24216
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15108 22568 15160 22574
rect 15108 22510 15160 22516
rect 15120 22438 15148 22510
rect 15108 22432 15160 22438
rect 15108 22374 15160 22380
rect 15200 22432 15252 22438
rect 15200 22374 15252 22380
rect 14740 22024 14792 22030
rect 14740 21966 14792 21972
rect 14924 22024 14976 22030
rect 14924 21966 14976 21972
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 14556 21956 14608 21962
rect 14556 21898 14608 21904
rect 14648 21956 14700 21962
rect 14648 21898 14700 21904
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13832 21622 13860 21830
rect 14568 21690 14596 21898
rect 14556 21684 14608 21690
rect 14556 21626 14608 21632
rect 13820 21616 13872 21622
rect 13872 21576 14136 21604
rect 13820 21558 13872 21564
rect 13820 21480 13872 21486
rect 13648 21428 13820 21434
rect 13648 21422 13872 21428
rect 13648 21406 13860 21422
rect 13544 21140 13596 21146
rect 13544 21082 13596 21088
rect 13544 20936 13596 20942
rect 13648 20890 13676 21406
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13912 21344 13964 21350
rect 13912 21286 13964 21292
rect 13596 20884 13676 20890
rect 13544 20878 13676 20884
rect 13556 20862 13676 20878
rect 13740 20874 13768 21286
rect 13924 21146 13952 21286
rect 13912 21140 13964 21146
rect 13912 21082 13964 21088
rect 13360 20800 13412 20806
rect 13360 20742 13412 20748
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12808 20460 12860 20466
rect 12728 20420 12808 20448
rect 12808 20402 12860 20408
rect 12716 20052 12768 20058
rect 12716 19994 12768 20000
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12636 19446 12664 19790
rect 12624 19440 12676 19446
rect 12624 19382 12676 19388
rect 12728 19378 12756 19994
rect 12820 19922 12848 20402
rect 12808 19916 12860 19922
rect 12808 19858 12860 19864
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12532 19236 12584 19242
rect 12532 19178 12584 19184
rect 12624 18624 12676 18630
rect 12624 18566 12676 18572
rect 12636 18290 12664 18566
rect 12912 18306 12940 20470
rect 13372 20262 13400 20742
rect 13360 20256 13412 20262
rect 13360 20198 13412 20204
rect 13268 19984 13320 19990
rect 13268 19926 13320 19932
rect 13280 19242 13308 19926
rect 13268 19236 13320 19242
rect 13268 19178 13320 19184
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 13004 18426 13032 18566
rect 12992 18420 13044 18426
rect 12992 18362 13044 18368
rect 12624 18284 12676 18290
rect 12912 18278 13032 18306
rect 12624 18226 12676 18232
rect 12636 18154 12664 18226
rect 12624 18148 12676 18154
rect 12624 18090 12676 18096
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12268 17270 12296 17478
rect 12256 17264 12308 17270
rect 12256 17206 12308 17212
rect 12452 17134 12480 17478
rect 12544 17270 12572 17546
rect 12532 17264 12584 17270
rect 12532 17206 12584 17212
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12268 16946 12296 17070
rect 12268 16918 12572 16946
rect 12544 16658 12572 16918
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12256 16584 12308 16590
rect 12256 16526 12308 16532
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12162 16144 12218 16153
rect 12162 16079 12164 16088
rect 12216 16079 12218 16088
rect 12164 16050 12216 16056
rect 12268 16046 12296 16526
rect 12532 16516 12584 16522
rect 12532 16458 12584 16464
rect 12256 16040 12308 16046
rect 12256 15982 12308 15988
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12348 15904 12400 15910
rect 12348 15846 12400 15852
rect 12084 15638 12112 15846
rect 12072 15632 12124 15638
rect 12072 15574 12124 15580
rect 11980 14884 12032 14890
rect 11980 14826 12032 14832
rect 11992 14414 12020 14826
rect 12084 14482 12112 15574
rect 12360 15502 12388 15846
rect 12348 15496 12400 15502
rect 12348 15438 12400 15444
rect 12544 15162 12572 16458
rect 12636 15178 12664 16526
rect 12728 16114 12756 16730
rect 12716 16108 12768 16114
rect 12716 16050 12768 16056
rect 12728 15638 12756 16050
rect 12716 15632 12768 15638
rect 12716 15574 12768 15580
rect 12820 15366 12848 16730
rect 12900 16584 12952 16590
rect 12900 16526 12952 16532
rect 12912 15502 12940 16526
rect 13004 16289 13032 18278
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 13188 17338 13216 17750
rect 13176 17332 13228 17338
rect 13176 17274 13228 17280
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12990 16280 13046 16289
rect 12990 16215 13046 16224
rect 12990 16144 13046 16153
rect 12990 16079 12992 16088
rect 13044 16079 13046 16088
rect 12992 16050 13044 16056
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 13004 15638 13032 15914
rect 12992 15632 13044 15638
rect 12992 15574 13044 15580
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 12808 15360 12860 15366
rect 12808 15302 12860 15308
rect 13004 15178 13032 15438
rect 13096 15366 13124 17138
rect 13280 17134 13308 18226
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13372 16590 13400 20198
rect 13648 19922 13676 20862
rect 13728 20868 13780 20874
rect 13728 20810 13780 20816
rect 14004 20800 14056 20806
rect 14002 20768 14004 20777
rect 14056 20768 14058 20777
rect 14002 20703 14058 20712
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 14108 19854 14136 21576
rect 14188 21548 14240 21554
rect 14188 21490 14240 21496
rect 14200 20942 14228 21490
rect 14372 21480 14424 21486
rect 14372 21422 14424 21428
rect 14384 21146 14412 21422
rect 14568 21146 14596 21626
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14556 21140 14608 21146
rect 14556 21082 14608 21088
rect 14188 20936 14240 20942
rect 14188 20878 14240 20884
rect 14752 19961 14780 21966
rect 14936 21010 14964 21966
rect 15028 21146 15056 21966
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 14924 21004 14976 21010
rect 14924 20946 14976 20952
rect 14936 20602 14964 20946
rect 14924 20596 14976 20602
rect 14924 20538 14976 20544
rect 15120 20534 15148 21966
rect 15212 21434 15240 22374
rect 15304 22234 15332 23122
rect 15856 22982 15884 23258
rect 16672 23180 16724 23186
rect 16672 23122 16724 23128
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 15844 22976 15896 22982
rect 15844 22918 15896 22924
rect 16040 22778 16068 23054
rect 16028 22772 16080 22778
rect 16028 22714 16080 22720
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15476 22636 15528 22642
rect 15476 22578 15528 22584
rect 15292 22228 15344 22234
rect 15292 22170 15344 22176
rect 15396 21554 15424 22578
rect 15488 22030 15516 22578
rect 15844 22568 15896 22574
rect 15844 22510 15896 22516
rect 15856 22094 15884 22510
rect 15856 22066 16068 22094
rect 15476 22024 15528 22030
rect 15476 21966 15528 21972
rect 15936 21888 15988 21894
rect 15936 21830 15988 21836
rect 15948 21554 15976 21830
rect 15384 21548 15436 21554
rect 15384 21490 15436 21496
rect 15568 21548 15620 21554
rect 15568 21490 15620 21496
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 15212 21406 15424 21434
rect 15396 21010 15424 21406
rect 15580 21146 15608 21490
rect 15660 21480 15712 21486
rect 15660 21422 15712 21428
rect 15568 21140 15620 21146
rect 15568 21082 15620 21088
rect 15384 21004 15436 21010
rect 15384 20946 15436 20952
rect 15672 20942 15700 21422
rect 16040 21010 16068 22066
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16224 21690 16252 21830
rect 16408 21690 16436 21966
rect 16684 21690 16712 23122
rect 16212 21684 16264 21690
rect 16212 21626 16264 21632
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16672 21684 16724 21690
rect 16672 21626 16724 21632
rect 16028 21004 16080 21010
rect 16028 20946 16080 20952
rect 15660 20936 15712 20942
rect 15660 20878 15712 20884
rect 15108 20528 15160 20534
rect 15108 20470 15160 20476
rect 15672 20466 15700 20878
rect 16040 20466 16068 20946
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 14738 19952 14794 19961
rect 14738 19887 14794 19896
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13556 19378 13584 19654
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13464 17338 13492 19110
rect 13452 17332 13504 17338
rect 13452 17274 13504 17280
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16794 13492 16934
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13188 15706 13216 16458
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16114 13400 16390
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13176 15700 13228 15706
rect 13176 15642 13228 15648
rect 13280 15570 13308 15846
rect 13372 15638 13400 16050
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 13556 15502 13584 19178
rect 14740 18828 14792 18834
rect 14740 18770 14792 18776
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 13648 16402 13676 18566
rect 14476 18426 14504 18566
rect 14568 18426 14596 18566
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14752 18290 14780 18770
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 14464 18284 14516 18290
rect 14464 18226 14516 18232
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 14476 18136 14504 18226
rect 14556 18148 14608 18154
rect 14476 18108 14556 18136
rect 13820 18080 13872 18086
rect 14292 18034 14320 18090
rect 13872 18028 14320 18034
rect 13820 18022 14320 18028
rect 13832 18006 14320 18022
rect 14476 17678 14504 18108
rect 14556 18090 14608 18096
rect 14752 17678 14780 18226
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14648 17672 14700 17678
rect 14648 17614 14700 17620
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 16794 13768 16934
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13728 16584 13780 16590
rect 14188 16584 14240 16590
rect 13780 16544 14188 16572
rect 13728 16526 13780 16532
rect 14188 16526 14240 16532
rect 13648 16374 13768 16402
rect 13634 16280 13690 16289
rect 13634 16215 13690 16224
rect 13544 15496 13596 15502
rect 13544 15438 13596 15444
rect 13084 15360 13136 15366
rect 13648 15314 13676 16215
rect 13740 15434 13768 16374
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13084 15302 13136 15308
rect 12532 15156 12584 15162
rect 12636 15150 13032 15178
rect 12532 15098 12584 15104
rect 12164 15020 12216 15026
rect 12164 14962 12216 14968
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 11980 14408 12032 14414
rect 11980 14350 12032 14356
rect 11980 13728 12032 13734
rect 11980 13670 12032 13676
rect 11992 13326 12020 13670
rect 12084 13530 12112 14418
rect 12176 14414 12204 14962
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12360 14414 12388 14554
rect 12544 14414 12572 15098
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12728 14929 12756 14962
rect 12714 14920 12770 14929
rect 12714 14855 12770 14864
rect 12900 14884 12952 14890
rect 12728 14482 12756 14855
rect 12900 14826 12952 14832
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12912 14414 12940 14826
rect 12164 14408 12216 14414
rect 12162 14376 12164 14385
rect 12348 14408 12400 14414
rect 12216 14376 12218 14385
rect 12348 14350 12400 14356
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 12900 14408 12952 14414
rect 13004 14385 13032 15150
rect 13464 15286 13676 15314
rect 13464 14958 13492 15286
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 12900 14350 12952 14356
rect 12990 14376 13046 14385
rect 12162 14311 12218 14320
rect 12808 14340 12860 14346
rect 12990 14311 13046 14320
rect 12808 14282 12860 14288
rect 12256 14272 12308 14278
rect 12256 14214 12308 14220
rect 12532 14272 12584 14278
rect 12532 14214 12584 14220
rect 12268 14074 12296 14214
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12360 13462 12388 13670
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 11980 13320 12032 13326
rect 11980 13262 12032 13268
rect 11992 12986 12020 13262
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12176 12442 12204 12582
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 11900 12238 11928 12378
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 11336 12232 11388 12238
rect 11520 12232 11572 12238
rect 11336 12174 11388 12180
rect 11518 12200 11520 12209
rect 11888 12232 11940 12238
rect 11572 12200 11574 12209
rect 10232 12164 10284 12170
rect 11888 12174 11940 12180
rect 11518 12135 11574 12144
rect 10232 12106 10284 12112
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11898 11652 12038
rect 11900 11898 11928 12174
rect 12360 12102 12388 13398
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12176 11898 12204 12038
rect 11612 11892 11664 11898
rect 11612 11834 11664 11840
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11900 11694 11928 11834
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 12176 11354 12204 11834
rect 12164 11348 12216 11354
rect 12164 11290 12216 11296
rect 12360 11082 12388 12038
rect 12452 11898 12480 12582
rect 12544 12238 12572 14214
rect 12716 13796 12768 13802
rect 12716 13738 12768 13744
rect 12728 13530 12756 13738
rect 12820 13530 12848 14282
rect 13096 14260 13124 14554
rect 13464 14482 13492 14894
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13556 14482 13584 14758
rect 13452 14476 13504 14482
rect 13452 14418 13504 14424
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13740 14414 13768 15370
rect 13832 15162 13860 15506
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 14476 14550 14504 17614
rect 14556 17604 14608 17610
rect 14556 17546 14608 17552
rect 14568 17066 14596 17546
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14568 16590 14596 17002
rect 14660 16794 14688 17614
rect 14844 17542 14872 18226
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 17338 14872 17478
rect 14832 17332 14884 17338
rect 14832 17274 14884 17280
rect 14648 16788 14700 16794
rect 14648 16730 14700 16736
rect 14844 16697 14872 17274
rect 15120 17202 15148 18226
rect 15212 17746 15240 18362
rect 15304 17882 15332 18702
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15200 17740 15252 17746
rect 15200 17682 15252 17688
rect 15200 17604 15252 17610
rect 15200 17546 15252 17552
rect 15212 17338 15240 17546
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 14924 17196 14976 17202
rect 14924 17138 14976 17144
rect 15108 17196 15160 17202
rect 15108 17138 15160 17144
rect 14830 16688 14886 16697
rect 14830 16623 14886 16632
rect 14844 16590 14872 16623
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14832 16584 14884 16590
rect 14832 16526 14884 16532
rect 14648 16448 14700 16454
rect 14648 16390 14700 16396
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14464 14544 14516 14550
rect 14464 14486 14516 14492
rect 13636 14408 13688 14414
rect 13634 14376 13636 14385
rect 13728 14408 13780 14414
rect 13688 14376 13690 14385
rect 13360 14340 13412 14346
rect 13728 14350 13780 14356
rect 13634 14311 13690 14320
rect 13820 14340 13872 14346
rect 13360 14282 13412 14288
rect 13820 14282 13872 14288
rect 13004 14232 13124 14260
rect 13176 14272 13228 14278
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12624 13524 12676 13530
rect 12624 13466 12676 13472
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12636 13394 12664 13466
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12808 13388 12860 13394
rect 12808 13330 12860 13336
rect 12820 12918 12848 13330
rect 12912 12986 12940 13670
rect 13004 13326 13032 14232
rect 13176 14214 13228 14220
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 13096 13870 13124 13942
rect 13188 13938 13216 14214
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13372 13802 13400 14282
rect 13832 14249 13860 14282
rect 13818 14240 13874 14249
rect 13818 14175 13874 14184
rect 13452 14068 13504 14074
rect 13504 14028 13768 14056
rect 13452 14010 13504 14016
rect 13450 13968 13506 13977
rect 13740 13938 13768 14028
rect 14568 14006 14596 14554
rect 14660 14521 14688 16390
rect 14844 16250 14872 16526
rect 14832 16244 14884 16250
rect 14832 16186 14884 16192
rect 14936 15026 14964 17138
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15120 15570 15148 16526
rect 15396 16250 15424 19314
rect 16592 18426 16620 19314
rect 16684 18766 16712 19722
rect 16776 19242 16804 24210
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16868 23322 16896 24142
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 16856 23316 16908 23322
rect 16856 23258 16908 23264
rect 17132 22976 17184 22982
rect 17132 22918 17184 22924
rect 17144 22778 17172 22918
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17224 22568 17276 22574
rect 17224 22510 17276 22516
rect 16856 21548 16908 21554
rect 16856 21490 16908 21496
rect 16868 21146 16896 21490
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 16960 19242 16988 19926
rect 17040 19712 17092 19718
rect 17040 19654 17092 19660
rect 17052 19514 17080 19654
rect 17040 19508 17092 19514
rect 17040 19450 17092 19456
rect 17132 19304 17184 19310
rect 17132 19246 17184 19252
rect 16764 19236 16816 19242
rect 16764 19178 16816 19184
rect 16948 19236 17000 19242
rect 16948 19178 17000 19184
rect 16960 18834 16988 19178
rect 17144 18970 17172 19246
rect 17236 18970 17264 22510
rect 18156 22234 18184 24006
rect 19352 22778 19380 24754
rect 19812 24750 19840 24806
rect 19800 24744 19852 24750
rect 19800 24686 19852 24692
rect 19996 24682 20024 25162
rect 20364 25140 20392 25230
rect 20732 25140 20760 25248
rect 20812 25230 20864 25236
rect 20364 25112 20760 25140
rect 20812 25152 20864 25158
rect 20812 25094 20864 25100
rect 19984 24676 20036 24682
rect 19984 24618 20036 24624
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 20824 23866 20852 25094
rect 20916 24750 20944 25298
rect 20996 25288 21048 25294
rect 20996 25230 21048 25236
rect 21008 24954 21036 25230
rect 20996 24948 21048 24954
rect 20996 24890 21048 24896
rect 20904 24744 20956 24750
rect 20904 24686 20956 24692
rect 20812 23860 20864 23866
rect 20812 23802 20864 23808
rect 20628 23724 20680 23730
rect 20628 23666 20680 23672
rect 21088 23724 21140 23730
rect 21088 23666 21140 23672
rect 20444 23656 20496 23662
rect 20444 23598 20496 23604
rect 20456 23322 20484 23598
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19444 22778 19472 23122
rect 20456 23118 20484 23258
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19340 22772 19392 22778
rect 19340 22714 19392 22720
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19996 22642 20024 23054
rect 20640 23050 20668 23666
rect 21100 23254 21128 23666
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 21916 23656 21968 23662
rect 21916 23598 21968 23604
rect 21180 23588 21232 23594
rect 21180 23530 21232 23536
rect 21088 23248 21140 23254
rect 21088 23190 21140 23196
rect 21192 23186 21220 23530
rect 21180 23180 21232 23186
rect 21180 23122 21232 23128
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20720 22976 20772 22982
rect 20720 22918 20772 22924
rect 19984 22636 20036 22642
rect 19984 22578 20036 22584
rect 18328 22568 18380 22574
rect 18328 22510 18380 22516
rect 18788 22568 18840 22574
rect 18788 22510 18840 22516
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18248 22030 18276 22374
rect 18340 22030 18368 22510
rect 18800 22094 18828 22510
rect 19996 22234 20024 22578
rect 19984 22228 20036 22234
rect 19984 22170 20036 22176
rect 18800 22066 18920 22094
rect 18892 22030 18920 22066
rect 18236 22024 18288 22030
rect 18236 21966 18288 21972
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 17408 21888 17460 21894
rect 17408 21830 17460 21836
rect 17420 21690 17448 21830
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17420 21418 17448 21626
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 17604 21486 17632 21558
rect 17592 21480 17644 21486
rect 17592 21422 17644 21428
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 18144 21344 18196 21350
rect 18144 21286 18196 21292
rect 18236 21344 18288 21350
rect 18236 21286 18288 21292
rect 18156 20942 18184 21286
rect 18248 21146 18276 21286
rect 18236 21140 18288 21146
rect 18236 21082 18288 21088
rect 17684 20936 17736 20942
rect 17684 20878 17736 20884
rect 18144 20936 18196 20942
rect 18144 20878 18196 20884
rect 17696 20398 17724 20878
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17972 20398 18000 20742
rect 18156 20398 18184 20878
rect 18248 20602 18276 21082
rect 18892 20602 18920 21966
rect 19996 21894 20024 22170
rect 20168 22160 20220 22166
rect 20168 22102 20220 22108
rect 20180 22030 20208 22102
rect 20168 22024 20220 22030
rect 20168 21966 20220 21972
rect 19984 21888 20036 21894
rect 19984 21830 20036 21836
rect 20536 21888 20588 21894
rect 20536 21830 20588 21836
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21146 20024 21830
rect 20548 21146 20576 21830
rect 20732 21554 20760 22918
rect 21468 22234 21496 23598
rect 21928 23322 21956 23598
rect 21916 23316 21968 23322
rect 21916 23258 21968 23264
rect 22112 23118 22140 25638
rect 23032 25430 23060 25638
rect 23020 25424 23072 25430
rect 23020 25366 23072 25372
rect 23124 25294 23152 25774
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23124 23798 23152 25230
rect 23676 23866 23704 25230
rect 24136 24410 24164 25842
rect 33244 25838 33272 27406
rect 33336 26450 33364 29582
rect 34888 29572 34940 29578
rect 34888 29514 34940 29520
rect 34900 29209 34928 29514
rect 34886 29200 34942 29209
rect 34886 29135 34942 29144
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34888 27396 34940 27402
rect 34888 27338 34940 27344
rect 34900 27033 34928 27338
rect 34886 27024 34942 27033
rect 34886 26959 34942 26968
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 33324 26444 33376 26450
rect 33324 26386 33376 26392
rect 24400 25832 24452 25838
rect 24400 25774 24452 25780
rect 33232 25832 33284 25838
rect 33232 25774 33284 25780
rect 24412 25498 24440 25774
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 24400 25492 24452 25498
rect 24400 25434 24452 25440
rect 24124 24404 24176 24410
rect 24124 24346 24176 24352
rect 23664 23860 23716 23866
rect 23664 23802 23716 23808
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23020 23724 23072 23730
rect 23020 23666 23072 23672
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23032 23526 23060 23666
rect 23020 23520 23072 23526
rect 23020 23462 23072 23468
rect 23032 23322 23060 23462
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 22100 23112 22152 23118
rect 22100 23054 22152 23060
rect 22652 23112 22704 23118
rect 22652 23054 22704 23060
rect 22560 22636 22612 22642
rect 22560 22578 22612 22584
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21088 22160 21140 22166
rect 21088 22102 21140 22108
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 21008 21690 21036 21830
rect 21100 21690 21128 22102
rect 21732 22092 21784 22098
rect 21732 22034 21784 22040
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 21088 21684 21140 21690
rect 21088 21626 21140 21632
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 19984 21004 20036 21010
rect 19984 20946 20036 20952
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19248 20868 19300 20874
rect 19248 20810 19300 20816
rect 19156 20800 19208 20806
rect 19156 20742 19208 20748
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18880 20596 18932 20602
rect 18880 20538 18932 20544
rect 19168 20534 19196 20742
rect 19156 20528 19208 20534
rect 19156 20470 19208 20476
rect 19260 20398 19288 20810
rect 19444 20602 19472 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 20946
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19444 20448 19472 20538
rect 19524 20460 19576 20466
rect 19444 20420 19524 20448
rect 19524 20402 19576 20408
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 18144 20392 18196 20398
rect 18144 20334 18196 20340
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17132 18964 17184 18970
rect 17132 18906 17184 18912
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17604 18902 17632 19382
rect 17696 18970 17724 20334
rect 17972 19514 18000 20334
rect 18236 20324 18288 20330
rect 18236 20266 18288 20272
rect 18052 19848 18104 19854
rect 18052 19790 18104 19796
rect 17960 19508 18012 19514
rect 17960 19450 18012 19456
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 17592 18896 17644 18902
rect 17592 18838 17644 18844
rect 16948 18828 17000 18834
rect 16948 18770 17000 18776
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16580 18420 16632 18426
rect 16580 18362 16632 18368
rect 15568 18284 15620 18290
rect 15568 18226 15620 18232
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15580 17678 15608 18226
rect 15672 17678 15700 18226
rect 16684 17814 16712 18702
rect 17788 18698 17816 19110
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 17880 18426 17908 18702
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 16672 17808 16724 17814
rect 16672 17750 16724 17756
rect 18064 17678 18092 19790
rect 18248 19786 18276 20266
rect 18236 19780 18288 19786
rect 18236 19722 18288 19728
rect 18972 19780 19024 19786
rect 18972 19722 19024 19728
rect 18248 19378 18276 19722
rect 18236 19372 18288 19378
rect 18236 19314 18288 19320
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18524 18154 18552 19314
rect 18984 19310 19012 19722
rect 19432 19712 19484 19718
rect 19432 19654 19484 19660
rect 19444 19378 19472 19654
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19996 19514 20024 20402
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18970 19380 19110
rect 19340 18964 19392 18970
rect 19340 18906 19392 18912
rect 19720 18766 19748 19314
rect 19340 18760 19392 18766
rect 19340 18702 19392 18708
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 18512 18148 18564 18154
rect 18512 18090 18564 18096
rect 19352 17882 19380 18702
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 20088 17882 20116 20878
rect 21008 18902 21036 21490
rect 21284 21486 21312 21966
rect 21744 21690 21772 22034
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 21732 21684 21784 21690
rect 21732 21626 21784 21632
rect 22480 21622 22508 21830
rect 22572 21622 22600 22578
rect 22468 21616 22520 21622
rect 22468 21558 22520 21564
rect 22560 21616 22612 21622
rect 22560 21558 22612 21564
rect 21272 21480 21324 21486
rect 21272 21422 21324 21428
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 20720 18828 20772 18834
rect 20720 18770 20772 18776
rect 19340 17876 19392 17882
rect 19340 17818 19392 17824
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20444 17808 20496 17814
rect 20444 17750 20496 17756
rect 20456 17678 20484 17750
rect 20732 17678 20760 18770
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20824 17882 20852 18702
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20996 17808 21048 17814
rect 20996 17750 21048 17756
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15660 17672 15712 17678
rect 18052 17672 18104 17678
rect 15660 17614 15712 17620
rect 17972 17620 18052 17626
rect 17972 17614 18104 17620
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 17972 17598 18092 17614
rect 17972 17202 18000 17598
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18064 17134 18092 17478
rect 18616 17202 18644 17478
rect 18892 17270 18920 17614
rect 20168 17536 20220 17542
rect 20168 17478 20220 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18052 17128 18104 17134
rect 18052 17070 18104 17076
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 19340 16992 19392 16998
rect 19340 16934 19392 16940
rect 15672 16794 15700 16934
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 15488 16522 15516 16662
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16304 16584 16356 16590
rect 16304 16526 16356 16532
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15384 16244 15436 16250
rect 15384 16186 15436 16192
rect 16316 15910 16344 16526
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 14924 15020 14976 15026
rect 14924 14962 14976 14968
rect 14646 14512 14702 14521
rect 14646 14447 14702 14456
rect 14660 14414 14688 14447
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14556 14000 14608 14006
rect 14370 13968 14426 13977
rect 13450 13903 13452 13912
rect 13504 13903 13506 13912
rect 13728 13932 13780 13938
rect 13452 13874 13504 13880
rect 13728 13874 13780 13880
rect 14096 13932 14148 13938
rect 14556 13942 14608 13948
rect 15120 13938 15148 15506
rect 15304 14958 15332 15642
rect 15672 15502 15700 15846
rect 16408 15638 16436 16594
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18800 16250 18828 16526
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16500 15638 16528 15914
rect 16592 15706 16620 16186
rect 16764 15904 16816 15910
rect 16764 15846 16816 15852
rect 16776 15706 16804 15846
rect 16580 15700 16632 15706
rect 16764 15700 16816 15706
rect 16632 15660 16712 15688
rect 16580 15642 16632 15648
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16488 15632 16540 15638
rect 16488 15574 16540 15580
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15396 15026 15424 15438
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15304 14074 15332 14350
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15672 13938 15700 14758
rect 16408 14550 16436 15574
rect 16580 15360 16632 15366
rect 16580 15302 16632 15308
rect 16592 15162 16620 15302
rect 16684 15162 16712 15660
rect 16764 15642 16816 15648
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16672 15156 16724 15162
rect 16672 15098 16724 15104
rect 16776 14958 16804 15302
rect 16764 14952 16816 14958
rect 16764 14894 16816 14900
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 18064 14618 18092 14894
rect 18236 14816 18288 14822
rect 18236 14758 18288 14764
rect 18248 14618 18276 14758
rect 18052 14612 18104 14618
rect 18052 14554 18104 14560
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15764 14074 15792 14214
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 14370 13903 14372 13912
rect 14096 13874 14148 13880
rect 14424 13903 14426 13912
rect 15108 13932 15160 13938
rect 14372 13874 14424 13880
rect 15108 13874 15160 13880
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 14108 13802 14136 13874
rect 13360 13796 13412 13802
rect 13360 13738 13412 13744
rect 14096 13796 14148 13802
rect 14096 13738 14148 13744
rect 13912 13728 13964 13734
rect 13912 13670 13964 13676
rect 14924 13728 14976 13734
rect 14924 13670 14976 13676
rect 13728 13456 13780 13462
rect 13728 13398 13780 13404
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 13556 12646 13584 13126
rect 13740 12646 13768 13398
rect 13924 12850 13952 13670
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 12986 14044 13126
rect 14108 12986 14136 13262
rect 14936 12986 14964 13670
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 16040 12918 16068 13126
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 13912 12844 13964 12850
rect 14372 12844 14424 12850
rect 13964 12804 14228 12832
rect 13912 12786 13964 12792
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13728 12640 13780 12646
rect 13728 12582 13780 12588
rect 13556 12238 13584 12582
rect 13740 12306 13768 12582
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 14200 12238 14228 12804
rect 14372 12786 14424 12792
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14384 12238 14412 12786
rect 14568 12434 14596 12786
rect 14936 12442 14964 12786
rect 16132 12714 16160 14350
rect 18800 14346 18828 16186
rect 19260 16182 19288 16662
rect 19352 16658 19380 16934
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19248 16176 19300 16182
rect 19248 16118 19300 16124
rect 19444 15162 19472 16526
rect 20180 16522 20208 17478
rect 20640 17134 20668 17614
rect 20916 17202 20944 17614
rect 21008 17202 21036 17750
rect 22008 17740 22060 17746
rect 22008 17682 22060 17688
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21180 17536 21232 17542
rect 21180 17478 21232 17484
rect 21192 17270 21220 17478
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20904 17196 20956 17202
rect 20904 17138 20956 17144
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 20628 17128 20680 17134
rect 20628 17070 20680 17076
rect 20640 16590 20668 17070
rect 20824 16794 20852 17138
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20916 16590 20944 17138
rect 21008 16590 21036 17138
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21192 16794 21220 16934
rect 21180 16788 21232 16794
rect 21180 16730 21232 16736
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19996 16250 20024 16390
rect 19984 16244 20036 16250
rect 19984 16186 20036 16192
rect 20260 16244 20312 16250
rect 20260 16186 20312 16192
rect 20272 16114 20300 16186
rect 20076 16108 20128 16114
rect 20260 16108 20312 16114
rect 20128 16068 20260 16096
rect 20076 16050 20128 16056
rect 20260 16050 20312 16056
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 18972 14952 19024 14958
rect 18972 14894 19024 14900
rect 18788 14340 18840 14346
rect 18788 14282 18840 14288
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 18880 14272 18932 14278
rect 18880 14214 18932 14220
rect 16304 13728 16356 13734
rect 16304 13670 16356 13676
rect 16120 12708 16172 12714
rect 16120 12650 16172 12656
rect 15752 12640 15804 12646
rect 15752 12582 15804 12588
rect 14476 12406 14596 12434
rect 14924 12436 14976 12442
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 14200 11830 14228 12174
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14384 11762 14412 12174
rect 14476 12102 14504 12406
rect 14924 12378 14976 12384
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14476 11558 14504 12038
rect 15672 11898 15700 12038
rect 15764 11898 15792 12582
rect 16316 12209 16344 13670
rect 17052 13326 17080 14214
rect 18892 14074 18920 14214
rect 18984 14074 19012 14894
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 19260 14006 19288 15030
rect 19352 14822 19380 15098
rect 19340 14816 19392 14822
rect 19340 14758 19392 14764
rect 19352 14618 19380 14758
rect 19996 14618 20024 15302
rect 20088 14958 20116 16050
rect 20456 15570 20484 16050
rect 20444 15564 20496 15570
rect 20444 15506 20496 15512
rect 20548 15502 20576 16050
rect 20916 15978 20944 16526
rect 21008 16232 21036 16526
rect 21284 16522 21312 17614
rect 22020 17338 22048 17682
rect 22008 17332 22060 17338
rect 22008 17274 22060 17280
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21088 16244 21140 16250
rect 21008 16204 21088 16232
rect 21088 16186 21140 16192
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 20904 15972 20956 15978
rect 20904 15914 20956 15920
rect 22020 15706 22048 16050
rect 22480 15706 22508 16050
rect 22008 15700 22060 15706
rect 22008 15642 22060 15648
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 20720 15564 20772 15570
rect 20720 15506 20772 15512
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20076 14952 20128 14958
rect 20076 14894 20128 14900
rect 20352 14884 20404 14890
rect 20352 14826 20404 14832
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 18880 13932 18932 13938
rect 18880 13874 18932 13880
rect 17972 13530 18000 13874
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 17960 13320 18012 13326
rect 17960 13262 18012 13268
rect 17052 12986 17080 13262
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17132 12912 17184 12918
rect 17132 12854 17184 12860
rect 16672 12844 16724 12850
rect 16948 12844 17000 12850
rect 16724 12804 16804 12832
rect 16672 12786 16724 12792
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16592 12442 16620 12718
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 16302 12200 16358 12209
rect 16302 12135 16358 12144
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16132 11898 16160 12038
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16316 11762 16344 12135
rect 16684 11762 16712 12582
rect 16776 12170 16804 12804
rect 16948 12786 17000 12792
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16960 12170 16988 12786
rect 17052 12442 17080 12786
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17144 12238 17172 12854
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17512 12238 17540 12786
rect 17880 12782 17908 13126
rect 17972 12782 18000 13262
rect 18064 12986 18092 13806
rect 18892 13462 18920 13874
rect 19352 13734 19380 14350
rect 19444 13870 19472 14418
rect 20364 14414 20392 14826
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 13728 19392 13734
rect 19340 13670 19392 13676
rect 19352 13530 19380 13670
rect 19444 13530 19472 13806
rect 19340 13524 19392 13530
rect 19340 13466 19392 13472
rect 19432 13524 19484 13530
rect 19432 13466 19484 13472
rect 18880 13456 18932 13462
rect 18880 13398 18932 13404
rect 19628 13326 19656 13874
rect 19996 13530 20024 14214
rect 20272 14074 20300 14350
rect 20456 14074 20484 14758
rect 20732 14550 20760 15506
rect 20996 14884 21048 14890
rect 20996 14826 21048 14832
rect 20720 14544 20772 14550
rect 20720 14486 20772 14492
rect 20732 14278 20760 14486
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20824 14346 20852 14418
rect 21008 14414 21036 14826
rect 22480 14618 22508 15642
rect 22468 14612 22520 14618
rect 22468 14554 22520 14560
rect 22560 14476 22612 14482
rect 22560 14418 22612 14424
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 22468 14408 22520 14414
rect 22468 14350 22520 14356
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20720 14272 20772 14278
rect 20720 14214 20772 14220
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 14074 21312 14214
rect 22480 14074 22508 14350
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22572 13938 22600 14418
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 21732 13796 21784 13802
rect 21732 13738 21784 13744
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 21468 13326 21496 13670
rect 21744 13326 21772 13738
rect 22572 13530 22600 13874
rect 22664 13530 22692 23054
rect 23032 22778 23060 23258
rect 23400 22778 23428 23666
rect 24136 22778 24164 24346
rect 24676 24132 24728 24138
rect 24676 24074 24728 24080
rect 24952 24132 25004 24138
rect 24952 24074 25004 24080
rect 24688 23866 24716 24074
rect 24964 23866 24992 24074
rect 24676 23860 24728 23866
rect 24676 23802 24728 23808
rect 24952 23860 25004 23866
rect 24952 23802 25004 23808
rect 25516 23526 25544 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 33140 25288 33192 25294
rect 33140 25230 33192 25236
rect 33152 24070 33180 25230
rect 34336 25220 34388 25226
rect 34336 25162 34388 25168
rect 34348 24857 34376 25162
rect 34334 24848 34390 24857
rect 34334 24783 34390 24792
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 33140 24064 33192 24070
rect 33140 24006 33192 24012
rect 25504 23520 25556 23526
rect 25504 23462 25556 23468
rect 23020 22772 23072 22778
rect 23020 22714 23072 22720
rect 23388 22772 23440 22778
rect 23388 22714 23440 22720
rect 24124 22772 24176 22778
rect 24124 22714 24176 22720
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 22940 22166 22968 22578
rect 22928 22160 22980 22166
rect 22928 22102 22980 22108
rect 23216 22030 23244 22578
rect 23204 22024 23256 22030
rect 23204 21966 23256 21972
rect 23216 21690 23244 21966
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 23296 21548 23348 21554
rect 23296 21490 23348 21496
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 23204 21344 23256 21350
rect 23204 21286 23256 21292
rect 22848 21146 22876 21286
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 23216 20806 23244 21286
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 23216 17882 23244 20742
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23308 17610 23336 21490
rect 24136 21146 24164 22714
rect 25516 22642 25544 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 33152 22778 33180 23054
rect 34888 23044 34940 23050
rect 34888 22986 34940 22992
rect 33140 22772 33192 22778
rect 33140 22714 33192 22720
rect 34900 22681 34928 22986
rect 34886 22672 34942 22681
rect 25504 22636 25556 22642
rect 34886 22607 34942 22616
rect 25504 22578 25556 22584
rect 24216 22568 24268 22574
rect 24216 22510 24268 22516
rect 24228 22234 24256 22510
rect 24216 22228 24268 22234
rect 24216 22170 24268 22176
rect 25516 22094 25544 22578
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 25424 22066 25544 22094
rect 24124 21140 24176 21146
rect 24124 21082 24176 21088
rect 24136 20942 24164 21082
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24136 17882 24164 20878
rect 25136 20868 25188 20874
rect 25136 20810 25188 20816
rect 25148 20602 25176 20810
rect 25424 20602 25452 22066
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34336 20868 34388 20874
rect 34336 20810 34388 20816
rect 25136 20596 25188 20602
rect 25136 20538 25188 20544
rect 25412 20596 25464 20602
rect 25412 20538 25464 20544
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24136 17678 24164 17818
rect 24124 17672 24176 17678
rect 24124 17614 24176 17620
rect 23296 17604 23348 17610
rect 23296 17546 23348 17552
rect 23112 17536 23164 17542
rect 23112 17478 23164 17484
rect 23124 16250 23152 17478
rect 23308 17338 23336 17546
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 23308 16250 23336 17274
rect 23112 16244 23164 16250
rect 23112 16186 23164 16192
rect 23296 16244 23348 16250
rect 23296 16186 23348 16192
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22848 14618 22876 16050
rect 24136 16046 24164 17614
rect 25136 17604 25188 17610
rect 25136 17546 25188 17552
rect 25148 17338 25176 17546
rect 25424 17338 25452 20538
rect 34348 20505 34376 20810
rect 34334 20496 34390 20505
rect 34334 20431 34390 20440
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33152 17542 33180 18702
rect 34888 18692 34940 18698
rect 34888 18634 34940 18640
rect 34900 18329 34928 18634
rect 34886 18320 34942 18329
rect 34886 18255 34942 18264
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 33140 17536 33192 17542
rect 33140 17478 33192 17484
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 25412 17332 25464 17338
rect 25412 17274 25464 17280
rect 25424 16114 25452 17274
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 33140 16584 33192 16590
rect 33140 16526 33192 16532
rect 33152 16250 33180 16526
rect 34888 16516 34940 16522
rect 34888 16458 34940 16464
rect 33140 16244 33192 16250
rect 33140 16186 33192 16192
rect 34900 16153 34928 16458
rect 34886 16144 34942 16153
rect 25412 16108 25464 16114
rect 25412 16050 25464 16056
rect 26056 16108 26108 16114
rect 34886 16079 34942 16088
rect 26056 16050 26108 16056
rect 24124 16040 24176 16046
rect 24124 15982 24176 15988
rect 24136 15706 24164 15982
rect 24124 15700 24176 15706
rect 24124 15642 24176 15648
rect 22836 14612 22888 14618
rect 22836 14554 22888 14560
rect 24136 14074 24164 15642
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 24136 13870 24164 14010
rect 26068 14006 26096 16050
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 33140 14408 33192 14414
rect 33140 14350 33192 14356
rect 33152 14074 33180 14350
rect 34888 14340 34940 14346
rect 34888 14282 34940 14288
rect 33140 14068 33192 14074
rect 33140 14010 33192 14016
rect 26056 14000 26108 14006
rect 34900 13977 34928 14282
rect 26056 13942 26108 13948
rect 34886 13968 34942 13977
rect 34886 13903 34942 13912
rect 23480 13864 23532 13870
rect 23480 13806 23532 13812
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 25044 13864 25096 13870
rect 25044 13806 25096 13812
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22652 13524 22704 13530
rect 22652 13466 22704 13472
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18616 12782 18644 13126
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 22112 12782 22140 13126
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 18604 12776 18656 12782
rect 18604 12718 18656 12724
rect 22100 12776 22152 12782
rect 22100 12718 22152 12724
rect 17880 12442 17908 12718
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 17132 12232 17184 12238
rect 17132 12174 17184 12180
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16776 11898 16804 12106
rect 16764 11892 16816 11898
rect 16764 11834 16816 11840
rect 16868 11830 16896 12106
rect 17512 12102 17540 12174
rect 17500 12096 17552 12102
rect 17500 12038 17552 12044
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 16856 11824 16908 11830
rect 16856 11766 16908 11772
rect 17512 11762 17540 12038
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 20732 11558 20760 12038
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 20720 11552 20772 11558
rect 20720 11494 20772 11500
rect 12636 11354 12664 11494
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 20732 11082 20760 11494
rect 12348 11076 12400 11082
rect 12348 11018 12400 11024
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10742 12664 10950
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 14464 10736 14516 10742
rect 14464 10678 14516 10684
rect 14476 10266 14504 10678
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10266 15240 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 10048 8900 10100 8906
rect 10048 8842 10100 8848
rect 9956 8832 10008 8838
rect 9956 8774 10008 8780
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 9968 3398 9996 8774
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 20732 3738 20760 11018
rect 21364 10464 21416 10470
rect 21364 10406 21416 10412
rect 21376 5710 21404 10406
rect 21652 5778 21680 12310
rect 22204 12306 22232 13262
rect 22468 13252 22520 13258
rect 22468 13194 22520 13200
rect 22480 12850 22508 13194
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22480 12442 22508 12786
rect 22468 12436 22520 12442
rect 22468 12378 22520 12384
rect 23492 12322 23520 13806
rect 23572 12640 23624 12646
rect 23572 12582 23624 12588
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 23308 12294 23520 12322
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 22008 12096 22060 12102
rect 22008 12038 22060 12044
rect 21836 11626 21864 12038
rect 22020 11694 22048 12038
rect 23308 11694 23336 12294
rect 23584 11830 23612 12582
rect 24400 12096 24452 12102
rect 24400 12038 24452 12044
rect 24952 12096 25004 12102
rect 25056 12084 25084 13806
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 33140 12232 33192 12238
rect 33140 12174 33192 12180
rect 25004 12056 25084 12084
rect 24952 12038 25004 12044
rect 24412 11830 24440 12038
rect 23572 11824 23624 11830
rect 23572 11766 23624 11772
rect 24400 11824 24452 11830
rect 24400 11766 24452 11772
rect 22008 11688 22060 11694
rect 22008 11630 22060 11636
rect 23296 11688 23348 11694
rect 23296 11630 23348 11636
rect 21824 11620 21876 11626
rect 21824 11562 21876 11568
rect 23308 11558 23336 11630
rect 23296 11552 23348 11558
rect 23296 11494 23348 11500
rect 23480 11552 23532 11558
rect 23480 11494 23532 11500
rect 23308 10606 23336 11494
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23296 10600 23348 10606
rect 23296 10542 23348 10548
rect 23400 10062 23428 10950
rect 23492 10742 23520 11494
rect 24964 11150 24992 12038
rect 33152 11898 33180 12174
rect 34888 12164 34940 12170
rect 34888 12106 34940 12112
rect 33140 11892 33192 11898
rect 33140 11834 33192 11840
rect 34900 11801 34928 12106
rect 34886 11792 34942 11801
rect 34886 11727 34942 11736
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 23480 10736 23532 10742
rect 23480 10678 23532 10684
rect 24872 10674 24900 11018
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 33140 10464 33192 10470
rect 33140 10406 33192 10412
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 23388 10056 23440 10062
rect 23388 9998 23440 10004
rect 23400 6914 23428 9998
rect 32968 8090 32996 10202
rect 33152 10062 33180 10406
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 33140 10056 33192 10062
rect 33140 9998 33192 10004
rect 34336 9988 34388 9994
rect 34336 9930 34388 9936
rect 34348 9625 34376 9930
rect 34334 9616 34390 9625
rect 34334 9551 34390 9560
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 34888 7812 34940 7818
rect 34888 7754 34940 7760
rect 34900 7449 34928 7754
rect 34886 7440 34942 7449
rect 34886 7375 34942 7384
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 23216 6886 23428 6914
rect 21640 5772 21692 5778
rect 21640 5714 21692 5720
rect 23216 5710 23244 6886
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 23204 5704 23256 5710
rect 23204 5646 23256 5652
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20720 3732 20772 3738
rect 20720 3674 20772 3680
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 9968 2514 9996 3334
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 20732 3194 20760 3674
rect 20824 3534 20852 5510
rect 23216 3534 23244 5646
rect 34336 5636 34388 5642
rect 34336 5578 34388 5584
rect 34348 5273 34376 5578
rect 34334 5264 34390 5273
rect 34334 5199 34390 5208
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23216 3398 23244 3470
rect 34888 3460 34940 3466
rect 34888 3402 34940 3408
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 20720 3188 20772 3194
rect 20720 3130 20772 3136
rect 23216 2514 23244 3334
rect 34900 3097 34928 3402
rect 34886 3088 34942 3097
rect 34886 3023 34942 3032
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 23204 2508 23256 2514
rect 23204 2450 23256 2456
rect 940 2440 992 2446
rect 940 2382 992 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 27344 2440 27396 2446
rect 27344 2382 27396 2388
rect 952 2009 980 2382
rect 938 2000 994 2009
rect 938 1935 994 1944
rect 9140 1306 9168 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 27356 1306 27384 2382
rect 9048 1278 9168 1306
rect 27264 1278 27384 1306
rect 9048 800 9076 1278
rect 27264 800 27292 1278
rect 9034 0 9090 800
rect 27250 0 27306 800
<< via2 >>
rect 938 36760 994 36816
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 938 34584 994 34640
rect 938 32408 994 32464
rect 1398 30232 1454 30288
rect 938 28056 994 28112
rect 1398 26152 1454 26208
rect 938 23704 994 23760
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 34334 35672 34390 35728
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34886 33496 34942 33552
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 938 21528 994 21584
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 938 19352 994 19408
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 938 17176 994 17232
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 1398 15136 1454 15192
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 938 12824 994 12880
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 1398 10920 1454 10976
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 938 8472 994 8528
rect 9310 19896 9366 19952
rect 9494 20748 9496 20768
rect 9496 20748 9548 20768
rect 9548 20748 9550 20768
rect 9494 20712 9550 20748
rect 9862 21412 9918 21448
rect 9862 21392 9864 21412
rect 9864 21392 9916 21412
rect 9916 21392 9918 21412
rect 8574 17040 8630 17096
rect 9586 17040 9642 17096
rect 10230 20576 10286 20632
rect 11610 21428 11612 21448
rect 11612 21428 11664 21448
rect 11664 21428 11666 21448
rect 11610 21392 11666 21428
rect 10230 16652 10286 16688
rect 10230 16632 10232 16652
rect 10232 16632 10284 16652
rect 10284 16632 10286 16652
rect 10690 14864 10746 14920
rect 11702 19372 11758 19408
rect 11702 19352 11704 19372
rect 11704 19352 11756 19372
rect 11756 19352 11758 19372
rect 11702 14456 11758 14512
rect 10966 14184 11022 14240
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 938 6296 994 6352
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 938 4120 994 4176
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11518 13912 11574 13968
rect 12714 24404 12770 24440
rect 12714 24384 12716 24404
rect 12716 24384 12768 24404
rect 12768 24384 12770 24404
rect 12070 19352 12126 19408
rect 15106 24404 15162 24440
rect 15106 24384 15108 24404
rect 15108 24384 15160 24404
rect 15160 24384 15162 24404
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 34334 31320 34390 31376
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 12162 16108 12218 16144
rect 12162 16088 12164 16108
rect 12164 16088 12216 16108
rect 12216 16088 12218 16108
rect 12990 16224 13046 16280
rect 12990 16108 13046 16144
rect 12990 16088 12992 16108
rect 12992 16088 13044 16108
rect 13044 16088 13046 16108
rect 14002 20748 14004 20768
rect 14004 20748 14056 20768
rect 14056 20748 14058 20768
rect 14002 20712 14058 20748
rect 14738 19896 14794 19952
rect 13634 16224 13690 16280
rect 12714 14864 12770 14920
rect 12162 14356 12164 14376
rect 12164 14356 12216 14376
rect 12216 14356 12218 14376
rect 12162 14320 12218 14356
rect 12990 14320 13046 14376
rect 11518 12180 11520 12200
rect 11520 12180 11572 12200
rect 11572 12180 11574 12200
rect 11518 12144 11574 12180
rect 14830 16632 14886 16688
rect 13634 14356 13636 14376
rect 13636 14356 13688 14376
rect 13688 14356 13690 14376
rect 13634 14320 13690 14356
rect 13818 14184 13874 14240
rect 13450 13932 13506 13968
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 34886 29144 34942 29200
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34886 26968 34942 27024
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 14646 14456 14702 14512
rect 13450 13912 13452 13932
rect 13452 13912 13504 13932
rect 13504 13912 13506 13932
rect 14370 13932 14426 13968
rect 14370 13912 14372 13932
rect 14372 13912 14424 13932
rect 14424 13912 14426 13932
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 16302 12144 16358 12200
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34334 24792 34390 24848
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34886 22616 34942 22672
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34334 20440 34390 20496
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34886 18264 34942 18320
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34886 16088 34942 16144
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34886 13912 34942 13968
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34886 11736 34942 11792
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34334 9560 34390 9616
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34886 7384 34942 7440
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34334 5208 34390 5264
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34886 3032 34942 3088
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 938 1944 994 2000
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 34329 35730 34395 35733
rect 35600 35730 36400 35760
rect 34329 35728 36400 35730
rect 34329 35672 34334 35728
rect 34390 35672 36400 35728
rect 34329 35670 36400 35672
rect 34329 35667 34395 35670
rect 35600 35640 36400 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 0 34642 800 34672
rect 933 34642 999 34645
rect 0 34640 999 34642
rect 0 34584 938 34640
rect 994 34584 999 34640
rect 0 34582 999 34584
rect 0 34552 800 34582
rect 933 34579 999 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 34881 33554 34947 33557
rect 35600 33554 36400 33584
rect 34881 33552 36400 33554
rect 34881 33496 34886 33552
rect 34942 33496 36400 33552
rect 34881 33494 36400 33496
rect 34881 33491 34947 33494
rect 35600 33464 36400 33494
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 0 32466 800 32496
rect 933 32466 999 32469
rect 0 32464 999 32466
rect 0 32408 938 32464
rect 994 32408 999 32464
rect 0 32406 999 32408
rect 0 32376 800 32406
rect 933 32403 999 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 34329 31378 34395 31381
rect 35600 31378 36400 31408
rect 34329 31376 36400 31378
rect 34329 31320 34334 31376
rect 34390 31320 36400 31376
rect 34329 31318 36400 31320
rect 34329 31315 34395 31318
rect 35600 31288 36400 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 30290 800 30320
rect 1393 30290 1459 30293
rect 0 30288 1459 30290
rect 0 30232 1398 30288
rect 1454 30232 1459 30288
rect 0 30230 1459 30232
rect 0 30200 800 30230
rect 1393 30227 1459 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 34881 29202 34947 29205
rect 35600 29202 36400 29232
rect 34881 29200 36400 29202
rect 34881 29144 34886 29200
rect 34942 29144 36400 29200
rect 34881 29142 36400 29144
rect 34881 29139 34947 29142
rect 35600 29112 36400 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 0 28114 800 28144
rect 933 28114 999 28117
rect 0 28112 999 28114
rect 0 28056 938 28112
rect 994 28056 999 28112
rect 0 28054 999 28056
rect 0 28024 800 28054
rect 933 28051 999 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 34881 27026 34947 27029
rect 35600 27026 36400 27056
rect 34881 27024 36400 27026
rect 34881 26968 34886 27024
rect 34942 26968 36400 27024
rect 34881 26966 36400 26968
rect 34881 26963 34947 26966
rect 35600 26936 36400 26966
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1393 26210 1459 26213
rect 798 26208 1459 26210
rect 798 26152 1398 26208
rect 1454 26152 1459 26208
rect 798 26150 1459 26152
rect 798 25968 858 26150
rect 1393 26147 1459 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25878 858 25968
rect 0 25848 800 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 34329 24850 34395 24853
rect 35600 24850 36400 24880
rect 34329 24848 36400 24850
rect 34329 24792 34334 24848
rect 34390 24792 36400 24848
rect 34329 24790 36400 24792
rect 34329 24787 34395 24790
rect 35600 24760 36400 24790
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 12709 24442 12775 24445
rect 15101 24442 15167 24445
rect 12709 24440 15167 24442
rect 12709 24384 12714 24440
rect 12770 24384 15106 24440
rect 15162 24384 15167 24440
rect 12709 24382 15167 24384
rect 12709 24379 12775 24382
rect 15101 24379 15167 24382
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 0 23762 800 23792
rect 933 23762 999 23765
rect 0 23760 999 23762
rect 0 23704 938 23760
rect 994 23704 999 23760
rect 0 23702 999 23704
rect 0 23672 800 23702
rect 933 23699 999 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 34881 22674 34947 22677
rect 35600 22674 36400 22704
rect 34881 22672 36400 22674
rect 34881 22616 34886 22672
rect 34942 22616 36400 22672
rect 34881 22614 36400 22616
rect 34881 22611 34947 22614
rect 35600 22584 36400 22614
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 0 21586 800 21616
rect 933 21586 999 21589
rect 0 21584 999 21586
rect 0 21528 938 21584
rect 994 21528 999 21584
rect 0 21526 999 21528
rect 0 21496 800 21526
rect 933 21523 999 21526
rect 9857 21450 9923 21453
rect 11605 21450 11671 21453
rect 9857 21448 11671 21450
rect 9857 21392 9862 21448
rect 9918 21392 11610 21448
rect 11666 21392 11671 21448
rect 9857 21390 11671 21392
rect 9857 21387 9923 21390
rect 11605 21387 11671 21390
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 9489 20770 9555 20773
rect 13997 20770 14063 20773
rect 9489 20768 14063 20770
rect 9489 20712 9494 20768
rect 9550 20712 14002 20768
rect 14058 20712 14063 20768
rect 9489 20710 14063 20712
rect 9489 20707 9555 20710
rect 10182 20637 10242 20710
rect 13997 20707 14063 20710
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 10182 20632 10291 20637
rect 10182 20576 10230 20632
rect 10286 20576 10291 20632
rect 10182 20574 10291 20576
rect 10225 20571 10291 20574
rect 34329 20498 34395 20501
rect 35600 20498 36400 20528
rect 34329 20496 36400 20498
rect 34329 20440 34334 20496
rect 34390 20440 36400 20496
rect 34329 20438 36400 20440
rect 34329 20435 34395 20438
rect 35600 20408 36400 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 9305 19954 9371 19957
rect 14733 19954 14799 19957
rect 9305 19952 14799 19954
rect 9305 19896 9310 19952
rect 9366 19896 14738 19952
rect 14794 19896 14799 19952
rect 9305 19894 14799 19896
rect 9305 19891 9371 19894
rect 14733 19891 14799 19894
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 11697 19410 11763 19413
rect 12065 19410 12131 19413
rect 11697 19408 12131 19410
rect 11697 19352 11702 19408
rect 11758 19352 12070 19408
rect 12126 19352 12131 19408
rect 11697 19350 12131 19352
rect 11697 19347 11763 19350
rect 12065 19347 12131 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 34881 18322 34947 18325
rect 35600 18322 36400 18352
rect 34881 18320 36400 18322
rect 34881 18264 34886 18320
rect 34942 18264 36400 18320
rect 34881 18262 36400 18264
rect 34881 18259 34947 18262
rect 35600 18232 36400 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 0 17234 800 17264
rect 933 17234 999 17237
rect 0 17232 999 17234
rect 0 17176 938 17232
rect 994 17176 999 17232
rect 0 17174 999 17176
rect 0 17144 800 17174
rect 933 17171 999 17174
rect 8569 17098 8635 17101
rect 9581 17098 9647 17101
rect 8569 17096 9647 17098
rect 8569 17040 8574 17096
rect 8630 17040 9586 17096
rect 9642 17040 9647 17096
rect 8569 17038 9647 17040
rect 8569 17035 8635 17038
rect 9581 17035 9647 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 10225 16690 10291 16693
rect 14825 16690 14891 16693
rect 10225 16688 14891 16690
rect 10225 16632 10230 16688
rect 10286 16632 14830 16688
rect 14886 16632 14891 16688
rect 10225 16630 14891 16632
rect 10225 16627 10291 16630
rect 14825 16627 14891 16630
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 12985 16282 13051 16285
rect 13629 16282 13695 16285
rect 12985 16280 13695 16282
rect 12985 16224 12990 16280
rect 13046 16224 13634 16280
rect 13690 16224 13695 16280
rect 12985 16222 13695 16224
rect 12985 16219 13051 16222
rect 13629 16219 13695 16222
rect 12157 16146 12223 16149
rect 12985 16146 13051 16149
rect 12157 16144 13051 16146
rect 12157 16088 12162 16144
rect 12218 16088 12990 16144
rect 13046 16088 13051 16144
rect 12157 16086 13051 16088
rect 12157 16083 12223 16086
rect 12985 16083 13051 16086
rect 34881 16146 34947 16149
rect 35600 16146 36400 16176
rect 34881 16144 36400 16146
rect 34881 16088 34886 16144
rect 34942 16088 36400 16144
rect 34881 16086 36400 16088
rect 34881 16083 34947 16086
rect 35600 16056 36400 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 1393 15194 1459 15197
rect 798 15192 1459 15194
rect 798 15136 1398 15192
rect 1454 15136 1459 15192
rect 798 15134 1459 15136
rect 798 15088 858 15134
rect 1393 15131 1459 15134
rect 0 14998 858 15088
rect 0 14968 800 14998
rect 10685 14922 10751 14925
rect 12709 14922 12775 14925
rect 10685 14920 12775 14922
rect 10685 14864 10690 14920
rect 10746 14864 12714 14920
rect 12770 14864 12775 14920
rect 10685 14862 12775 14864
rect 10685 14859 10751 14862
rect 12709 14859 12775 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 11697 14514 11763 14517
rect 14641 14514 14707 14517
rect 11697 14512 14707 14514
rect 11697 14456 11702 14512
rect 11758 14456 14646 14512
rect 14702 14456 14707 14512
rect 11697 14454 14707 14456
rect 11697 14451 11763 14454
rect 14641 14451 14707 14454
rect 12157 14378 12223 14381
rect 12985 14378 13051 14381
rect 13629 14378 13695 14381
rect 12157 14376 13695 14378
rect 12157 14320 12162 14376
rect 12218 14320 12990 14376
rect 13046 14320 13634 14376
rect 13690 14320 13695 14376
rect 12157 14318 13695 14320
rect 12157 14315 12223 14318
rect 12985 14315 13051 14318
rect 13629 14315 13695 14318
rect 10961 14242 11027 14245
rect 13813 14242 13879 14245
rect 10961 14240 13879 14242
rect 10961 14184 10966 14240
rect 11022 14184 13818 14240
rect 13874 14184 13879 14240
rect 10961 14182 13879 14184
rect 10961 14179 11027 14182
rect 13813 14179 13879 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 11513 13970 11579 13973
rect 13445 13970 13511 13973
rect 14365 13970 14431 13973
rect 11513 13968 14431 13970
rect 11513 13912 11518 13968
rect 11574 13912 13450 13968
rect 13506 13912 14370 13968
rect 14426 13912 14431 13968
rect 11513 13910 14431 13912
rect 11513 13907 11579 13910
rect 13445 13907 13511 13910
rect 14365 13907 14431 13910
rect 34881 13970 34947 13973
rect 35600 13970 36400 14000
rect 34881 13968 36400 13970
rect 34881 13912 34886 13968
rect 34942 13912 36400 13968
rect 34881 13910 36400 13912
rect 34881 13907 34947 13910
rect 35600 13880 36400 13910
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 11513 12202 11579 12205
rect 16297 12202 16363 12205
rect 11513 12200 16363 12202
rect 11513 12144 11518 12200
rect 11574 12144 16302 12200
rect 16358 12144 16363 12200
rect 11513 12142 16363 12144
rect 11513 12139 11579 12142
rect 16297 12139 16363 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 34881 11794 34947 11797
rect 35600 11794 36400 11824
rect 34881 11792 36400 11794
rect 34881 11736 34886 11792
rect 34942 11736 36400 11792
rect 34881 11734 36400 11736
rect 34881 11731 34947 11734
rect 35600 11704 36400 11734
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 1393 10978 1459 10981
rect 798 10976 1459 10978
rect 798 10920 1398 10976
rect 1454 10920 1459 10976
rect 798 10918 1459 10920
rect 798 10736 858 10918
rect 1393 10915 1459 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 0 10646 858 10736
rect 0 10616 800 10646
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 34329 9618 34395 9621
rect 35600 9618 36400 9648
rect 34329 9616 36400 9618
rect 34329 9560 34334 9616
rect 34390 9560 36400 9616
rect 34329 9558 36400 9560
rect 34329 9555 34395 9558
rect 35600 9528 36400 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 0 8530 800 8560
rect 933 8530 999 8533
rect 0 8528 999 8530
rect 0 8472 938 8528
rect 994 8472 999 8528
rect 0 8470 999 8472
rect 0 8440 800 8470
rect 933 8467 999 8470
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 34881 7442 34947 7445
rect 35600 7442 36400 7472
rect 34881 7440 36400 7442
rect 34881 7384 34886 7440
rect 34942 7384 36400 7440
rect 34881 7382 36400 7384
rect 34881 7379 34947 7382
rect 35600 7352 36400 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 34329 5266 34395 5269
rect 35600 5266 36400 5296
rect 34329 5264 36400 5266
rect 34329 5208 34334 5264
rect 34390 5208 36400 5264
rect 34329 5206 36400 5208
rect 34329 5203 34395 5206
rect 35600 5176 36400 5206
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 34881 3090 34947 3093
rect 35600 3090 36400 3120
rect 34881 3088 36400 3090
rect 34881 3032 34886 3088
rect 34942 3032 36400 3088
rect 34881 3030 36400 3032
rect 34881 3027 34947 3030
rect 35600 3000 36400 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 0 2002 800 2032
rect 933 2002 999 2005
rect 0 2000 999 2002
rect 0 1944 938 2000
rect 994 1944 999 2000
rect 0 1942 999 1944
rect 0 1912 800 1942
rect 933 1939 999 1942
<< via3 >>
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 36480 4528 36496
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 35936 19888 36496
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 36480 35248 36496
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__inv_2  _413_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _414_
timestamp 1688980957
transform 1 0 9936 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _415_
timestamp 1688980957
transform -1 0 22908 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _416_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10672 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _417_
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _418_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _419_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _420_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7176 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _421_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_4  _422_
timestamp 1688980957
transform 1 0 6440 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_2  _423_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _424_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _425_
timestamp 1688980957
transform 1 0 7544 0 -1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__o22a_1  _426_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12604 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _427_
timestamp 1688980957
transform 1 0 9476 0 1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _428_
timestamp 1688980957
transform 1 0 9384 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _429_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _430_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _431_
timestamp 1688980957
transform 1 0 7360 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _432_
timestamp 1688980957
transform 1 0 7360 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _433_
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_4  _434_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5060 0 1 19584
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_4  _435_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _436_
timestamp 1688980957
transform 1 0 6348 0 1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _437_
timestamp 1688980957
transform -1 0 10856 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _438_
timestamp 1688980957
transform -1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _439_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11408 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _440_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11316 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _441_
timestamp 1688980957
transform 1 0 11408 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o311a_4  _443_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_4  _444_
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _445_
timestamp 1688980957
transform 1 0 6072 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_2  _446_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _447_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_4  _448_
timestamp 1688980957
transform 1 0 6164 0 1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_4  _449_
timestamp 1688980957
transform 1 0 6348 0 1 17408
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _450_
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_2  _451_
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _452_
timestamp 1688980957
transform 1 0 10488 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_2  _453_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _454_
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _455_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12328 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _456_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _457_
timestamp 1688980957
transform -1 0 15088 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _458_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16560 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _459_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _460_
timestamp 1688980957
transform 1 0 15640 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _461_
timestamp 1688980957
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_1  _462_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _463_
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _464_
timestamp 1688980957
transform 1 0 17296 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _465_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21804 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _466_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _467_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 6808 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _468_
timestamp 1688980957
transform 1 0 6808 0 1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1688980957
transform 1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _470_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_4  _471_
timestamp 1688980957
transform 1 0 7728 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _472_
timestamp 1688980957
transform -1 0 8372 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _473_
timestamp 1688980957
transform 1 0 7268 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _474_
timestamp 1688980957
transform 1 0 12880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _475_
timestamp 1688980957
transform 1 0 16100 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _476_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _477_
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _478_
timestamp 1688980957
transform -1 0 15640 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _479_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _480_
timestamp 1688980957
transform 1 0 12420 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _481_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _482_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _483_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _484_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _485_
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _486_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _487_
timestamp 1688980957
transform -1 0 19044 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _488_
timestamp 1688980957
transform 1 0 20332 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _489_
timestamp 1688980957
transform -1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _490_
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _491_
timestamp 1688980957
transform 1 0 21528 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _492_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22448 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _493_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _494_
timestamp 1688980957
transform 1 0 14628 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _495_
timestamp 1688980957
transform 1 0 16192 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _496_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13432 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _497_
timestamp 1688980957
transform 1 0 13616 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _498_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13616 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _499_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _500_
timestamp 1688980957
transform -1 0 17940 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_2  _501_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17480 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_1  _502_
timestamp 1688980957
transform 1 0 17296 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _503_
timestamp 1688980957
transform 1 0 18768 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _504_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _505_
timestamp 1688980957
transform -1 0 20332 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _506_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8004 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _507_
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _508_
timestamp 1688980957
transform 1 0 8372 0 -1 25024
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_1  _509_
timestamp 1688980957
transform 1 0 12972 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _510_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9568 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _511_
timestamp 1688980957
transform 1 0 13524 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _512_
timestamp 1688980957
transform -1 0 10120 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _513_
timestamp 1688980957
transform 1 0 7728 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _514_
timestamp 1688980957
transform 1 0 7636 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__or4_1  _515_
timestamp 1688980957
transform 1 0 12328 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _516_
timestamp 1688980957
transform -1 0 9292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _517_
timestamp 1688980957
transform 1 0 13340 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _518_
timestamp 1688980957
transform 1 0 15272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _519_
timestamp 1688980957
transform -1 0 15824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _520_
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _521_
timestamp 1688980957
transform -1 0 16928 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _522_
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _523_
timestamp 1688980957
transform 1 0 17112 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _524_
timestamp 1688980957
transform -1 0 20700 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _525_
timestamp 1688980957
transform -1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _526_
timestamp 1688980957
transform 1 0 21068 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _527_
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _528_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a2111o_1  _529_
timestamp 1688980957
transform -1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _530_
timestamp 1688980957
transform 1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _531_
timestamp 1688980957
transform 1 0 16008 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_1  _532_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15732 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2a_1  _533_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _534_
timestamp 1688980957
transform -1 0 19780 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _535_
timestamp 1688980957
transform 1 0 18676 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _536_
timestamp 1688980957
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_2  _537_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _538_
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _539_
timestamp 1688980957
transform -1 0 12052 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _540_
timestamp 1688980957
transform 1 0 12512 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _541_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _542_
timestamp 1688980957
transform -1 0 13248 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _543_
timestamp 1688980957
transform -1 0 12972 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _544_
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _545_
timestamp 1688980957
transform 1 0 13616 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _546_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10856 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_2  _547_
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _548_
timestamp 1688980957
transform 1 0 5888 0 1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_2  _549_
timestamp 1688980957
transform 1 0 10856 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _550_
timestamp 1688980957
transform -1 0 13340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _551_
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _552_
timestamp 1688980957
transform -1 0 12604 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _553_
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _554_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _555_
timestamp 1688980957
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _556_
timestamp 1688980957
transform 1 0 16192 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _557_
timestamp 1688980957
transform 1 0 16744 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _558_
timestamp 1688980957
transform 1 0 19872 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _559_
timestamp 1688980957
transform 1 0 20792 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _560_
timestamp 1688980957
transform 1 0 21252 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _561_
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _562_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23184 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _563_
timestamp 1688980957
transform 1 0 20148 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _564_
timestamp 1688980957
transform 1 0 19320 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _565_
timestamp 1688980957
transform 1 0 15640 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _566_
timestamp 1688980957
transform -1 0 8188 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_4  _567_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6624 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  _568_
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_2  _569_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 11592 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _570_
timestamp 1688980957
transform -1 0 10856 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _571_
timestamp 1688980957
transform 1 0 10120 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _572_
timestamp 1688980957
transform -1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nand4_1  _573_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _574_
timestamp 1688980957
transform 1 0 10672 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _575_
timestamp 1688980957
transform -1 0 13984 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _576_
timestamp 1688980957
transform -1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _577_
timestamp 1688980957
transform -1 0 13800 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _578_
timestamp 1688980957
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_2  _579_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13524 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _580_
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_4  _581_
timestamp 1688980957
transform -1 0 8832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_1  _582_
timestamp 1688980957
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _583_
timestamp 1688980957
transform -1 0 5888 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_4  _584_
timestamp 1688980957
transform 1 0 6256 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__or4b_4  _585_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10304 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__a2bb2o_1  _586_
timestamp 1688980957
transform -1 0 8556 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _587_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _588_
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _589_
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _590_
timestamp 1688980957
transform 1 0 11868 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _591_
timestamp 1688980957
transform -1 0 11868 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _592_
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _593_
timestamp 1688980957
transform 1 0 12236 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _594_
timestamp 1688980957
transform -1 0 12604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _595_
timestamp 1688980957
transform 1 0 13156 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _596_
timestamp 1688980957
transform -1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _597_
timestamp 1688980957
transform -1 0 19136 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _598_
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _599_
timestamp 1688980957
transform 1 0 18400 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _600_
timestamp 1688980957
transform -1 0 19136 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _601_
timestamp 1688980957
transform 1 0 21344 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _602_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _603_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21344 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _604_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _605_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _606_
timestamp 1688980957
transform 1 0 23184 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _607_
timestamp 1688980957
transform 1 0 12696 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _608_
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _609_
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _610_
timestamp 1688980957
transform -1 0 16008 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _611_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9844 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _612_
timestamp 1688980957
transform -1 0 10948 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _613_
timestamp 1688980957
transform -1 0 10304 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _614_
timestamp 1688980957
transform 1 0 9384 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _615_
timestamp 1688980957
transform -1 0 13432 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _616_
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _617_
timestamp 1688980957
transform 1 0 14168 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _618_
timestamp 1688980957
transform 1 0 16008 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _619_
timestamp 1688980957
transform 1 0 15364 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _620_
timestamp 1688980957
transform -1 0 15272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _621_
timestamp 1688980957
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _622_
timestamp 1688980957
transform -1 0 10212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _623_
timestamp 1688980957
transform -1 0 10580 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a32oi_4  _624_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10212 0 1 15232
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _625_
timestamp 1688980957
transform 1 0 10948 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _626_
timestamp 1688980957
transform 1 0 10580 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _627_
timestamp 1688980957
transform 1 0 10212 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _628_
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _629_
timestamp 1688980957
transform 1 0 17480 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _630_
timestamp 1688980957
transform 1 0 16836 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _631_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _632_
timestamp 1688980957
transform 1 0 18400 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _633_
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _634_
timestamp 1688980957
transform 1 0 19504 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _635_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _636_
timestamp 1688980957
transform 1 0 20424 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _637_
timestamp 1688980957
transform -1 0 21160 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _638_
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _639_
timestamp 1688980957
transform 1 0 22264 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _640_
timestamp 1688980957
transform 1 0 22724 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and4bb_1  _641_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__o22a_1  _642_
timestamp 1688980957
transform -1 0 12696 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _643_
timestamp 1688980957
transform 1 0 13156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _644_
timestamp 1688980957
transform -1 0 20056 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _645_
timestamp 1688980957
transform 1 0 14352 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _646_
timestamp 1688980957
transform -1 0 15640 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _647_
timestamp 1688980957
transform 1 0 15364 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _648_
timestamp 1688980957
transform -1 0 11408 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _649_
timestamp 1688980957
transform -1 0 11040 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _650_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _651_
timestamp 1688980957
transform 1 0 10304 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand3b_1  _652_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _653_
timestamp 1688980957
transform -1 0 14168 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _654_
timestamp 1688980957
transform 1 0 16100 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _655_
timestamp 1688980957
transform -1 0 16468 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _656_
timestamp 1688980957
transform 1 0 17480 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _657_
timestamp 1688980957
transform -1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2oi_1  _658_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15180 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _659_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15088 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _660_
timestamp 1688980957
transform 1 0 8740 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _661_
timestamp 1688980957
transform -1 0 9936 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  _662_
timestamp 1688980957
transform -1 0 10580 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _663_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13248 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _664_
timestamp 1688980957
transform -1 0 14536 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _665_
timestamp 1688980957
transform 1 0 15548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _666_
timestamp 1688980957
transform -1 0 15548 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _667_
timestamp 1688980957
transform 1 0 17572 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _668_
timestamp 1688980957
transform -1 0 18308 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _669_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_1  _670_
timestamp 1688980957
transform -1 0 18400 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _671_
timestamp 1688980957
transform -1 0 19780 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _672_
timestamp 1688980957
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _673_
timestamp 1688980957
transform -1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _674_
timestamp 1688980957
transform -1 0 20700 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _675_
timestamp 1688980957
transform 1 0 20424 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _676_
timestamp 1688980957
transform -1 0 20424 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _677_
timestamp 1688980957
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _678_
timestamp 1688980957
transform 1 0 21620 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _679_
timestamp 1688980957
transform -1 0 23460 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _680_
timestamp 1688980957
transform -1 0 21528 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _681_
timestamp 1688980957
transform -1 0 11592 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _682_
timestamp 1688980957
transform -1 0 15456 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _683_
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _684_
timestamp 1688980957
transform -1 0 17480 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _685_
timestamp 1688980957
transform 1 0 16560 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _686_
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _687_
timestamp 1688980957
transform -1 0 15272 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _688_
timestamp 1688980957
transform 1 0 15272 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _689_
timestamp 1688980957
transform -1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _690_
timestamp 1688980957
transform 1 0 16560 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _691_
timestamp 1688980957
transform 1 0 16652 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _692_
timestamp 1688980957
transform 1 0 18216 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _693_
timestamp 1688980957
transform 1 0 17572 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _694_
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _695_
timestamp 1688980957
transform 1 0 18492 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _696_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19780 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _697_
timestamp 1688980957
transform 1 0 19596 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _698_
timestamp 1688980957
transform -1 0 12512 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _699_
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _700_
timestamp 1688980957
transform -1 0 12880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _701_
timestamp 1688980957
transform -1 0 13432 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _702_
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _703_
timestamp 1688980957
transform -1 0 13708 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _704_
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _705_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _706_
timestamp 1688980957
transform 1 0 20424 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _707_
timestamp 1688980957
transform 1 0 20608 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _708_
timestamp 1688980957
transform 1 0 21160 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _709_
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _710_
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _711_
timestamp 1688980957
transform 1 0 20884 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o41a_1  _712_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15732 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21boi_1  _713_
timestamp 1688980957
transform 1 0 16008 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _714_
timestamp 1688980957
transform -1 0 16008 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _715_
timestamp 1688980957
transform 1 0 16744 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _716_
timestamp 1688980957
transform -1 0 17664 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _717_
timestamp 1688980957
transform 1 0 16744 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _718_
timestamp 1688980957
transform 1 0 18216 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _719_
timestamp 1688980957
transform -1 0 19136 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _720_
timestamp 1688980957
transform 1 0 17940 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _721_
timestamp 1688980957
transform 1 0 19688 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _722_
timestamp 1688980957
transform 1 0 19044 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _723_
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o22ai_1  _724_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12144 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _725_
timestamp 1688980957
transform -1 0 12236 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _726_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10304 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _727_
timestamp 1688980957
transform 1 0 11040 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _728_
timestamp 1688980957
transform 1 0 10580 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _729_
timestamp 1688980957
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _730_
timestamp 1688980957
transform 1 0 11684 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _731_
timestamp 1688980957
transform 1 0 11592 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _732_
timestamp 1688980957
transform 1 0 12144 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _733_
timestamp 1688980957
transform 1 0 12788 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _734_
timestamp 1688980957
transform 1 0 13616 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _735_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13984 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _736_
timestamp 1688980957
transform 1 0 14444 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _737_
timestamp 1688980957
transform -1 0 21436 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _738_
timestamp 1688980957
transform 1 0 19688 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _739_
timestamp 1688980957
transform 1 0 20332 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _740_
timestamp 1688980957
transform 1 0 21344 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _741_
timestamp 1688980957
transform 1 0 23460 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _742_
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _743_
timestamp 1688980957
transform -1 0 12604 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _744_
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _745_
timestamp 1688980957
transform -1 0 13064 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _746_
timestamp 1688980957
transform 1 0 12144 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _747_
timestamp 1688980957
transform -1 0 13248 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _748_
timestamp 1688980957
transform 1 0 11868 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _749_
timestamp 1688980957
transform -1 0 12604 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _750_
timestamp 1688980957
transform 1 0 12328 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _751_
timestamp 1688980957
transform -1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _752_
timestamp 1688980957
transform -1 0 15364 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _753_
timestamp 1688980957
transform -1 0 14904 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _754_
timestamp 1688980957
transform 1 0 17112 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _755_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor4_1  _756_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18308 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _757_
timestamp 1688980957
transform 1 0 20056 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _758_
timestamp 1688980957
transform -1 0 21344 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _759_
timestamp 1688980957
transform 1 0 20700 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _760_
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _761_
timestamp 1688980957
transform -1 0 16008 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2b_1  _762_
timestamp 1688980957
transform 1 0 15456 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _763_
timestamp 1688980957
transform -1 0 16284 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _764_
timestamp 1688980957
transform -1 0 14352 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _765_
timestamp 1688980957
transform 1 0 13616 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _766_
timestamp 1688980957
transform 1 0 14168 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _767_
timestamp 1688980957
transform -1 0 13432 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _768_
timestamp 1688980957
transform -1 0 14904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _769_
timestamp 1688980957
transform 1 0 13984 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _770_
timestamp 1688980957
transform 1 0 15364 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _771_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _772_
timestamp 1688980957
transform -1 0 16284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _773_
timestamp 1688980957
transform 1 0 16928 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _774_
timestamp 1688980957
transform -1 0 18492 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _775_
timestamp 1688980957
transform -1 0 17572 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _776_
timestamp 1688980957
transform 1 0 17848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _777_
timestamp 1688980957
transform 1 0 20148 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _778_
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _779_
timestamp 1688980957
transform -1 0 19872 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _780_
timestamp 1688980957
transform 1 0 19872 0 -1 27200
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _781_
timestamp 1688980957
transform -1 0 15640 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _782_
timestamp 1688980957
transform -1 0 16008 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _783_
timestamp 1688980957
transform 1 0 15732 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _784_
timestamp 1688980957
transform -1 0 18032 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _785_
timestamp 1688980957
transform -1 0 17480 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _786_
timestamp 1688980957
transform 1 0 18308 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _787_
timestamp 1688980957
transform -1 0 15824 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _788_
timestamp 1688980957
transform -1 0 19228 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _789_
timestamp 1688980957
transform -1 0 22724 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _790_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _791_
timestamp 1688980957
transform -1 0 22080 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _792_
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _793_
timestamp 1688980957
transform 1 0 22816 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _794_
timestamp 1688980957
transform -1 0 23092 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _795_
timestamp 1688980957
transform 1 0 23276 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _796_
timestamp 1688980957
transform 1 0 22816 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _797_
timestamp 1688980957
transform 1 0 23276 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _798_
timestamp 1688980957
transform 1 0 22816 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _799_
timestamp 1688980957
transform 1 0 22632 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _800_
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _801_
timestamp 1688980957
transform 1 0 23184 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _802_
timestamp 1688980957
transform 1 0 22540 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _803_
timestamp 1688980957
transform 1 0 22080 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _804_
timestamp 1688980957
transform 1 0 21896 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _805_
timestamp 1688980957
transform -1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _806_
timestamp 1688980957
transform 1 0 12052 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _807_
timestamp 1688980957
transform -1 0 20976 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _808_
timestamp 1688980957
transform -1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _809_
timestamp 1688980957
transform 1 0 20056 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _810_
timestamp 1688980957
transform -1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _811_
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _812_
timestamp 1688980957
transform 1 0 24472 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _813_
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _814_
timestamp 1688980957
transform -1 0 25852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _815_
timestamp 1688980957
transform -1 0 25944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _816_
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _817_
timestamp 1688980957
transform 1 0 24932 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _818_
timestamp 1688980957
transform -1 0 26036 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _819_
timestamp 1688980957
transform 1 0 24840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _820_
timestamp 1688980957
transform -1 0 26220 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _821_
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _822_
timestamp 1688980957
transform 1 0 25392 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _823_
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _824_
timestamp 1688980957
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _825_
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _826_
timestamp 1688980957
transform 1 0 4876 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _827_
timestamp 1688980957
transform 1 0 5060 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _828_
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _829_
timestamp 1688980957
transform 1 0 4784 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _830_
timestamp 1688980957
transform 1 0 4968 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _831_
timestamp 1688980957
transform 1 0 4600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _832_
timestamp 1688980957
transform -1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _833_
timestamp 1688980957
transform 1 0 5152 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _834_
timestamp 1688980957
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _835_
timestamp 1688980957
transform 1 0 5060 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _836_
timestamp 1688980957
transform 1 0 4416 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _837_
timestamp 1688980957
transform 1 0 5152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _838_
timestamp 1688980957
transform 1 0 5888 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _839_
timestamp 1688980957
transform 1 0 5244 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _840_
timestamp 1688980957
transform -1 0 5796 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _841_
timestamp 1688980957
transform -1 0 5612 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _842_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _843_
timestamp 1688980957
transform 1 0 21344 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _844_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13432 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _845_
timestamp 1688980957
transform 1 0 23460 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _846_
timestamp 1688980957
transform 1 0 23368 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _847_
timestamp 1688980957
transform 1 0 23736 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _848_
timestamp 1688980957
transform 1 0 23828 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _849_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _850_
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _851_
timestamp 1688980957
transform 1 0 23920 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _852_
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _853_
timestamp 1688980957
transform 1 0 24104 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _854_
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _855_
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _856_
timestamp 1688980957
transform 1 0 21896 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _857_
timestamp 1688980957
transform 1 0 23828 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _858_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3956 0 1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _859_
timestamp 1688980957
transform 1 0 3864 0 1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _860_
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _861_
timestamp 1688980957
transform 1 0 3864 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _862_
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _863_
timestamp 1688980957
transform 1 0 3956 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _864_
timestamp 1688980957
transform 1 0 3864 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _865_
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _866_
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _867_
timestamp 1688980957
transform 1 0 4232 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _868_
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _869_
timestamp 1688980957
transform 1 0 3864 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _870_
timestamp 1688980957
transform 1 0 4140 0 1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _871_
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _872_
timestamp 1688980957
transform 1 0 4232 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _873_
timestamp 1688980957
transform 1 0 4140 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _874_
timestamp 1688980957
transform 1 0 4048 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA__415__A pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__429__B1
timestamp 1688980957
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__439__B1
timestamp 1688980957
transform -1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__442__A1
timestamp 1688980957
transform -1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__465__A1
timestamp 1688980957
transform 1 0 21620 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__492__A1
timestamp 1688980957
transform -1 0 22816 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__528__A1
timestamp 1688980957
transform 1 0 22172 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__549__B
timestamp 1688980957
transform -1 0 10396 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__562__A1
timestamp 1688980957
transform 1 0 22264 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__C
timestamp 1688980957
transform 1 0 9844 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__585__D_N
timestamp 1688980957
transform 1 0 10488 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__A2_N
timestamp 1688980957
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__586__B1
timestamp 1688980957
transform -1 0 6348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__606__A1
timestamp 1688980957
transform 1 0 23000 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__620__B
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__A2
timestamp 1688980957
transform -1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__622__B1
timestamp 1688980957
transform -1 0 9844 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__624__A3
timestamp 1688980957
transform 1 0 9292 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__640__A1
timestamp 1688980957
transform 1 0 23276 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__A2_N
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__658__B1
timestamp 1688980957
transform 1 0 13432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__659__A2
timestamp 1688980957
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__679__A1
timestamp 1688980957
transform 1 0 22540 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__A2
timestamp 1688980957
transform 1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__687__B1
timestamp 1688980957
transform 1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__699__B
timestamp 1688980957
transform 1 0 12420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__710__A1
timestamp 1688980957
transform 1 0 22448 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__714__C1
timestamp 1688980957
transform -1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__726__C
timestamp 1688980957
transform -1 0 9936 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__726__D_N
timestamp 1688980957
transform 1 0 9936 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__727__A2_N
timestamp 1688980957
transform 1 0 11040 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__727__B1
timestamp 1688980957
transform 1 0 10120 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__741__A
timestamp 1688980957
transform -1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__742__B
timestamp 1688980957
transform -1 0 16836 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__744__C_N
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__760__A1
timestamp 1688980957
transform 1 0 21988 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__761__B
timestamp 1688980957
transform -1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__762__B
timestamp 1688980957
transform 1 0 15640 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__763__A1
timestamp 1688980957
transform 1 0 15272 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__782__A2
timestamp 1688980957
transform -1 0 15272 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__782__C1
timestamp 1688980957
transform 1 0 14720 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__787__B1
timestamp 1688980957
transform -1 0 15088 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__789__A1
timestamp 1688980957
transform -1 0 22816 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__791__A1
timestamp 1688980957
transform -1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__807__A
timestamp 1688980957
transform 1 0 20516 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__807__B
timestamp 1688980957
transform 1 0 21160 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__810__A
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__811__A
timestamp 1688980957
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__812__A
timestamp 1688980957
transform 1 0 24932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__813__A
timestamp 1688980957
transform 1 0 24840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__814__A
timestamp 1688980957
transform 1 0 26036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__815__A
timestamp 1688980957
transform 1 0 26128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__816__A
timestamp 1688980957
transform 1 0 25208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__817__A
timestamp 1688980957
transform 1 0 25392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__818__A
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__819__A
timestamp 1688980957
transform 1 0 25300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__820__A
timestamp 1688980957
transform 1 0 26404 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__821__A
timestamp 1688980957
transform 1 0 25852 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__822__A
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__823__A
timestamp 1688980957
transform 1 0 23368 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__824__A
timestamp 1688980957
transform 1 0 24288 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__825__A
timestamp 1688980957
transform 1 0 5428 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__826__A
timestamp 1688980957
transform 1 0 5336 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__827__A
timestamp 1688980957
transform 1 0 5520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__828__A
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__829__A
timestamp 1688980957
transform 1 0 5244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__830__A
timestamp 1688980957
transform 1 0 4784 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__831__A
timestamp 1688980957
transform 1 0 4416 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__832__A
timestamp 1688980957
transform 1 0 5980 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__833__A
timestamp 1688980957
transform 1 0 5612 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__834__A
timestamp 1688980957
transform 1 0 5612 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__835__A
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__836__A
timestamp 1688980957
transform -1 0 4416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__837__A
timestamp 1688980957
transform 1 0 5612 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__838__A
timestamp 1688980957
transform 1 0 6532 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__839__A
timestamp 1688980957
transform 1 0 6348 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__840__A
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__841__A
timestamp 1688980957
transform 1 0 5796 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__842__CLK
timestamp 1688980957
transform 1 0 20424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__842__D
timestamp 1688980957
transform -1 0 20792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__843__CLK
timestamp 1688980957
transform 1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__844__CLK
timestamp 1688980957
transform 1 0 13248 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__845__CLK
timestamp 1688980957
transform 1 0 23276 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__846__CLK
timestamp 1688980957
transform 1 0 23184 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__847__CLK
timestamp 1688980957
transform 1 0 23552 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__848__CLK
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__849__CLK
timestamp 1688980957
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__850__CLK
timestamp 1688980957
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__851__CLK
timestamp 1688980957
transform 1 0 23736 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__852__CLK
timestamp 1688980957
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__853__CLK
timestamp 1688980957
transform 1 0 23920 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__854__CLK
timestamp 1688980957
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__855__CLK
timestamp 1688980957
transform 1 0 23828 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__856__CLK
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__857__CLK
timestamp 1688980957
transform -1 0 23828 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__858__CLK
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__859__CLK
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__860__CLK
timestamp 1688980957
transform 1 0 6348 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__861__CLK
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__862__CLK
timestamp 1688980957
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__863__CLK
timestamp 1688980957
transform 1 0 6072 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__864__CLK
timestamp 1688980957
transform 1 0 6532 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__865__CLK
timestamp 1688980957
transform 1 0 5520 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__866__CLK
timestamp 1688980957
transform 1 0 6440 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__867__CLK
timestamp 1688980957
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__868__CLK
timestamp 1688980957
transform 1 0 6164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__869__CLK
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__870__CLK
timestamp 1688980957
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__871__CLK
timestamp 1688980957
transform 1 0 7176 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__872__CLK
timestamp 1688980957
transform 1 0 6532 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__873__CLK
timestamp 1688980957
transform 1 0 6440 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__874__CLK
timestamp 1688980957
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_A
timestamp 1688980957
transform 1 0 32936 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_99
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_281 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_301 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_211
timestamp 1688980957
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_214
timestamp 1688980957
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_222
timestamp 1688980957
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_367
timestamp 1688980957
transform 1 0 34868 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_212
timestamp 1688980957
transform 1 0 20608 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_237
timestamp 1688980957
transform 1 0 22908 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_241
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 24012 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_367
timestamp 1688980957
transform 1 0 34868 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_18
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_367
timestamp 1688980957
transform 1 0 34868 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_217
timestamp 1688980957
transform 1 0 21068 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_243
timestamp 1688980957
transform 1 0 23460 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_247
timestamp 1688980957
transform 1 0 23828 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_367
timestamp 1688980957
transform 1 0 34868 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 1688980957
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1688980957
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1688980957
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_367
timestamp 1688980957
transform 1 0 34868 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_49
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_367
timestamp 1688980957
transform 1 0 34868 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 1688980957
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1688980957
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_54
timestamp 1688980957
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_58
timestamp 1688980957
transform 1 0 6440 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_70
timestamp 1688980957
transform 1 0 7544 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_367
timestamp 1688980957
transform 1 0 34868 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_147
timestamp 1688980957
transform 1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_151
timestamp 1688980957
transform 1 0 14996 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_163
timestamp 1688980957
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_175
timestamp 1688980957
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_187
timestamp 1688980957
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_43
timestamp 1688980957
transform 1 0 5060 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_47
timestamp 1688980957
transform 1 0 5428 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_131
timestamp 1688980957
transform 1 0 13156 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_155
timestamp 1688980957
transform 1 0 15364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_263
timestamp 1688980957
transform 1 0 25300 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_275
timestamp 1688980957
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_367
timestamp 1688980957
transform 1 0 34868 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_6
timestamp 1688980957
transform 1 0 1656 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_18
timestamp 1688980957
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_26
timestamp 1688980957
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_33
timestamp 1688980957
transform 1 0 4140 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_57
timestamp 1688980957
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_61
timestamp 1688980957
transform 1 0 6716 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_73
timestamp 1688980957
transform 1 0 7820 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_126
timestamp 1688980957
transform 1 0 12696 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_257
timestamp 1688980957
transform 1 0 24748 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_273
timestamp 1688980957
transform 1 0 26220 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_285
timestamp 1688980957
transform 1 0 27324 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_297
timestamp 1688980957
transform 1 0 28428 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 1688980957
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_47
timestamp 1688980957
transform 1 0 5428 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_126
timestamp 1688980957
transform 1 0 12696 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_138
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_150
timestamp 1688980957
transform 1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_159
timestamp 1688980957
transform 1 0 15732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_175
timestamp 1688980957
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_179
timestamp 1688980957
transform 1 0 17572 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_191
timestamp 1688980957
transform 1 0 18676 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_203
timestamp 1688980957
transform 1 0 19780 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_213
timestamp 1688980957
transform 1 0 20700 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_221
timestamp 1688980957
transform 1 0 21436 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_233
timestamp 1688980957
transform 1 0 22540 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_239
timestamp 1688980957
transform 1 0 23092 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_262
timestamp 1688980957
transform 1 0 25208 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_274
timestamp 1688980957
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_367
timestamp 1688980957
transform 1 0 34868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_56
timestamp 1688980957
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_60
timestamp 1688980957
transform 1 0 6624 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_72
timestamp 1688980957
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_103
timestamp 1688980957
transform 1 0 10580 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_107
timestamp 1688980957
transform 1 0 10948 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_127
timestamp 1688980957
transform 1 0 12788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_174
timestamp 1688980957
transform 1 0 17112 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_183
timestamp 1688980957
transform 1 0 17940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_205
timestamp 1688980957
transform 1 0 19964 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_216
timestamp 1688980957
transform 1 0 20976 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_220
timestamp 1688980957
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_256
timestamp 1688980957
transform 1 0 24656 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_260
timestamp 1688980957
transform 1 0 25024 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_272
timestamp 1688980957
transform 1 0 26128 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_284
timestamp 1688980957
transform 1 0 27232 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_296
timestamp 1688980957
transform 1 0 28336 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_46
timestamp 1688980957
transform 1 0 5336 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_50
timestamp 1688980957
transform 1 0 5704 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_65
timestamp 1688980957
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_88
timestamp 1688980957
transform 1 0 9200 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_96
timestamp 1688980957
transform 1 0 9936 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_116
timestamp 1688980957
transform 1 0 11776 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_122
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_142
timestamp 1688980957
transform 1 0 14168 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_152
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_191
timestamp 1688980957
transform 1 0 18676 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_203
timestamp 1688980957
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_215
timestamp 1688980957
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_235
timestamp 1688980957
transform 1 0 22724 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_247
timestamp 1688980957
transform 1 0 23828 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_259
timestamp 1688980957
transform 1 0 24932 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_271
timestamp 1688980957
transform 1 0 26036 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_367
timestamp 1688980957
transform 1 0 34868 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_6
timestamp 1688980957
transform 1 0 1656 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_18
timestamp 1688980957
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_55
timestamp 1688980957
transform 1 0 6164 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_59
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_137
timestamp 1688980957
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_146
timestamp 1688980957
transform 1 0 14536 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_158
timestamp 1688980957
transform 1 0 15640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_170
timestamp 1688980957
transform 1 0 16744 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_187
timestamp 1688980957
transform 1 0 18308 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_191
timestamp 1688980957
transform 1 0 18676 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_206
timestamp 1688980957
transform 1 0 20056 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_218
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_225
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_232
timestamp 1688980957
transform 1 0 22448 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_236
timestamp 1688980957
transform 1 0 22816 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_248
timestamp 1688980957
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_31
timestamp 1688980957
transform 1 0 3956 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_61
timestamp 1688980957
transform 1 0 6716 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_67
timestamp 1688980957
transform 1 0 7268 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_90
timestamp 1688980957
transform 1 0 9384 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_102
timestamp 1688980957
transform 1 0 10488 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_109
timestamp 1688980957
transform 1 0 11132 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_123
timestamp 1688980957
transform 1 0 12420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_151
timestamp 1688980957
transform 1 0 14996 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_159
timestamp 1688980957
transform 1 0 15732 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_189
timestamp 1688980957
transform 1 0 18492 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_222
timestamp 1688980957
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_232
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_240
timestamp 1688980957
transform 1 0 23184 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_269
timestamp 1688980957
transform 1 0 25852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_367
timestamp 1688980957
transform 1 0 34868 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_57
timestamp 1688980957
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_61
timestamp 1688980957
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_71
timestamp 1688980957
transform 1 0 7636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_99
timestamp 1688980957
transform 1 0 10212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_116
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_125
timestamp 1688980957
transform 1 0 12604 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_167
timestamp 1688980957
transform 1 0 16468 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_179
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_191
timestamp 1688980957
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_206
timestamp 1688980957
transform 1 0 20056 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_220
timestamp 1688980957
transform 1 0 21344 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_228
timestamp 1688980957
transform 1 0 22080 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_235
timestamp 1688980957
transform 1 0 22724 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_247
timestamp 1688980957
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_31
timestamp 1688980957
transform 1 0 3956 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_91
timestamp 1688980957
transform 1 0 9476 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_95
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_158
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_172
timestamp 1688980957
transform 1 0 16928 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_188
timestamp 1688980957
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_203
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_215
timestamp 1688980957
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_367
timestamp 1688980957
transform 1 0 34868 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_6
timestamp 1688980957
transform 1 0 1656 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_18
timestamp 1688980957
transform 1 0 2760 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1688980957
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_66
timestamp 1688980957
transform 1 0 7176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_70
timestamp 1688980957
transform 1 0 7544 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_81
timestamp 1688980957
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_134
timestamp 1688980957
transform 1 0 13432 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_168
timestamp 1688980957
transform 1 0 16560 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_172
timestamp 1688980957
transform 1 0 16928 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_184
timestamp 1688980957
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_213
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_217
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_229
timestamp 1688980957
transform 1 0 22172 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_232
timestamp 1688980957
transform 1 0 22448 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_244
timestamp 1688980957
transform 1 0 23552 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_33
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_79
timestamp 1688980957
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_100
timestamp 1688980957
transform 1 0 10304 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_138
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_146
timestamp 1688980957
transform 1 0 14536 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_160
timestamp 1688980957
transform 1 0 15824 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_172
timestamp 1688980957
transform 1 0 16928 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_184
timestamp 1688980957
transform 1 0 18032 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_196
timestamp 1688980957
transform 1 0 19136 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_270
timestamp 1688980957
transform 1 0 25944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_274
timestamp 1688980957
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_367
timestamp 1688980957
transform 1 0 34868 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_106
timestamp 1688980957
transform 1 0 10856 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_118
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_128
timestamp 1688980957
transform 1 0 12880 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 14444 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_157
timestamp 1688980957
transform 1 0 15548 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_204
timestamp 1688980957
transform 1 0 19872 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_212
timestamp 1688980957
transform 1 0 20608 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_219
timestamp 1688980957
transform 1 0 21252 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_231
timestamp 1688980957
transform 1 0 22356 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_243
timestamp 1688980957
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_44
timestamp 1688980957
transform 1 0 5152 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_48
timestamp 1688980957
transform 1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_52
timestamp 1688980957
transform 1 0 5888 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_96
timestamp 1688980957
transform 1 0 9936 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_108
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_126
timestamp 1688980957
transform 1 0 12696 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_130
timestamp 1688980957
transform 1 0 13064 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_139
timestamp 1688980957
transform 1 0 13892 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_147
timestamp 1688980957
transform 1 0 14628 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_154
timestamp 1688980957
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_195
timestamp 1688980957
transform 1 0 19044 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_207
timestamp 1688980957
transform 1 0 20148 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_228
timestamp 1688980957
transform 1 0 22080 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_236
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_240
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_252
timestamp 1688980957
transform 1 0 24288 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_256
timestamp 1688980957
transform 1 0 24656 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_260
timestamp 1688980957
transform 1 0 25024 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_264
timestamp 1688980957
transform 1 0 25392 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_276
timestamp 1688980957
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_367
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_6
timestamp 1688980957
transform 1 0 1656 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_18
timestamp 1688980957
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1688980957
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_79
timestamp 1688980957
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_92
timestamp 1688980957
transform 1 0 9568 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_110
timestamp 1688980957
transform 1 0 11224 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_125
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1688980957
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_146
timestamp 1688980957
transform 1 0 14536 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_152
timestamp 1688980957
transform 1 0 15088 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_161
timestamp 1688980957
transform 1 0 15916 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_173
timestamp 1688980957
transform 1 0 17020 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_185
timestamp 1688980957
transform 1 0 18124 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_205
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_246
timestamp 1688980957
transform 1 0 23736 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_273
timestamp 1688980957
transform 1 0 26220 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_285
timestamp 1688980957
transform 1 0 27324 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_297
timestamp 1688980957
transform 1 0 28428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_305
timestamp 1688980957
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_44
timestamp 1688980957
transform 1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_52
timestamp 1688980957
transform 1 0 5888 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_79
timestamp 1688980957
transform 1 0 8372 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_98
timestamp 1688980957
transform 1 0 10120 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_132
timestamp 1688980957
transform 1 0 13248 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_162
timestamp 1688980957
transform 1 0 16008 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_183
timestamp 1688980957
transform 1 0 17940 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_195
timestamp 1688980957
transform 1 0 19044 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_207
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_219
timestamp 1688980957
transform 1 0 21252 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_367
timestamp 1688980957
transform 1 0 34868 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_145
timestamp 1688980957
transform 1 0 14444 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_161
timestamp 1688980957
transform 1 0 15916 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_176
timestamp 1688980957
transform 1 0 17296 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_183
timestamp 1688980957
transform 1 0 17940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_207
timestamp 1688980957
transform 1 0 20148 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_217
timestamp 1688980957
transform 1 0 21068 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_229
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_241
timestamp 1688980957
transform 1 0 23276 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_249
timestamp 1688980957
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_47
timestamp 1688980957
transform 1 0 5428 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_92
timestamp 1688980957
transform 1 0 9568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_104
timestamp 1688980957
transform 1 0 10672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_140
timestamp 1688980957
transform 1 0 13984 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_152
timestamp 1688980957
transform 1 0 15088 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_164
timestamp 1688980957
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_187
timestamp 1688980957
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_206
timestamp 1688980957
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_218
timestamp 1688980957
transform 1 0 21160 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_367
timestamp 1688980957
transform 1 0 34868 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_6
timestamp 1688980957
transform 1 0 1656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_18
timestamp 1688980957
transform 1 0 2760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 1688980957
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_95
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_119
timestamp 1688980957
transform 1 0 12052 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1688980957
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_154
timestamp 1688980957
transform 1 0 15272 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_166
timestamp 1688980957
transform 1 0 16376 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_174
timestamp 1688980957
transform 1 0 17112 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_186
timestamp 1688980957
transform 1 0 18216 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_194
timestamp 1688980957
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_202
timestamp 1688980957
transform 1 0 19688 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_214
timestamp 1688980957
transform 1 0 20792 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_226
timestamp 1688980957
transform 1 0 21896 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_238
timestamp 1688980957
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_250
timestamp 1688980957
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_79
timestamp 1688980957
transform 1 0 8372 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_83
timestamp 1688980957
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_92
timestamp 1688980957
transform 1 0 9568 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_107
timestamp 1688980957
transform 1 0 10948 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_121
timestamp 1688980957
transform 1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_132
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_144
timestamp 1688980957
transform 1 0 14352 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_152
timestamp 1688980957
transform 1 0 15088 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_177
timestamp 1688980957
transform 1 0 17388 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_188
timestamp 1688980957
transform 1 0 18400 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_196
timestamp 1688980957
transform 1 0 19136 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_203
timestamp 1688980957
transform 1 0 19780 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_215
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 1688980957
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_257
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_262
timestamp 1688980957
transform 1 0 25208 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_266
timestamp 1688980957
transform 1 0 25576 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_278
timestamp 1688980957
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_367
timestamp 1688980957
transform 1 0 34868 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_43
timestamp 1688980957
transform 1 0 5060 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_47
timestamp 1688980957
transform 1 0 5428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_55
timestamp 1688980957
transform 1 0 6164 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_71
timestamp 1688980957
transform 1 0 7636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_93
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_112
timestamp 1688980957
transform 1 0 11408 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_124
timestamp 1688980957
transform 1 0 12512 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_147
timestamp 1688980957
transform 1 0 14628 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_158
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_167
timestamp 1688980957
transform 1 0 16468 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_179
timestamp 1688980957
transform 1 0 17572 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_192
timestamp 1688980957
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_213
timestamp 1688980957
transform 1 0 20700 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_225
timestamp 1688980957
transform 1 0 21804 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_241
timestamp 1688980957
transform 1 0 23276 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_273
timestamp 1688980957
transform 1 0 26220 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_285
timestamp 1688980957
transform 1 0 27324 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_297
timestamp 1688980957
transform 1 0 28428 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_305
timestamp 1688980957
transform 1 0 29164 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_52
timestamp 1688980957
transform 1 0 5888 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_65
timestamp 1688980957
transform 1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_89
timestamp 1688980957
transform 1 0 9292 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_134
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_160
timestamp 1688980957
transform 1 0 15824 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_187
timestamp 1688980957
transform 1 0 18308 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_199
timestamp 1688980957
transform 1 0 19412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_211
timestamp 1688980957
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_239
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_243
timestamp 1688980957
transform 1 0 23460 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_255
timestamp 1688980957
transform 1 0 24564 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_267
timestamp 1688980957
transform 1 0 25668 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1688980957
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_367
timestamp 1688980957
transform 1 0 34868 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_6
timestamp 1688980957
transform 1 0 1656 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_18
timestamp 1688980957
transform 1 0 2760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_26
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_79
timestamp 1688980957
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_114
timestamp 1688980957
transform 1 0 11592 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_130
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_134
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_147
timestamp 1688980957
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_156
timestamp 1688980957
transform 1 0 15456 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_162
timestamp 1688980957
transform 1 0 16008 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_167
timestamp 1688980957
transform 1 0 16468 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_179
timestamp 1688980957
transform 1 0 17572 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_185
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_190
timestamp 1688980957
transform 1 0 18584 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_203
timestamp 1688980957
transform 1 0 19780 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_215
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_222
timestamp 1688980957
transform 1 0 21528 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_230
timestamp 1688980957
transform 1 0 22264 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_243
timestamp 1688980957
transform 1 0 23460 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_65
timestamp 1688980957
transform 1 0 7084 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_103
timestamp 1688980957
transform 1 0 10580 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_143
timestamp 1688980957
transform 1 0 14260 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_177
timestamp 1688980957
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_196
timestamp 1688980957
transform 1 0 19136 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_203
timestamp 1688980957
transform 1 0 19780 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_215
timestamp 1688980957
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_243
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_271
timestamp 1688980957
transform 1 0 26036 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_275
timestamp 1688980957
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_367
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_37
timestamp 1688980957
transform 1 0 4508 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_45
timestamp 1688980957
transform 1 0 5244 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_50
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_56
timestamp 1688980957
transform 1 0 6256 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_69
timestamp 1688980957
transform 1 0 7452 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_79
timestamp 1688980957
transform 1 0 8372 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_113
timestamp 1688980957
transform 1 0 11500 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_134
timestamp 1688980957
transform 1 0 13432 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_160
timestamp 1688980957
transform 1 0 15824 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_175
timestamp 1688980957
transform 1 0 17204 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_187
timestamp 1688980957
transform 1 0 18308 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_208
timestamp 1688980957
transform 1 0 20240 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_217
timestamp 1688980957
transform 1 0 21068 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_224
timestamp 1688980957
transform 1 0 21712 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_234
timestamp 1688980957
transform 1 0 22632 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_246
timestamp 1688980957
transform 1 0 23736 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1688980957
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_88
timestamp 1688980957
transform 1 0 9200 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_124
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_134
timestamp 1688980957
transform 1 0 13432 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_140
timestamp 1688980957
transform 1 0 13984 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_152
timestamp 1688980957
transform 1 0 15088 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_164
timestamp 1688980957
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_209
timestamp 1688980957
transform 1 0 20332 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_221
timestamp 1688980957
transform 1 0 21436 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_232
timestamp 1688980957
transform 1 0 22448 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_248
timestamp 1688980957
transform 1 0 23920 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_256
timestamp 1688980957
transform 1 0 24656 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_265
timestamp 1688980957
transform 1 0 25484 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_277
timestamp 1688980957
transform 1 0 26588 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_367
timestamp 1688980957
transform 1 0 34868 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_6
timestamp 1688980957
transform 1 0 1656 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_18
timestamp 1688980957
transform 1 0 2760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_26
timestamp 1688980957
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_56
timestamp 1688980957
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_92
timestamp 1688980957
transform 1 0 9568 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_104
timestamp 1688980957
transform 1 0 10672 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_108
timestamp 1688980957
transform 1 0 11040 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_128
timestamp 1688980957
transform 1 0 12880 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_146
timestamp 1688980957
transform 1 0 14536 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_152
timestamp 1688980957
transform 1 0 15088 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_156
timestamp 1688980957
transform 1 0 15456 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_160
timestamp 1688980957
transform 1 0 15824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_168
timestamp 1688980957
transform 1 0 16560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_180
timestamp 1688980957
transform 1 0 17664 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_249
timestamp 1688980957
transform 1 0 24012 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_273
timestamp 1688980957
transform 1 0 26220 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_285
timestamp 1688980957
transform 1 0 27324 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_297
timestamp 1688980957
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_305
timestamp 1688980957
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_43
timestamp 1688980957
transform 1 0 5060 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_47
timestamp 1688980957
transform 1 0 5428 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_101
timestamp 1688980957
transform 1 0 10396 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_106
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1688980957
transform 1 0 11224 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_121
timestamp 1688980957
transform 1 0 12236 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_128
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_150
timestamp 1688980957
transform 1 0 14904 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_221
timestamp 1688980957
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_367
timestamp 1688980957
transform 1 0 34868 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_56
timestamp 1688980957
transform 1 0 6256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_60
timestamp 1688980957
transform 1 0 6624 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_93
timestamp 1688980957
transform 1 0 9660 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_96
timestamp 1688980957
transform 1 0 9936 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_128
timestamp 1688980957
transform 1 0 12880 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_147
timestamp 1688980957
transform 1 0 14628 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_150
timestamp 1688980957
transform 1 0 14904 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_167
timestamp 1688980957
transform 1 0 16468 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_171
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_179
timestamp 1688980957
transform 1 0 17572 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1688980957
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_201
timestamp 1688980957
transform 1 0 19596 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_227
timestamp 1688980957
transform 1 0 21988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_235
timestamp 1688980957
transform 1 0 22724 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_246
timestamp 1688980957
transform 1 0 23736 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_33
timestamp 1688980957
transform 1 0 4140 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_61
timestamp 1688980957
transform 1 0 6716 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_73
timestamp 1688980957
transform 1 0 7820 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_85
timestamp 1688980957
transform 1 0 8924 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_98
timestamp 1688980957
transform 1 0 10120 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_102
timestamp 1688980957
transform 1 0 10488 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_108
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_119
timestamp 1688980957
transform 1 0 12052 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_134
timestamp 1688980957
transform 1 0 13432 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_144
timestamp 1688980957
transform 1 0 14352 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_152
timestamp 1688980957
transform 1 0 15088 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_162
timestamp 1688980957
transform 1 0 16008 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_173
timestamp 1688980957
transform 1 0 17020 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_211
timestamp 1688980957
transform 1 0 20516 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_220
timestamp 1688980957
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_246
timestamp 1688980957
transform 1 0 23736 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_277
timestamp 1688980957
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 1688980957
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_367
timestamp 1688980957
transform 1 0 34868 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_6
timestamp 1688980957
transform 1 0 1656 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_18
timestamp 1688980957
transform 1 0 2760 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_26
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_51
timestamp 1688980957
transform 1 0 5796 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_55
timestamp 1688980957
transform 1 0 6164 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_59
timestamp 1688980957
transform 1 0 6532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_71
timestamp 1688980957
transform 1 0 7636 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_118
timestamp 1688980957
transform 1 0 11960 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_125
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1688980957
transform 1 0 13708 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_145
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_160
timestamp 1688980957
transform 1 0 15824 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_171
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_179
timestamp 1688980957
transform 1 0 17572 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_185
timestamp 1688980957
transform 1 0 18124 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1688980957
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_239
timestamp 1688980957
transform 1 0 23092 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_247
timestamp 1688980957
transform 1 0 23828 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_273
timestamp 1688980957
transform 1 0 26220 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_285
timestamp 1688980957
transform 1 0 27324 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_297
timestamp 1688980957
transform 1 0 28428 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_305
timestamp 1688980957
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_53
timestamp 1688980957
transform 1 0 5980 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_61
timestamp 1688980957
transform 1 0 6716 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_73
timestamp 1688980957
transform 1 0 7820 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_85
timestamp 1688980957
transform 1 0 8924 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_97
timestamp 1688980957
transform 1 0 10028 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_109
timestamp 1688980957
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_134
timestamp 1688980957
transform 1 0 13432 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_158
timestamp 1688980957
transform 1 0 15640 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_166
timestamp 1688980957
transform 1 0 16376 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_189
timestamp 1688980957
transform 1 0 18492 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_222
timestamp 1688980957
transform 1 0 21528 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_232
timestamp 1688980957
transform 1 0 22448 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_236
timestamp 1688980957
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_254
timestamp 1688980957
transform 1 0 24472 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_260
timestamp 1688980957
transform 1 0 25024 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_267
timestamp 1688980957
transform 1 0 25668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_271
timestamp 1688980957
transform 1 0 26036 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_275
timestamp 1688980957
transform 1 0 26404 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_367
timestamp 1688980957
transform 1 0 34868 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_35
timestamp 1688980957
transform 1 0 4324 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_68
timestamp 1688980957
transform 1 0 7360 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_80
timestamp 1688980957
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_132
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_144
timestamp 1688980957
transform 1 0 14352 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_150
timestamp 1688980957
transform 1 0 14904 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_162
timestamp 1688980957
transform 1 0 16008 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_174
timestamp 1688980957
transform 1 0 17112 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_186
timestamp 1688980957
transform 1 0 18216 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_190
timestamp 1688980957
transform 1 0 18584 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_204
timestamp 1688980957
transform 1 0 19872 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_216
timestamp 1688980957
transform 1 0 20976 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_235
timestamp 1688980957
transform 1 0 22724 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_240
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_244
timestamp 1688980957
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_273
timestamp 1688980957
transform 1 0 26220 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_285
timestamp 1688980957
transform 1 0 27324 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_297
timestamp 1688980957
transform 1 0 28428 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_305
timestamp 1688980957
transform 1 0 29164 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_61
timestamp 1688980957
transform 1 0 6716 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_73
timestamp 1688980957
transform 1 0 7820 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_85
timestamp 1688980957
transform 1 0 8924 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_97
timestamp 1688980957
transform 1 0 10028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_109
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_221
timestamp 1688980957
transform 1 0 21436 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_268
timestamp 1688980957
transform 1 0 25760 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_367
timestamp 1688980957
transform 1 0 34868 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_6
timestamp 1688980957
transform 1 0 1656 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_18
timestamp 1688980957
transform 1 0 2760 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_247
timestamp 1688980957
transform 1 0 23828 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_367
timestamp 1688980957
transform 1 0 34868 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_367
timestamp 1688980957
transform 1 0 34868 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_6
timestamp 1688980957
transform 1 0 1656 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_18
timestamp 1688980957
transform 1 0 2760 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_367
timestamp 1688980957
transform 1 0 34868 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_367
timestamp 1688980957
transform 1 0 34868 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_6
timestamp 1688980957
transform 1 0 1656 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_18
timestamp 1688980957
transform 1 0 2760 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_26
timestamp 1688980957
transform 1 0 3496 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_367
timestamp 1688980957
transform 1 0 34868 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_367
timestamp 1688980957
transform 1 0 34868 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_6
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_18
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 1688980957
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_367
timestamp 1688980957
transform 1 0 34868 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_6
timestamp 1688980957
transform 1 0 1656 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_18
timestamp 1688980957
transform 1 0 2760 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_69
timestamp 1688980957
transform 1 0 7452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_81
timestamp 1688980957
transform 1 0 8556 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_113
timestamp 1688980957
transform 1 0 11500 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_125
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_169
timestamp 1688980957
transform 1 0 16652 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_181
timestamp 1688980957
transform 1 0 17756 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_225
timestamp 1688980957
transform 1 0 21804 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_237
timestamp 1688980957
transform 1 0 22908 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_249
timestamp 1688980957
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_281
timestamp 1688980957
transform 1 0 26956 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_293
timestamp 1688980957
transform 1 0 28060 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_305
timestamp 1688980957
transform 1 0 29164 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_337
timestamp 1688980957
transform 1 0 32108 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 1656 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform -1 0 1656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform -1 0 1656 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform -1 0 1656 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input17 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  input19 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27324 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output20
timestamp 1688980957
transform 1 0 33120 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 1688980957
transform 1 0 33120 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 1688980957
transform 1 0 33120 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 1688980957
transform 1 0 33120 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 1688980957
transform 1 0 33120 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 1688980957
transform 1 0 33120 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 1688980957
transform 1 0 33120 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 1688980957
transform 1 0 33120 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 1688980957
transform 1 0 33120 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 1688980957
transform 1 0 33120 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 1688980957
transform 1 0 33120 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 1688980957
transform 1 0 33120 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 1688980957
transform 1 0 33120 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 1688980957
transform 1 0 33120 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output35
timestamp 1688980957
transform 1 0 33120 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 35236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 35236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 35236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 35236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 35236 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 35236 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 35236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 35236 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 35236 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 35236 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 35236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 35236 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 35236 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 35236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 35236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 35236 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 35236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 35236 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 35236 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 35236 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 35236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 35236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 35236 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 35236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 35236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 35236 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 35236 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 35236 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 35236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 35236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 35236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 35236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 35236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 35236 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 35236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 35236 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 35236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 35236 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 35236 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 35236 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 35236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 35236 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 35236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 35236 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 35236 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 35236 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 35236 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 35236 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 35236 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 35236 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 35236 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 35236 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 35236 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 35236 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 35236 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 35236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 35236 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 35236 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 6256 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 11408 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 21712 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 26864 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 32016 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
<< labels >>
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 a[0]
port 0 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 a[1]
port 1 nsew signal input
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 a[2]
port 2 nsew signal input
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 a[3]
port 3 nsew signal input
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 a[4]
port 4 nsew signal input
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 a[5]
port 5 nsew signal input
flabel metal3 s 0 30200 800 30320 0 FreeSans 480 0 0 0 a[6]
port 6 nsew signal input
flabel metal3 s 0 34552 800 34672 0 FreeSans 480 0 0 0 a[7]
port 7 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 b[0]
port 8 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 b[1]
port 9 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 b[2]
port 10 nsew signal input
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 b[3]
port 11 nsew signal input
flabel metal3 s 0 23672 800 23792 0 FreeSans 480 0 0 0 b[4]
port 12 nsew signal input
flabel metal3 s 0 28024 800 28144 0 FreeSans 480 0 0 0 b[5]
port 13 nsew signal input
flabel metal3 s 0 32376 800 32496 0 FreeSans 480 0 0 0 b[6]
port 14 nsew signal input
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 b[7]
port 15 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 clk
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 control
port 17 nsew signal input
flabel metal3 s 35600 3000 36400 3120 0 FreeSans 480 0 0 0 p[0]
port 18 nsew signal tristate
flabel metal3 s 35600 24760 36400 24880 0 FreeSans 480 0 0 0 p[10]
port 19 nsew signal tristate
flabel metal3 s 35600 26936 36400 27056 0 FreeSans 480 0 0 0 p[11]
port 20 nsew signal tristate
flabel metal3 s 35600 29112 36400 29232 0 FreeSans 480 0 0 0 p[12]
port 21 nsew signal tristate
flabel metal3 s 35600 31288 36400 31408 0 FreeSans 480 0 0 0 p[13]
port 22 nsew signal tristate
flabel metal3 s 35600 33464 36400 33584 0 FreeSans 480 0 0 0 p[14]
port 23 nsew signal tristate
flabel metal3 s 35600 35640 36400 35760 0 FreeSans 480 0 0 0 p[15]
port 24 nsew signal tristate
flabel metal3 s 35600 5176 36400 5296 0 FreeSans 480 0 0 0 p[1]
port 25 nsew signal tristate
flabel metal3 s 35600 7352 36400 7472 0 FreeSans 480 0 0 0 p[2]
port 26 nsew signal tristate
flabel metal3 s 35600 9528 36400 9648 0 FreeSans 480 0 0 0 p[3]
port 27 nsew signal tristate
flabel metal3 s 35600 11704 36400 11824 0 FreeSans 480 0 0 0 p[4]
port 28 nsew signal tristate
flabel metal3 s 35600 13880 36400 14000 0 FreeSans 480 0 0 0 p[5]
port 29 nsew signal tristate
flabel metal3 s 35600 16056 36400 16176 0 FreeSans 480 0 0 0 p[6]
port 30 nsew signal tristate
flabel metal3 s 35600 18232 36400 18352 0 FreeSans 480 0 0 0 p[7]
port 31 nsew signal tristate
flabel metal3 s 35600 20408 36400 20528 0 FreeSans 480 0 0 0 p[8]
port 32 nsew signal tristate
flabel metal3 s 35600 22584 36400 22704 0 FreeSans 480 0 0 0 p[9]
port 33 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 rst
port 34 nsew signal input
flabel metal4 s 4208 2128 4528 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 34928 2128 35248 36496 0 FreeSans 1920 90 0 0 vccd1
port 35 nsew power bidirectional
flabel metal4 s 19568 2128 19888 36496 0 FreeSans 1920 90 0 0 vssd1
port 36 nsew ground bidirectional
rlabel metal1 18176 36448 18176 36448 0 vccd1
rlabel metal1 18170 35904 18170 35904 0 vssd1
rlabel metal1 10856 12206 10856 12206 0 FA0.q
rlabel metal2 8050 19142 8050 19142 0 FA1.q
rlabel metal2 7130 16014 7130 16014 0 FA2.q
rlabel metal1 6946 18292 6946 18292 0 FA3.q
rlabel metal1 8832 21522 8832 21522 0 FA4.q
rlabel metal2 7958 22848 7958 22848 0 FA5.q
rlabel metal1 6302 21998 6302 21998 0 FA6.q
rlabel metal1 6072 19890 6072 19890 0 FA7.q
rlabel metal1 10718 12172 10718 12172 0 FB0.q
rlabel metal2 7314 12002 7314 12002 0 FB1.q
rlabel metal2 7682 14416 7682 14416 0 FB2.q
rlabel metal2 6854 16320 6854 16320 0 FB3.q
rlabel metal2 8050 23936 8050 23936 0 FB4.q
rlabel metal1 7084 25262 7084 25262 0 FB5.q
rlabel via1 6946 25262 6946 25262 0 FB6.q
rlabel metal1 6716 14994 6716 14994 0 FB7.q
rlabel metal1 6900 20910 6900 20910 0 FC.q
rlabel metal1 20930 3570 20930 3570 0 FP0.d
rlabel metal1 21160 12342 21160 12342 0 FP1.d
rlabel metal1 24288 23630 24288 23630 0 FP10.d
rlabel metal1 23874 25466 23874 25466 0 FP11.d
rlabel metal1 24196 26010 24196 26010 0 FP12.d
rlabel metal1 23552 26894 23552 26894 0 FP13.d
rlabel metal2 22218 27812 22218 27812 0 FP14.d
rlabel metal2 22678 27744 22678 27744 0 FP15.d
rlabel metal1 13202 10710 13202 10710 0 FP2.d
rlabel metal1 23644 10710 23644 10710 0 FP3.d
rlabel metal1 23644 11798 23644 11798 0 FP4.d
rlabel metal1 23138 13906 23138 13906 0 FP5.d
rlabel metal1 23966 16218 23966 16218 0 FP6.d
rlabel metal1 23920 17714 23920 17714 0 FP7.d
rlabel metal1 23966 20978 23966 20978 0 FP8.d
rlabel metal1 23782 22202 23782 22202 0 FP9.d
rlabel metal1 22547 3434 22547 3434 0 _000_
rlabel metal1 23099 5610 23099 5610 0 _001_
rlabel metal2 14490 10472 14490 10472 0 _002_
rlabel metal2 24886 10846 24886 10846 0 _003_
rlabel metal2 24426 11934 24426 11934 0 _004_
rlabel metal1 25491 13974 25491 13974 0 _005_
rlabel metal1 25583 16150 25583 16150 0 _006_
rlabel metal1 25024 17306 25024 17306 0 _007_
rlabel metal1 25116 20570 25116 20570 0 _008_
rlabel metal1 25675 22678 25675 22678 0 _009_
rlabel metal2 24978 23970 24978 23970 0 _010_
rlabel metal1 25859 25942 25859 25942 0 _011_
rlabel metal2 25254 26520 25254 26520 0 _012_
rlabel metal1 25484 27098 25484 27098 0 _013_
rlabel metal1 23000 27574 23000 27574 0 _014_
rlabel metal1 24518 27302 24518 27302 0 _015_
rlabel metal1 5060 8602 5060 8602 0 _016_
rlabel metal1 4968 18394 4968 18394 0 _017_
rlabel metal1 5152 12954 5152 12954 0 _018_
rlabel metal1 4968 17306 4968 17306 0 _019_
rlabel metal1 4876 21114 4876 21114 0 _020_
rlabel metal1 5060 23290 5060 23290 0 _021_
rlabel metal2 4738 27166 4738 27166 0 _022_
rlabel metal1 5389 22678 5389 22678 0 _023_
rlabel metal1 5244 11866 5244 11866 0 _024_
rlabel metal1 5428 10778 5428 10778 0 _025_
rlabel metal1 5152 14586 5152 14586 0 _026_
rlabel metal1 4600 16218 4600 16218 0 _027_
rlabel metal1 5244 24582 5244 24582 0 _028_
rlabel metal1 5980 27846 5980 27846 0 _029_
rlabel metal2 5566 26112 5566 26112 0 _030_
rlabel metal1 5566 25371 5566 25371 0 _031_
rlabel metal2 5474 14076 5474 14076 0 _032_
rlabel metal1 9522 16558 9522 16558 0 _033_
rlabel metal1 14674 14008 14674 14008 0 _034_
rlabel metal1 13846 13906 13846 13906 0 _035_
rlabel metal1 7268 18258 7268 18258 0 _036_
rlabel metal1 14858 14416 14858 14416 0 _037_
rlabel metal1 13570 14314 13570 14314 0 _038_
rlabel metal2 14582 14280 14582 14280 0 _039_
rlabel via2 13478 13923 13478 13923 0 _040_
rlabel metal1 14168 12206 14168 12206 0 _041_
rlabel metal2 14490 11798 14490 11798 0 _042_
rlabel metal1 12650 11764 12650 11764 0 _043_
rlabel metal1 15824 12206 15824 12206 0 _044_
rlabel metal1 16721 12342 16721 12342 0 _045_
rlabel metal1 16882 12784 16882 12784 0 _046_
rlabel metal1 12742 12274 12742 12274 0 _047_
rlabel metal1 15962 11730 15962 11730 0 _048_
rlabel metal2 16790 12002 16790 12002 0 _049_
rlabel metal2 17526 11968 17526 11968 0 _050_
rlabel metal1 17020 11730 17020 11730 0 _051_
rlabel metal1 19734 11662 19734 11662 0 _052_
rlabel metal1 22402 12818 22402 12818 0 _053_
rlabel metal1 7130 15674 7130 15674 0 _054_
rlabel metal1 6854 24310 6854 24310 0 _055_
rlabel metal2 9338 20978 9338 20978 0 _056_
rlabel metal1 11178 24718 11178 24718 0 _057_
rlabel metal1 16100 15402 16100 15402 0 _058_
rlabel metal1 8372 21998 8372 21998 0 _059_
rlabel metal1 7958 21930 7958 21930 0 _060_
rlabel metal1 12742 16626 12742 16626 0 _061_
rlabel metal1 15916 15470 15916 15470 0 _062_
rlabel metal1 16422 15674 16422 15674 0 _063_
rlabel metal1 16652 14994 16652 14994 0 _064_
rlabel metal1 19458 14586 19458 14586 0 _065_
rlabel metal2 15686 14348 15686 14348 0 _066_
rlabel metal1 13616 13158 13616 13158 0 _067_
rlabel metal1 13708 12274 13708 12274 0 _068_
rlabel metal1 13662 12750 13662 12750 0 _069_
rlabel metal1 14444 12342 14444 12342 0 _070_
rlabel metal1 14582 12274 14582 12274 0 _071_
rlabel via1 17158 12206 17158 12206 0 _072_
rlabel metal1 18998 13260 18998 13260 0 _073_
rlabel metal1 19412 13838 19412 13838 0 _074_
rlabel metal1 19734 14348 19734 14348 0 _075_
rlabel metal1 21022 13872 21022 13872 0 _076_
rlabel metal1 22034 13838 22034 13838 0 _077_
rlabel metal1 21528 13294 21528 13294 0 _078_
rlabel metal1 22126 13226 22126 13226 0 _079_
rlabel metal1 22678 13906 22678 13906 0 _080_
rlabel metal1 18722 16524 18722 16524 0 _081_
rlabel metal1 16238 14348 16238 14348 0 _082_
rlabel metal1 17342 13294 17342 13294 0 _083_
rlabel metal1 12972 12886 12972 12886 0 _084_
rlabel metal1 13524 12818 13524 12818 0 _085_
rlabel metal2 16054 13022 16054 13022 0 _086_
rlabel metal1 17710 12716 17710 12716 0 _087_
rlabel metal1 17848 12750 17848 12750 0 _088_
rlabel metal1 18952 13906 18952 13906 0 _089_
rlabel metal1 18446 13906 18446 13906 0 _090_
rlabel metal2 18906 14144 18906 14144 0 _091_
rlabel metal1 20148 14246 20148 14246 0 _092_
rlabel metal1 20240 14382 20240 14382 0 _093_
rlabel metal2 9246 24514 9246 24514 0 _094_
rlabel metal1 9246 20978 9246 20978 0 _095_
rlabel metal1 12558 19380 12558 19380 0 _096_
rlabel metal1 13754 19788 13754 19788 0 _097_
rlabel metal1 13754 19414 13754 19414 0 _098_
rlabel metal1 15456 16082 15456 16082 0 _099_
rlabel metal2 8602 22372 8602 22372 0 _100_
rlabel metal1 9246 16626 9246 16626 0 _101_
rlabel metal2 8786 16966 8786 16966 0 _102_
rlabel metal2 13386 16252 13386 16252 0 _103_
rlabel metal1 13570 16150 13570 16150 0 _104_
rlabel metal1 14536 16082 14536 16082 0 _105_
rlabel metal1 16514 16014 16514 16014 0 _106_
rlabel metal1 15962 16150 15962 16150 0 _107_
rlabel metal1 16836 15470 16836 15470 0 _108_
rlabel metal1 17020 14926 17020 14926 0 _109_
rlabel metal1 18768 14382 18768 14382 0 _110_
rlabel metal1 20424 14382 20424 14382 0 _111_
rlabel metal1 21298 14416 21298 14416 0 _112_
rlabel metal1 21022 15504 21022 15504 0 _113_
rlabel metal1 21942 13906 21942 13906 0 _114_
rlabel metal1 22448 13838 22448 13838 0 _115_
rlabel metal1 22908 16082 22908 16082 0 _116_
rlabel metal1 20424 15470 20424 15470 0 _117_
rlabel metal1 21482 15674 21482 15674 0 _118_
rlabel metal1 15991 14382 15991 14382 0 _119_
rlabel metal1 15502 13974 15502 13974 0 _120_
rlabel metal1 18492 14994 18492 14994 0 _121_
rlabel metal1 19044 14042 19044 14042 0 _122_
rlabel metal2 20102 15504 20102 15504 0 _123_
rlabel metal1 16560 16558 16560 16558 0 _124_
rlabel metal1 7222 25126 7222 25126 0 _125_
rlabel metal1 10902 19788 10902 19788 0 _126_
rlabel metal1 10718 20366 10718 20366 0 _127_
rlabel metal1 13064 20298 13064 20298 0 _128_
rlabel metal1 12972 19278 12972 19278 0 _129_
rlabel metal1 13708 16558 13708 16558 0 _130_
rlabel metal1 13570 19890 13570 19890 0 _131_
rlabel metal1 13570 17170 13570 17170 0 _132_
rlabel metal2 13754 16864 13754 16864 0 _133_
rlabel metal2 10442 15266 10442 15266 0 _134_
rlabel metal1 6256 21658 6256 21658 0 _135_
rlabel metal1 8004 15538 8004 15538 0 _136_
rlabel metal1 11362 15470 11362 15470 0 _137_
rlabel metal1 12926 15538 12926 15538 0 _138_
rlabel metal1 11592 15878 11592 15878 0 _139_
rlabel metal1 12328 15470 12328 15470 0 _140_
rlabel metal1 13892 16626 13892 16626 0 _141_
rlabel metal1 16054 16524 16054 16524 0 _142_
rlabel metal1 15870 16592 15870 16592 0 _143_
rlabel metal1 16790 16626 16790 16626 0 _144_
rlabel metal1 19918 16116 19918 16116 0 _145_
rlabel metal1 20654 16014 20654 16014 0 _146_
rlabel metal1 21206 17748 21206 17748 0 _147_
rlabel metal1 21804 16014 21804 16014 0 _148_
rlabel metal1 22678 16048 22678 16048 0 _149_
rlabel metal1 23276 17646 23276 17646 0 _150_
rlabel metal1 21022 16626 21022 16626 0 _151_
rlabel metal1 19504 16558 19504 16558 0 _152_
rlabel metal1 18630 17102 18630 17102 0 _153_
rlabel metal2 7682 24412 7682 24412 0 _154_
rlabel metal1 15502 25330 15502 25330 0 _155_
rlabel metal1 15732 24378 15732 24378 0 _156_
rlabel metal1 11224 20842 11224 20842 0 _157_
rlabel metal1 10212 20774 10212 20774 0 _158_
rlabel metal2 10074 21114 10074 21114 0 _159_
rlabel metal1 9982 21556 9982 21556 0 _160_
rlabel metal1 13386 21420 13386 21420 0 _161_
rlabel metal1 12926 21386 12926 21386 0 _162_
rlabel metal2 13570 21556 13570 21556 0 _163_
rlabel metal2 13110 21590 13110 21590 0 _164_
rlabel metal1 13800 21522 13800 21522 0 _165_
rlabel metal1 13984 19890 13984 19890 0 _166_
rlabel metal2 14214 21216 14214 21216 0 _167_
rlabel metal1 18170 17646 18170 17646 0 _168_
rlabel metal1 8602 17238 8602 17238 0 _169_
rlabel metal1 9338 17170 9338 17170 0 _170_
rlabel metal2 5382 21420 5382 21420 0 _171_
rlabel metal1 13156 16762 13156 16762 0 _172_
rlabel metal2 9062 16660 9062 16660 0 _173_
rlabel metal2 8878 16422 8878 16422 0 _174_
rlabel metal1 9706 17578 9706 17578 0 _175_
rlabel metal2 11454 17408 11454 17408 0 _176_
rlabel metal1 10810 17646 10810 17646 0 _177_
rlabel via1 12282 17510 12282 17510 0 _178_
rlabel metal1 12466 17578 12466 17578 0 _179_
rlabel metal1 12804 17238 12804 17238 0 _180_
rlabel metal1 13386 17136 13386 17136 0 _181_
rlabel metal1 13202 17238 13202 17238 0 _182_
rlabel metal1 15824 17102 15824 17102 0 _183_
rlabel metal1 18538 17782 18538 17782 0 _184_
rlabel metal1 18906 17714 18906 17714 0 _185_
rlabel metal1 18446 17102 18446 17102 0 _186_
rlabel metal1 19136 16626 19136 16626 0 _187_
rlabel metal1 20240 17646 20240 17646 0 _188_
rlabel metal1 20838 17238 20838 17238 0 _189_
rlabel metal1 20838 16524 20838 16524 0 _190_
rlabel metal1 22034 17204 22034 17204 0 _191_
rlabel metal1 21850 17136 21850 17136 0 _192_
rlabel metal2 22034 17510 22034 17510 0 _193_
rlabel metal1 23046 20910 23046 20910 0 _194_
rlabel metal1 20838 21522 20838 21522 0 _195_
rlabel metal2 20838 18292 20838 18292 0 _196_
rlabel metal1 19550 18734 19550 18734 0 _197_
rlabel metal1 15962 20434 15962 20434 0 _198_
rlabel metal1 10166 20434 10166 20434 0 _199_
rlabel metal1 10350 20536 10350 20536 0 _200_
rlabel metal1 10350 20944 10350 20944 0 _201_
rlabel metal1 11730 21454 11730 21454 0 _202_
rlabel metal1 12282 21481 12282 21481 0 _203_
rlabel metal1 13938 21556 13938 21556 0 _204_
rlabel metal1 15594 20434 15594 20434 0 _205_
rlabel metal1 17204 21590 17204 21590 0 _206_
rlabel metal1 18354 19346 18354 19346 0 _207_
rlabel metal1 17296 18258 17296 18258 0 _208_
rlabel metal1 10764 16422 10764 16422 0 _209_
rlabel metal1 10258 15674 10258 15674 0 _210_
rlabel metal1 10074 17646 10074 17646 0 _211_
rlabel metal1 10672 17714 10672 17714 0 _212_
rlabel metal2 10994 18054 10994 18054 0 _213_
rlabel metal1 10672 17850 10672 17850 0 _214_
rlabel metal1 12834 18224 12834 18224 0 _215_
rlabel metal1 16606 18190 16606 18190 0 _216_
rlabel metal1 18078 19380 18078 19380 0 _217_
rlabel metal1 18584 19346 18584 19346 0 _218_
rlabel metal1 19504 19346 19504 19346 0 _219_
rlabel metal1 19826 19380 19826 19380 0 _220_
rlabel metal1 19504 18802 19504 18802 0 _221_
rlabel metal1 20562 18836 20562 18836 0 _222_
rlabel metal2 20102 19380 20102 19380 0 _223_
rlabel metal1 21068 21522 21068 21522 0 _224_
rlabel metal1 21022 21930 21022 21930 0 _225_
rlabel metal1 22264 21522 22264 21522 0 _226_
rlabel metal1 22770 21318 22770 21318 0 _227_
rlabel metal1 23138 21998 23138 21998 0 _228_
rlabel metal2 13386 22848 13386 22848 0 _229_
rlabel metal1 12926 23086 12926 23086 0 _230_
rlabel metal1 20332 21930 20332 21930 0 _231_
rlabel metal1 19872 20434 19872 20434 0 _232_
rlabel metal1 15410 22644 15410 22644 0 _233_
rlabel metal2 15594 21318 15594 21318 0 _234_
rlabel metal1 16330 21522 16330 21522 0 _235_
rlabel metal1 10810 20842 10810 20842 0 _236_
rlabel metal1 10856 20910 10856 20910 0 _237_
rlabel metal1 10534 20944 10534 20944 0 _238_
rlabel metal1 13662 21556 13662 21556 0 _239_
rlabel metal2 14582 21522 14582 21522 0 _240_
rlabel metal1 15962 21454 15962 21454 0 _241_
rlabel metal2 17434 21760 17434 21760 0 _242_
rlabel metal1 16698 21454 16698 21454 0 _243_
rlabel metal1 18308 20910 18308 20910 0 _244_
rlabel metal1 18354 21114 18354 21114 0 _245_
rlabel metal1 14766 16762 14766 16762 0 _246_
rlabel metal2 15318 18292 15318 18292 0 _247_
rlabel metal1 9890 17578 9890 17578 0 _248_
rlabel metal1 10350 17680 10350 17680 0 _249_
rlabel metal2 12650 18428 12650 18428 0 _250_
rlabel metal1 15456 18598 15456 18598 0 _251_
rlabel metal1 14766 18734 14766 18734 0 _252_
rlabel metal1 17802 18632 17802 18632 0 _253_
rlabel metal1 17204 19278 17204 19278 0 _254_
rlabel metal2 17710 19652 17710 19652 0 _255_
rlabel metal1 17894 20366 17894 20366 0 _256_
rlabel metal2 19182 20638 19182 20638 0 _257_
rlabel metal1 18492 20366 18492 20366 0 _258_
rlabel metal1 19826 20774 19826 20774 0 _259_
rlabel metal1 19826 20944 19826 20944 0 _260_
rlabel metal1 20148 21114 20148 21114 0 _261_
rlabel metal1 20616 21862 20616 21862 0 _262_
rlabel metal1 21160 21590 21160 21590 0 _263_
rlabel metal1 21298 22032 21298 22032 0 _264_
rlabel metal1 21712 21658 21712 21658 0 _265_
rlabel metal1 23046 22066 23046 22066 0 _266_
rlabel metal1 23460 23698 23460 23698 0 _267_
rlabel metal1 21436 23630 21436 23630 0 _268_
rlabel metal1 15180 22610 15180 22610 0 _269_
rlabel metal1 15364 22202 15364 22202 0 _270_
rlabel metal1 16100 23018 16100 23018 0 _271_
rlabel metal1 16744 21658 16744 21658 0 _272_
rlabel metal1 17480 22610 17480 22610 0 _273_
rlabel metal1 15594 18292 15594 18292 0 _274_
rlabel metal1 15318 17714 15318 17714 0 _275_
rlabel metal1 16790 18734 16790 18734 0 _276_
rlabel metal1 17020 19210 17020 19210 0 _277_
rlabel metal1 17020 19346 17020 19346 0 _278_
rlabel metal1 17480 22542 17480 22542 0 _279_
rlabel metal2 18262 22202 18262 22202 0 _280_
rlabel metal1 18400 21998 18400 21998 0 _281_
rlabel metal1 18722 21998 18722 21998 0 _282_
rlabel metal1 19519 22610 19519 22610 0 _283_
rlabel metal1 19320 24786 19320 24786 0 _284_
rlabel metal1 20286 23290 20286 23290 0 _285_
rlabel metal1 12558 24106 12558 24106 0 _286_
rlabel metal1 12696 24922 12696 24922 0 _287_
rlabel metal1 13202 23766 13202 23766 0 _288_
rlabel metal1 13754 23630 13754 23630 0 _289_
rlabel metal1 12926 25874 12926 25874 0 _290_
rlabel metal1 13984 24650 13984 24650 0 _291_
rlabel metal1 13938 23834 13938 23834 0 _292_
rlabel metal1 17572 23698 17572 23698 0 _293_
rlabel metal1 21068 23562 21068 23562 0 _294_
rlabel metal1 21252 23222 21252 23222 0 _295_
rlabel metal1 21804 23290 21804 23290 0 _296_
rlabel metal1 22632 23698 22632 23698 0 _297_
rlabel metal1 23092 25262 23092 25262 0 _298_
rlabel metal1 20884 25126 20884 25126 0 _299_
rlabel metal1 15870 22746 15870 22746 0 _300_
rlabel metal1 16928 24174 16928 24174 0 _301_
rlabel metal1 16284 18394 16284 18394 0 _302_
rlabel metal1 16928 24242 16928 24242 0 _303_
rlabel metal1 17756 25194 17756 25194 0 _304_
rlabel metal1 18170 24208 18170 24208 0 _305_
rlabel metal1 18262 24174 18262 24174 0 _306_
rlabel metal1 18630 25432 18630 25432 0 _307_
rlabel metal1 18860 24718 18860 24718 0 _308_
rlabel metal1 18952 25330 18952 25330 0 _309_
rlabel metal1 20792 24786 20792 24786 0 _310_
rlabel metal1 13478 25806 13478 25806 0 _311_
rlabel metal1 11960 25262 11960 25262 0 _312_
rlabel metal2 11822 25670 11822 25670 0 _313_
rlabel metal1 13846 25908 13846 25908 0 _314_
rlabel metal1 10948 25466 10948 25466 0 _315_
rlabel metal1 11684 25942 11684 25942 0 _316_
rlabel metal1 13202 26452 13202 26452 0 _317_
rlabel metal1 12006 26418 12006 26418 0 _318_
rlabel metal1 12190 25874 12190 25874 0 _319_
rlabel metal1 12742 25806 12742 25806 0 _320_
rlabel metal1 13892 24718 13892 24718 0 _321_
rlabel metal1 14122 27370 14122 27370 0 _322_
rlabel metal1 14674 24718 14674 24718 0 _323_
rlabel metal1 19596 25194 19596 25194 0 _324_
rlabel metal1 21068 25262 21068 25262 0 _325_
rlabel metal1 20240 25262 20240 25262 0 _326_
rlabel metal2 20930 25024 20930 25024 0 _327_
rlabel metal1 22954 25364 22954 25364 0 _328_
rlabel metal2 23046 25534 23046 25534 0 _329_
rlabel metal1 17572 26214 17572 26214 0 _330_
rlabel metal1 12098 26894 12098 26894 0 _331_
rlabel metal2 13018 26214 13018 26214 0 _332_
rlabel metal1 12558 26894 12558 26894 0 _333_
rlabel metal1 13163 27030 13163 27030 0 _334_
rlabel metal1 13018 27336 13018 27336 0 _335_
rlabel metal2 12558 27268 12558 27268 0 _336_
rlabel metal1 12512 26554 12512 26554 0 _337_
rlabel metal1 14306 27472 14306 27472 0 _338_
rlabel metal1 14674 27404 14674 27404 0 _339_
rlabel metal1 14904 27098 14904 27098 0 _340_
rlabel metal1 17250 26384 17250 26384 0 _341_
rlabel metal2 18262 25466 18262 25466 0 _342_
rlabel metal1 20608 25262 20608 25262 0 _343_
rlabel metal1 19274 25874 19274 25874 0 _344_
rlabel metal1 20700 25874 20700 25874 0 _345_
rlabel metal1 21160 25466 21160 25466 0 _346_
rlabel metal1 21298 25806 21298 25806 0 _347_
rlabel metal1 22126 26962 22126 26962 0 _348_
rlabel metal2 16054 26690 16054 26690 0 _349_
rlabel metal1 15916 24718 15916 24718 0 _350_
rlabel metal1 15962 26316 15962 26316 0 _351_
rlabel metal1 15272 25874 15272 25874 0 _352_
rlabel metal1 14122 26010 14122 26010 0 _353_
rlabel metal1 14260 26962 14260 26962 0 _354_
rlabel metal1 13708 26962 13708 26962 0 _355_
rlabel metal1 15594 26996 15594 26996 0 _356_
rlabel metal1 15410 26894 15410 26894 0 _357_
rlabel metal1 16514 26282 16514 26282 0 _358_
rlabel metal1 17342 26894 17342 26894 0 _359_
rlabel metal1 16606 26350 16606 26350 0 _360_
rlabel metal1 17572 26282 17572 26282 0 _361_
rlabel metal1 17480 26826 17480 26826 0 _362_
rlabel metal1 17710 26350 17710 26350 0 _363_
rlabel metal1 19366 26758 19366 26758 0 _364_
rlabel metal1 21421 26962 21421 26962 0 _365_
rlabel metal1 21068 27030 21068 27030 0 _366_
rlabel metal2 19274 27268 19274 27268 0 _367_
rlabel metal1 21482 26894 21482 26894 0 _368_
rlabel metal1 15732 26010 15732 26010 0 _369_
rlabel metal1 15916 25466 15916 25466 0 _370_
rlabel metal1 17434 27030 17434 27030 0 _371_
rlabel metal1 18308 26962 18308 26962 0 _372_
rlabel metal1 17802 26758 17802 26758 0 _373_
rlabel metal1 18906 27506 18906 27506 0 _374_
rlabel metal1 17250 26554 17250 26554 0 _375_
rlabel metal2 19182 27200 19182 27200 0 _376_
rlabel metal1 21574 27472 21574 27472 0 _377_
rlabel metal1 23276 25806 23276 25806 0 _378_
rlabel metal1 23506 25942 23506 25942 0 _379_
rlabel metal1 12512 11186 12512 11186 0 _380_
rlabel metal1 20286 12240 20286 12240 0 _381_
rlabel metal1 15042 12206 15042 12206 0 _382_
rlabel metal1 12558 19754 12558 19754 0 _383_
rlabel metal1 12236 14382 12236 14382 0 _384_
rlabel metal1 10856 12410 10856 12410 0 _385_
rlabel metal1 9844 23698 9844 23698 0 _386_
rlabel metal1 7912 13294 7912 13294 0 _387_
rlabel metal1 9575 12886 9575 12886 0 _388_
rlabel metal1 8372 15470 8372 15470 0 _389_
rlabel metal1 8694 22066 8694 22066 0 _390_
rlabel metal1 7413 19346 7413 19346 0 _391_
rlabel metal1 9798 20366 9798 20366 0 _392_
rlabel via1 9522 19299 9522 19299 0 _393_
rlabel metal1 11730 12172 11730 12172 0 _394_
rlabel metal1 21988 12274 21988 12274 0 _395_
rlabel metal1 11960 12206 11960 12206 0 _396_
rlabel metal1 12190 11798 12190 11798 0 _397_
rlabel metal1 7406 14858 7406 14858 0 _398_
rlabel metal1 8740 15062 8740 15062 0 _399_
rlabel metal2 8694 15436 8694 15436 0 _400_
rlabel metal2 12006 13498 12006 13498 0 _401_
rlabel metal2 7314 20128 7314 20128 0 _402_
rlabel via2 14030 20757 14030 20757 0 _403_
rlabel metal1 15594 14960 15594 14960 0 _404_
rlabel metal1 12190 13260 12190 13260 0 _405_
rlabel metal1 10810 12716 10810 12716 0 _406_
rlabel metal1 15594 13872 15594 13872 0 _407_
rlabel metal1 11408 12206 11408 12206 0 _408_
rlabel metal1 11822 11730 11822 11730 0 _409_
rlabel metal1 22126 11662 22126 11662 0 _410_
rlabel metal1 7130 16150 7130 16150 0 _411_
rlabel metal1 8510 14416 8510 14416 0 _412_
rlabel metal3 820 4148 820 4148 0 a[0]
rlabel metal3 820 8500 820 8500 0 a[1]
rlabel metal3 820 12852 820 12852 0 a[2]
rlabel metal3 820 17204 820 17204 0 a[3]
rlabel metal3 820 21556 820 21556 0 a[4]
rlabel metal3 751 25908 751 25908 0 a[5]
rlabel metal3 1050 30260 1050 30260 0 a[6]
rlabel metal3 820 34612 820 34612 0 a[7]
rlabel metal3 820 6324 820 6324 0 b[0]
rlabel metal3 751 10676 751 10676 0 b[1]
rlabel metal3 751 15028 751 15028 0 b[2]
rlabel metal3 820 19380 820 19380 0 b[3]
rlabel metal3 820 23732 820 23732 0 b[4]
rlabel metal3 820 28084 820 28084 0 b[5]
rlabel metal3 820 32436 820 32436 0 b[6]
rlabel metal3 820 36788 820 36788 0 b[7]
rlabel metal2 9062 1027 9062 1027 0 clk
rlabel metal3 820 1972 820 1972 0 control
rlabel metal1 3128 4794 3128 4794 0 net1
rlabel metal1 3082 11186 3082 11186 0 net10
rlabel metal2 4370 15198 4370 15198 0 net11
rlabel metal2 4646 18156 4646 18156 0 net12
rlabel metal1 1610 24072 1610 24072 0 net13
rlabel metal2 1610 28016 1610 28016 0 net14
rlabel metal1 3174 32742 3174 32742 0 net15
rlabel metal1 3128 36006 3128 36006 0 net16
rlabel metal1 20654 3502 20654 3502 0 net17
rlabel metal1 3174 2618 3174 2618 0 net18
rlabel metal2 23230 2924 23230 2924 0 net19
rlabel metal1 3220 9146 3220 9146 0 net2
rlabel metal1 23046 3400 23046 3400 0 net20
rlabel metal2 33166 24650 33166 24650 0 net21
rlabel metal2 33258 26622 33258 26622 0 net22
rlabel metal2 33350 28016 33350 28016 0 net23
rlabel metal2 33166 29546 33166 29546 0 net24
rlabel metal1 28428 33966 28428 33966 0 net25
rlabel metal1 29394 36142 29394 36142 0 net26
rlabel metal1 23598 5576 23598 5576 0 net27
rlabel metal2 15226 10336 15226 10336 0 net28
rlabel metal1 25737 10506 25737 10506 0 net29
rlabel metal1 2185 13158 2185 13158 0 net3
rlabel metal1 25691 11526 25691 11526 0 net30
rlabel metal2 33166 14212 33166 14212 0 net31
rlabel metal2 33166 16388 33166 16388 0 net32
rlabel metal2 33166 18122 33166 18122 0 net33
rlabel metal1 33166 20842 33166 20842 0 net34
rlabel metal1 33166 22644 33166 22644 0 net35
rlabel metal1 1610 17544 1610 17544 0 net4
rlabel metal1 1610 21624 1610 21624 0 net5
rlabel metal1 1610 26248 1610 26248 0 net6
rlabel metal2 4830 28730 4830 28730 0 net7
rlabel metal1 2760 34918 2760 34918 0 net8
rlabel metal1 3266 6630 3266 6630 0 net9
rlabel metal3 35336 3060 35336 3060 0 p[0]
rlabel metal3 35060 24820 35060 24820 0 p[10]
rlabel metal3 35336 26996 35336 26996 0 p[11]
rlabel metal3 35336 29172 35336 29172 0 p[12]
rlabel metal3 35060 31348 35060 31348 0 p[13]
rlabel metal3 35336 33524 35336 33524 0 p[14]
rlabel metal3 35060 35700 35060 35700 0 p[15]
rlabel metal3 35060 5236 35060 5236 0 p[1]
rlabel metal3 35336 7412 35336 7412 0 p[2]
rlabel metal3 35060 9588 35060 9588 0 p[3]
rlabel metal3 35336 11764 35336 11764 0 p[4]
rlabel metal3 35336 13940 35336 13940 0 p[5]
rlabel metal1 34638 16490 34638 16490 0 p[6]
rlabel metal3 35336 18292 35336 18292 0 p[7]
rlabel metal3 35060 20468 35060 20468 0 p[8]
rlabel metal3 35336 22644 35336 22644 0 p[9]
rlabel metal2 27278 1027 27278 1027 0 rst
<< properties >>
string FIXED_BBOX 0 0 36400 38800
<< end >>
