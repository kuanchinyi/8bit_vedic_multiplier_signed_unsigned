magic
tech sky130A
magscale 1 2
timestamp 1726899429
<< obsli1 >>
rect 1104 2159 35236 36465
<< obsm1 >>
rect 934 2128 35406 36496
<< metal2 >>
rect 938 0 994 800
rect 1950 0 2006 800
rect 2962 0 3018 800
rect 3974 0 4030 800
rect 4986 0 5042 800
rect 5998 0 6054 800
rect 7010 0 7066 800
rect 8022 0 8078 800
rect 9034 0 9090 800
rect 10046 0 10102 800
rect 11058 0 11114 800
rect 12070 0 12126 800
rect 13082 0 13138 800
rect 14094 0 14150 800
rect 15106 0 15162 800
rect 16118 0 16174 800
rect 17130 0 17186 800
rect 18142 0 18198 800
rect 19154 0 19210 800
rect 20166 0 20222 800
rect 21178 0 21234 800
rect 22190 0 22246 800
rect 23202 0 23258 800
rect 24214 0 24270 800
rect 25226 0 25282 800
rect 26238 0 26294 800
rect 27250 0 27306 800
rect 28262 0 28318 800
rect 29274 0 29330 800
rect 30286 0 30342 800
rect 31298 0 31354 800
rect 32310 0 32366 800
rect 33322 0 33378 800
rect 34334 0 34390 800
rect 35346 0 35402 800
<< obsm2 >>
rect 940 856 35400 36485
rect 1050 734 1894 856
rect 2062 734 2906 856
rect 3074 734 3918 856
rect 4086 734 4930 856
rect 5098 734 5942 856
rect 6110 734 6954 856
rect 7122 734 7966 856
rect 8134 734 8978 856
rect 9146 734 9990 856
rect 10158 734 11002 856
rect 11170 734 12014 856
rect 12182 734 13026 856
rect 13194 734 14038 856
rect 14206 734 15050 856
rect 15218 734 16062 856
rect 16230 734 17074 856
rect 17242 734 18086 856
rect 18254 734 19098 856
rect 19266 734 20110 856
rect 20278 734 21122 856
rect 21290 734 22134 856
rect 22302 734 23146 856
rect 23314 734 24158 856
rect 24326 734 25170 856
rect 25338 734 26182 856
rect 26350 734 27194 856
rect 27362 734 28206 856
rect 28374 734 29218 856
rect 29386 734 30230 856
rect 30398 734 31242 856
rect 31410 734 32254 856
rect 32422 734 33266 856
rect 33434 734 34278 856
rect 34446 734 35290 856
<< obsm3 >>
rect 4210 2143 35246 36481
<< metal4 >>
rect 4208 2128 4528 36496
rect 19568 2128 19888 36496
rect 34928 2128 35248 36496
<< obsm4 >>
rect 14411 7787 14477 11117
<< labels >>
rlabel metal2 s 938 0 994 800 6 a[0]
port 1 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 a[1]
port 2 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 a[2]
port 3 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 a[3]
port 4 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 a[4]
port 5 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 a[5]
port 6 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 a[6]
port 7 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 a[7]
port 8 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 b[0]
port 9 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 b[1]
port 10 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 b[2]
port 11 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 b[3]
port 12 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 b[4]
port 13 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 b[5]
port 14 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 b[6]
port 15 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 b[7]
port 16 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 clk
port 17 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 control
port 18 nsew signal input
rlabel metal2 s 17130 0 17186 800 6 p[0]
port 19 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 p[10]
port 20 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 p[11]
port 21 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 p[12]
port 22 nsew signal output
rlabel metal2 s 30286 0 30342 800 6 p[13]
port 23 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 p[14]
port 24 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 p[15]
port 25 nsew signal output
rlabel metal2 s 18142 0 18198 800 6 p[1]
port 26 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 p[2]
port 27 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 p[3]
port 28 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 p[4]
port 29 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 p[5]
port 30 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 p[6]
port 31 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 p[7]
port 32 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 p[8]
port 33 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 p[9]
port 34 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 rst
port 35 nsew signal input
rlabel metal4 s 4208 2128 4528 36496 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 36496 6 vccd1
port 36 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 36496 6 vssd1
port 37 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 36400 38800
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1917120
string GDS_FILE /home/cykuan/chinyi2/8bit_vedic_multiplier_signed_unsigned/openlane/vmsu_8bit_top/runs/24_09_21_14_16/results/signoff/vmsu_8bit_top.magic.gds
string GDS_START 631526
<< end >>

