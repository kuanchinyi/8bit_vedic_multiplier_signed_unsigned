// This is the unpowered netlist.
module vmsu_8bit_top (clk,
    control,
    rst,
    a,
    b,
    p);
 input clk;
 input control;
 input rst;
 input [7:0] a;
 input [7:0] b;
 output [15:0] p;

 wire \FA0.q ;
 wire \FA1.q ;
 wire \FA2.q ;
 wire \FA3.q ;
 wire \FA4.q ;
 wire \FA5.q ;
 wire \FA6.q ;
 wire \FA7.q ;
 wire \FB0.q ;
 wire \FB1.q ;
 wire \FB2.q ;
 wire \FB3.q ;
 wire \FB4.q ;
 wire \FB5.q ;
 wire \FB6.q ;
 wire \FB7.q ;
 wire \FC.q ;
 wire \FP0.d ;
 wire \FP1.d ;
 wire \FP10.d ;
 wire \FP11.d ;
 wire \FP12.d ;
 wire \FP13.d ;
 wire \FP14.d ;
 wire \FP15.d ;
 wire \FP2.d ;
 wire \FP3.d ;
 wire \FP4.d ;
 wire \FP5.d ;
 wire \FP6.d ;
 wire \FP7.d ;
 wire \FP8.d ;
 wire \FP9.d ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__515__B (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__551__C (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__551__D_N (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__552__A2_N (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__552__B1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__586__B (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__588__A2 (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__588__B1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__590__A3 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__A2_N (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__624__B1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__625__A2 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__653__A2 (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__653__B1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__665__B (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__680__C1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__692__C (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__692__D_N (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__693__A2_N (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__693__B1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__708__B (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__710__C_N (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__727__B (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__728__B (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__729__A1 (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__748__A2 (.DIODE(_068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__748__C1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__753__B1 (.DIODE(_104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__808__D (.DIODE(net18));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_95 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__inv_2 _380_ (.A(\FA0.q ),
    .Y(_250_));
 sky130_fd_sc_hd__inv_2 _381_ (.A(\FB0.q ),
    .Y(_261_));
 sky130_fd_sc_hd__nand2_1 _382_ (.A(\FA0.q ),
    .B(\FB0.q ),
    .Y(_272_));
 sky130_fd_sc_hd__inv_2 _383_ (.A(_272_),
    .Y(\FP0.d ));
 sky130_fd_sc_hd__and2_4 _384_ (.A(\FC.q ),
    .B(\FB7.q ),
    .X(_293_));
 sky130_fd_sc_hd__and3_4 _385_ (.A(\FC.q ),
    .B(\FB7.q ),
    .C(\FB0.q ),
    .X(_304_));
 sky130_fd_sc_hd__xor2_4 _386_ (.A(\FB1.q ),
    .B(_304_),
    .X(_314_));
 sky130_fd_sc_hd__xnor2_4 _387_ (.A(\FB1.q ),
    .B(_304_),
    .Y(_318_));
 sky130_fd_sc_hd__and2_4 _388_ (.A(\FC.q ),
    .B(\FA7.q ),
    .X(_322_));
 sky130_fd_sc_hd__and3_2 _389_ (.A(\FC.q ),
    .B(\FA7.q ),
    .C(\FA0.q ),
    .X(_323_));
 sky130_fd_sc_hd__xor2_2 _390_ (.A(\FA1.q ),
    .B(_323_),
    .X(_324_));
 sky130_fd_sc_hd__xnor2_4 _391_ (.A(\FA1.q ),
    .B(_323_),
    .Y(_325_));
 sky130_fd_sc_hd__o22a_1 _392_ (.A1(_250_),
    .A2(_318_),
    .B1(_325_),
    .B2(_261_),
    .X(_326_));
 sky130_fd_sc_hd__xor2_4 _393_ (.A(_293_),
    .B(_322_),
    .X(_327_));
 sky130_fd_sc_hd__xnor2_4 _394_ (.A(_293_),
    .B(_322_),
    .Y(_328_));
 sky130_fd_sc_hd__a21o_1 _395_ (.A1(_272_),
    .A2(_326_),
    .B1(_328_),
    .X(_329_));
 sky130_fd_sc_hd__o211a_4 _396_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .B1(\FC.q ),
    .C1(\FB7.q ),
    .X(_330_));
 sky130_fd_sc_hd__xor2_4 _397_ (.A(\FB2.q ),
    .B(_330_),
    .X(_331_));
 sky130_fd_sc_hd__xnor2_4 _398_ (.A(\FB2.q ),
    .B(_330_),
    .Y(_332_));
 sky130_fd_sc_hd__nand2_1 _399_ (.A(\FA0.q ),
    .B(_331_),
    .Y(_333_));
 sky130_fd_sc_hd__o211a_2 _400_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .B1(\FC.q ),
    .C1(\FA7.q ),
    .X(_334_));
 sky130_fd_sc_hd__xor2_2 _401_ (.A(\FA2.q ),
    .B(_334_),
    .X(_335_));
 sky130_fd_sc_hd__xnor2_4 _402_ (.A(\FA2.q ),
    .B(_334_),
    .Y(_336_));
 sky130_fd_sc_hd__nand2_1 _403_ (.A(\FB0.q ),
    .B(_335_),
    .Y(_337_));
 sky130_fd_sc_hd__nand2_1 _404_ (.A(_333_),
    .B(_337_),
    .Y(_338_));
 sky130_fd_sc_hd__a2111o_1 _405_ (.A1(_333_),
    .A2(_337_),
    .B1(\FP0.d ),
    .C1(_318_),
    .D1(_325_),
    .X(_339_));
 sky130_fd_sc_hd__a31o_1 _406_ (.A1(_272_),
    .A2(_314_),
    .A3(_324_),
    .B1(_338_),
    .X(_340_));
 sky130_fd_sc_hd__nand2_1 _407_ (.A(_339_),
    .B(_340_),
    .Y(_341_));
 sky130_fd_sc_hd__o21a_1 _408_ (.A1(_328_),
    .A2(_341_),
    .B1(_329_),
    .X(_342_));
 sky130_fd_sc_hd__o311a_4 _409_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .A3(\FB2.q ),
    .B1(\FB7.q ),
    .C1(\FC.q ),
    .X(_343_));
 sky130_fd_sc_hd__xor2_4 _410_ (.A(\FB3.q ),
    .B(_343_),
    .X(_344_));
 sky130_fd_sc_hd__xnor2_4 _411_ (.A(\FB3.q ),
    .B(_343_),
    .Y(_345_));
 sky130_fd_sc_hd__or4_2 _412_ (.A(_250_),
    .B(_325_),
    .C(_332_),
    .D(_345_),
    .X(_346_));
 sky130_fd_sc_hd__a22o_1 _413_ (.A1(_324_),
    .A2(_331_),
    .B1(_344_),
    .B2(\FA0.q ),
    .X(_347_));
 sky130_fd_sc_hd__o311a_2 _414_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .A3(\FA2.q ),
    .B1(\FA7.q ),
    .C1(\FC.q ),
    .X(_348_));
 sky130_fd_sc_hd__xor2_2 _415_ (.A(\FA3.q ),
    .B(_348_),
    .X(_349_));
 sky130_fd_sc_hd__xnor2_4 _416_ (.A(\FA3.q ),
    .B(_348_),
    .Y(_350_));
 sky130_fd_sc_hd__or4_2 _417_ (.A(_261_),
    .B(_318_),
    .C(_336_),
    .D(_350_),
    .X(_351_));
 sky130_fd_sc_hd__a22o_1 _418_ (.A1(_314_),
    .A2(_335_),
    .B1(_349_),
    .B2(\FB0.q ),
    .X(_352_));
 sky130_fd_sc_hd__nand4_2 _419_ (.A(_346_),
    .B(_347_),
    .C(_351_),
    .D(_352_),
    .Y(_353_));
 sky130_fd_sc_hd__a22o_1 _420_ (.A1(_346_),
    .A2(_347_),
    .B1(_351_),
    .B2(_352_),
    .X(_354_));
 sky130_fd_sc_hd__nor2_1 _421_ (.A(_333_),
    .B(_337_),
    .Y(_355_));
 sky130_fd_sc_hd__and3_1 _422_ (.A(_353_),
    .B(_354_),
    .C(_355_),
    .X(_356_));
 sky130_fd_sc_hd__a21o_1 _423_ (.A1(_353_),
    .A2(_354_),
    .B1(_355_),
    .X(_357_));
 sky130_fd_sc_hd__and2b_1 _424_ (.A_N(_356_),
    .B(_357_),
    .X(_358_));
 sky130_fd_sc_hd__and4_1 _425_ (.A(\FA0.q ),
    .B(\FB0.q ),
    .C(_314_),
    .D(_324_),
    .X(_359_));
 sky130_fd_sc_hd__inv_2 _426_ (.A(_359_),
    .Y(_360_));
 sky130_fd_sc_hd__nand2_1 _427_ (.A(_339_),
    .B(_360_),
    .Y(_361_));
 sky130_fd_sc_hd__and3b_1 _428_ (.A_N(_356_),
    .B(_357_),
    .C(_361_),
    .X(_362_));
 sky130_fd_sc_hd__nor2_1 _429_ (.A(_358_),
    .B(_361_),
    .Y(_363_));
 sky130_fd_sc_hd__nor2_1 _430_ (.A(_362_),
    .B(_363_),
    .Y(_364_));
 sky130_fd_sc_hd__a21bo_1 _431_ (.A1(_327_),
    .A2(_364_),
    .B1_N(_342_),
    .X(_365_));
 sky130_fd_sc_hd__or4_4 _432_ (.A(\FB0.q ),
    .B(\FB1.q ),
    .C(\FB2.q ),
    .D(\FB3.q ),
    .X(_366_));
 sky130_fd_sc_hd__nand2_2 _433_ (.A(_293_),
    .B(_366_),
    .Y(_367_));
 sky130_fd_sc_hd__xor2_4 _434_ (.A(\FB4.q ),
    .B(_367_),
    .X(_368_));
 sky130_fd_sc_hd__inv_2 _435_ (.A(_368_),
    .Y(_369_));
 sky130_fd_sc_hd__nor2_1 _436_ (.A(_250_),
    .B(_368_),
    .Y(_370_));
 sky130_fd_sc_hd__or4_4 _437_ (.A(\FA0.q ),
    .B(\FA1.q ),
    .C(\FA2.q ),
    .D(\FA3.q ),
    .X(_371_));
 sky130_fd_sc_hd__nand2_2 _438_ (.A(_322_),
    .B(_371_),
    .Y(_372_));
 sky130_fd_sc_hd__xor2_4 _439_ (.A(\FA4.q ),
    .B(_372_),
    .X(_373_));
 sky130_fd_sc_hd__nor2_1 _440_ (.A(_261_),
    .B(_373_),
    .Y(_374_));
 sky130_fd_sc_hd__nand2_2 _441_ (.A(_370_),
    .B(_374_),
    .Y(_375_));
 sky130_fd_sc_hd__or2_1 _442_ (.A(_370_),
    .B(_374_),
    .X(_376_));
 sky130_fd_sc_hd__nand2_1 _443_ (.A(_375_),
    .B(_376_),
    .Y(_377_));
 sky130_fd_sc_hd__nor2_1 _444_ (.A(_332_),
    .B(_336_),
    .Y(_378_));
 sky130_fd_sc_hd__or3b_2 _445_ (.A(_325_),
    .B(_345_),
    .C_N(_333_),
    .X(_379_));
 sky130_fd_sc_hd__or3b_2 _446_ (.A(_318_),
    .B(_350_),
    .C_N(_337_),
    .X(_000_));
 sky130_fd_sc_hd__and2_1 _447_ (.A(_379_),
    .B(_000_),
    .X(_001_));
 sky130_fd_sc_hd__xor2_2 _448_ (.A(_379_),
    .B(_000_),
    .X(_002_));
 sky130_fd_sc_hd__a21boi_1 _449_ (.A1(_354_),
    .A2(_355_),
    .B1_N(_353_),
    .Y(_003_));
 sky130_fd_sc_hd__xnor2_2 _450_ (.A(_002_),
    .B(_003_),
    .Y(_004_));
 sky130_fd_sc_hd__xor2_1 _451_ (.A(_362_),
    .B(_004_),
    .X(_005_));
 sky130_fd_sc_hd__and2_1 _452_ (.A(_378_),
    .B(_005_),
    .X(_006_));
 sky130_fd_sc_hd__nor2_1 _453_ (.A(_378_),
    .B(_005_),
    .Y(_007_));
 sky130_fd_sc_hd__or2_1 _454_ (.A(_006_),
    .B(_007_),
    .X(_008_));
 sky130_fd_sc_hd__nor2_1 _455_ (.A(_377_),
    .B(_008_),
    .Y(_009_));
 sky130_fd_sc_hd__and2_1 _456_ (.A(_377_),
    .B(_008_),
    .X(_010_));
 sky130_fd_sc_hd__nor2_1 _457_ (.A(_009_),
    .B(_010_),
    .Y(_011_));
 sky130_fd_sc_hd__a21oi_1 _458_ (.A1(_327_),
    .A2(_011_),
    .B1(_365_),
    .Y(_012_));
 sky130_fd_sc_hd__or4_1 _459_ (.A(_332_),
    .B(_336_),
    .C(_345_),
    .D(_350_),
    .X(_013_));
 sky130_fd_sc_hd__a22o_1 _460_ (.A1(_335_),
    .A2(_344_),
    .B1(_349_),
    .B2(_331_),
    .X(_014_));
 sky130_fd_sc_hd__nand2_1 _461_ (.A(_013_),
    .B(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__xnor2_1 _462_ (.A(_346_),
    .B(_351_),
    .Y(_016_));
 sky130_fd_sc_hd__o21a_1 _463_ (.A1(_379_),
    .A2(_000_),
    .B1(_353_),
    .X(_017_));
 sky130_fd_sc_hd__o21ai_2 _464_ (.A1(_001_),
    .A2(_017_),
    .B1(_016_),
    .Y(_018_));
 sky130_fd_sc_hd__nand3_1 _465_ (.A(_362_),
    .B(_004_),
    .C(_018_),
    .Y(_019_));
 sky130_fd_sc_hd__a21o_1 _466_ (.A1(_362_),
    .A2(_004_),
    .B1(_018_),
    .X(_020_));
 sky130_fd_sc_hd__nand3b_2 _467_ (.A_N(_015_),
    .B(_019_),
    .C(_020_),
    .Y(_021_));
 sky130_fd_sc_hd__a21bo_1 _468_ (.A1(_019_),
    .A2(_020_),
    .B1_N(_015_),
    .X(_022_));
 sky130_fd_sc_hd__nand2_1 _469_ (.A(_021_),
    .B(_022_),
    .Y(_023_));
 sky130_fd_sc_hd__nand3_1 _470_ (.A(_006_),
    .B(_021_),
    .C(_022_),
    .Y(_024_));
 sky130_fd_sc_hd__a21o_1 _471_ (.A1(_021_),
    .A2(_022_),
    .B1(_006_),
    .X(_025_));
 sky130_fd_sc_hd__o21ai_4 _472_ (.A1(\FB4.q ),
    .A2(_366_),
    .B1(_293_),
    .Y(_026_));
 sky130_fd_sc_hd__xnor2_1 _473_ (.A(\FB5.q ),
    .B(_026_),
    .Y(_027_));
 sky130_fd_sc_hd__xor2_4 _474_ (.A(\FB5.q ),
    .B(_026_),
    .X(_028_));
 sky130_fd_sc_hd__or4_1 _475_ (.A(_250_),
    .B(_325_),
    .C(_368_),
    .D(_028_),
    .X(_029_));
 sky130_fd_sc_hd__a2bb2o_1 _476_ (.A1_N(_325_),
    .A2_N(_368_),
    .B1(_027_),
    .B2(\FA0.q ),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _477_ (.A(_029_),
    .B(_030_),
    .X(_031_));
 sky130_fd_sc_hd__o21ai_4 _478_ (.A1(\FA4.q ),
    .A2(_371_),
    .B1(_322_),
    .Y(_032_));
 sky130_fd_sc_hd__xnor2_1 _479_ (.A(\FA5.q ),
    .B(_032_),
    .Y(_033_));
 sky130_fd_sc_hd__xor2_4 _480_ (.A(\FA5.q ),
    .B(_032_),
    .X(_034_));
 sky130_fd_sc_hd__or4_1 _481_ (.A(_261_),
    .B(_318_),
    .C(_373_),
    .D(_034_),
    .X(_035_));
 sky130_fd_sc_hd__a2bb2o_1 _482_ (.A1_N(_318_),
    .A2_N(_373_),
    .B1(_033_),
    .B2(\FB0.q ),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _483_ (.A(_035_),
    .B(_036_),
    .X(_037_));
 sky130_fd_sc_hd__nand2_1 _484_ (.A(_031_),
    .B(_037_),
    .Y(_038_));
 sky130_fd_sc_hd__nor2_1 _485_ (.A(_031_),
    .B(_037_),
    .Y(_039_));
 sky130_fd_sc_hd__inv_2 _486_ (.A(_039_),
    .Y(_040_));
 sky130_fd_sc_hd__nand2_1 _487_ (.A(_038_),
    .B(_040_),
    .Y(_041_));
 sky130_fd_sc_hd__xnor2_1 _488_ (.A(_375_),
    .B(_041_),
    .Y(_042_));
 sky130_fd_sc_hd__xor2_1 _489_ (.A(_375_),
    .B(_041_),
    .X(_043_));
 sky130_fd_sc_hd__a21o_1 _490_ (.A1(_024_),
    .A2(_025_),
    .B1(_043_),
    .X(_044_));
 sky130_fd_sc_hd__nand3_1 _491_ (.A(_024_),
    .B(_025_),
    .C(_043_),
    .Y(_045_));
 sky130_fd_sc_hd__nand2_1 _492_ (.A(_044_),
    .B(_045_),
    .Y(_046_));
 sky130_fd_sc_hd__xor2_1 _493_ (.A(_009_),
    .B(_046_),
    .X(_047_));
 sky130_fd_sc_hd__o21ai_1 _494_ (.A1(_328_),
    .A2(_047_),
    .B1(_012_),
    .Y(_048_));
 sky130_fd_sc_hd__a2111o_1 _495_ (.A1(_023_),
    .A2(_042_),
    .B1(_377_),
    .C1(_006_),
    .D1(_007_),
    .X(_049_));
 sky130_fd_sc_hd__nand2_1 _496_ (.A(_045_),
    .B(_049_),
    .Y(_050_));
 sky130_fd_sc_hd__nand3_1 _497_ (.A(_358_),
    .B(_359_),
    .C(_018_),
    .Y(_051_));
 sky130_fd_sc_hd__a211oi_1 _498_ (.A1(_339_),
    .A2(_378_),
    .B1(_350_),
    .C1(_345_),
    .Y(_052_));
 sky130_fd_sc_hd__o2bb2a_1 _499_ (.A1_N(_051_),
    .A2_N(_052_),
    .B1(_346_),
    .B2(_351_),
    .X(_053_));
 sky130_fd_sc_hd__a21bo_1 _500_ (.A1(_006_),
    .A2(_022_),
    .B1_N(_021_),
    .X(_054_));
 sky130_fd_sc_hd__xor2_1 _501_ (.A(_053_),
    .B(_054_),
    .X(_055_));
 sky130_fd_sc_hd__a21oi_1 _502_ (.A1(_375_),
    .A2(_038_),
    .B1(_039_),
    .Y(_056_));
 sky130_fd_sc_hd__o31a_2 _503_ (.A1(\FB5.q ),
    .A2(\FB4.q ),
    .A3(_366_),
    .B1(_293_),
    .X(_057_));
 sky130_fd_sc_hd__xnor2_4 _504_ (.A(\FB6.q ),
    .B(_057_),
    .Y(_058_));
 sky130_fd_sc_hd__or2_2 _505_ (.A(_250_),
    .B(_058_),
    .X(_059_));
 sky130_fd_sc_hd__or2_1 _506_ (.A(_336_),
    .B(_368_),
    .X(_060_));
 sky130_fd_sc_hd__o311a_1 _507_ (.A1(_325_),
    .A2(_370_),
    .A3(_028_),
    .B1(_059_),
    .C1(_060_),
    .X(_061_));
 sky130_fd_sc_hd__nor2_2 _508_ (.A(_059_),
    .B(_060_),
    .Y(_062_));
 sky130_fd_sc_hd__a2111o_1 _509_ (.A1(_059_),
    .A2(_060_),
    .B1(_325_),
    .C1(_370_),
    .D1(_028_),
    .X(_063_));
 sky130_fd_sc_hd__and2b_1 _510_ (.A_N(_061_),
    .B(_063_),
    .X(_064_));
 sky130_fd_sc_hd__inv_2 _511_ (.A(_064_),
    .Y(_065_));
 sky130_fd_sc_hd__or2_2 _512_ (.A(_332_),
    .B(_373_),
    .X(_066_));
 sky130_fd_sc_hd__o31a_2 _513_ (.A1(\FA5.q ),
    .A2(\FA4.q ),
    .A3(_371_),
    .B1(_322_),
    .X(_067_));
 sky130_fd_sc_hd__xnor2_4 _514_ (.A(\FA6.q ),
    .B(_067_),
    .Y(_068_));
 sky130_fd_sc_hd__or2_1 _515_ (.A(_261_),
    .B(_068_),
    .X(_069_));
 sky130_fd_sc_hd__o311a_1 _516_ (.A1(_318_),
    .A2(_374_),
    .A3(_034_),
    .B1(_066_),
    .C1(_069_),
    .X(_070_));
 sky130_fd_sc_hd__nor2_1 _517_ (.A(_066_),
    .B(_069_),
    .Y(_071_));
 sky130_fd_sc_hd__a2111o_1 _518_ (.A1(_066_),
    .A2(_069_),
    .B1(_318_),
    .C1(_374_),
    .D1(_034_),
    .X(_072_));
 sky130_fd_sc_hd__or3b_1 _519_ (.A(_070_),
    .B(_071_),
    .C_N(_072_),
    .X(_073_));
 sky130_fd_sc_hd__nor3_1 _520_ (.A(_062_),
    .B(_065_),
    .C(_073_),
    .Y(_074_));
 sky130_fd_sc_hd__o21ai_1 _521_ (.A1(_062_),
    .A2(_065_),
    .B1(_073_),
    .Y(_075_));
 sky130_fd_sc_hd__and2b_1 _522_ (.A_N(_074_),
    .B(_075_),
    .X(_076_));
 sky130_fd_sc_hd__xnor2_1 _523_ (.A(_056_),
    .B(_076_),
    .Y(_077_));
 sky130_fd_sc_hd__nand2_1 _524_ (.A(_055_),
    .B(_077_),
    .Y(_078_));
 sky130_fd_sc_hd__or2_1 _525_ (.A(_055_),
    .B(_077_),
    .X(_079_));
 sky130_fd_sc_hd__and2_1 _526_ (.A(_078_),
    .B(_079_),
    .X(_080_));
 sky130_fd_sc_hd__xnor2_1 _527_ (.A(_050_),
    .B(_080_),
    .Y(_081_));
 sky130_fd_sc_hd__o21ba_1 _528_ (.A1(_328_),
    .A2(_081_),
    .B1_N(_048_),
    .X(_082_));
 sky130_fd_sc_hd__a22o_1 _529_ (.A1(_045_),
    .A2(_049_),
    .B1(_055_),
    .B2(_077_),
    .X(_083_));
 sky130_fd_sc_hd__or2_1 _530_ (.A(_021_),
    .B(_053_),
    .X(_084_));
 sky130_fd_sc_hd__o21a_1 _531_ (.A1(_056_),
    .A2(_074_),
    .B1(_075_),
    .X(_085_));
 sky130_fd_sc_hd__or4_1 _532_ (.A(\FB5.q ),
    .B(\FB4.q ),
    .C(\FB6.q ),
    .D(_366_),
    .X(_086_));
 sky130_fd_sc_hd__a21boi_4 _533_ (.A1(\FC.q ),
    .A2(_086_),
    .B1_N(\FB7.q ),
    .Y(_087_));
 sky130_fd_sc_hd__inv_2 _534_ (.A(_087_),
    .Y(_088_));
 sky130_fd_sc_hd__or4b_4 _535_ (.A(_250_),
    .B(_325_),
    .C(_058_),
    .D_N(_087_),
    .X(_089_));
 sky130_fd_sc_hd__a2bb2o_1 _536_ (.A1_N(_325_),
    .A2_N(_058_),
    .B1(_087_),
    .B2(\FA0.q ),
    .X(_090_));
 sky130_fd_sc_hd__or4_2 _537_ (.A(_336_),
    .B(_350_),
    .C(_368_),
    .D(_028_),
    .X(_091_));
 sky130_fd_sc_hd__a2bb2o_1 _538_ (.A1_N(_350_),
    .A2_N(_368_),
    .B1(_027_),
    .B2(_335_),
    .X(_092_));
 sky130_fd_sc_hd__nand4_1 _539_ (.A(_089_),
    .B(_090_),
    .C(_091_),
    .D(_092_),
    .Y(_093_));
 sky130_fd_sc_hd__a22o_1 _540_ (.A1(_089_),
    .A2(_090_),
    .B1(_091_),
    .B2(_092_),
    .X(_094_));
 sky130_fd_sc_hd__and3_1 _541_ (.A(_062_),
    .B(_093_),
    .C(_094_),
    .X(_095_));
 sky130_fd_sc_hd__a21oi_1 _542_ (.A1(_093_),
    .A2(_094_),
    .B1(_062_),
    .Y(_096_));
 sky130_fd_sc_hd__nor2_1 _543_ (.A(_095_),
    .B(_096_),
    .Y(_097_));
 sky130_fd_sc_hd__nand2_2 _544_ (.A(_029_),
    .B(_063_),
    .Y(_098_));
 sky130_fd_sc_hd__or3b_1 _545_ (.A(_095_),
    .B(_096_),
    .C_N(_098_),
    .X(_099_));
 sky130_fd_sc_hd__xnor2_2 _546_ (.A(_097_),
    .B(_098_),
    .Y(_100_));
 sky130_fd_sc_hd__or4_4 _547_ (.A(_332_),
    .B(_345_),
    .C(_373_),
    .D(_034_),
    .X(_101_));
 sky130_fd_sc_hd__a2bb2o_1 _548_ (.A1_N(_345_),
    .A2_N(_373_),
    .B1(_033_),
    .B2(_331_),
    .X(_102_));
 sky130_fd_sc_hd__or4_1 _549_ (.A(\FA5.q ),
    .B(\FA4.q ),
    .C(\FA6.q ),
    .D(_371_),
    .X(_103_));
 sky130_fd_sc_hd__a21boi_4 _550_ (.A1(\FC.q ),
    .A2(_103_),
    .B1_N(\FA7.q ),
    .Y(_104_));
 sky130_fd_sc_hd__or4b_4 _551_ (.A(_261_),
    .B(_318_),
    .C(_068_),
    .D_N(_104_),
    .X(_105_));
 sky130_fd_sc_hd__a2bb2o_1 _552_ (.A1_N(_318_),
    .A2_N(_068_),
    .B1(_104_),
    .B2(\FB0.q ),
    .X(_106_));
 sky130_fd_sc_hd__and4_1 _553_ (.A(_101_),
    .B(_102_),
    .C(_105_),
    .D(_106_),
    .X(_107_));
 sky130_fd_sc_hd__nand4_1 _554_ (.A(_101_),
    .B(_102_),
    .C(_105_),
    .D(_106_),
    .Y(_108_));
 sky130_fd_sc_hd__a22o_1 _555_ (.A1(_101_),
    .A2(_102_),
    .B1(_105_),
    .B2(_106_),
    .X(_109_));
 sky130_fd_sc_hd__nand3_1 _556_ (.A(_071_),
    .B(_108_),
    .C(_109_),
    .Y(_110_));
 sky130_fd_sc_hd__a21o_1 _557_ (.A1(_108_),
    .A2(_109_),
    .B1(_071_),
    .X(_111_));
 sky130_fd_sc_hd__nand2_1 _558_ (.A(_035_),
    .B(_072_),
    .Y(_112_));
 sky130_fd_sc_hd__and3_2 _559_ (.A(_110_),
    .B(_111_),
    .C(_112_),
    .X(_113_));
 sky130_fd_sc_hd__a21oi_1 _560_ (.A1(_110_),
    .A2(_111_),
    .B1(_112_),
    .Y(_114_));
 sky130_fd_sc_hd__or2_1 _561_ (.A(_113_),
    .B(_114_),
    .X(_115_));
 sky130_fd_sc_hd__nor2_1 _562_ (.A(_100_),
    .B(_115_),
    .Y(_116_));
 sky130_fd_sc_hd__nand2_1 _563_ (.A(_100_),
    .B(_115_),
    .Y(_117_));
 sky130_fd_sc_hd__xor2_1 _564_ (.A(_100_),
    .B(_115_),
    .X(_118_));
 sky130_fd_sc_hd__xnor2_1 _565_ (.A(_085_),
    .B(_118_),
    .Y(_119_));
 sky130_fd_sc_hd__a31o_1 _566_ (.A1(_013_),
    .A2(_051_),
    .A3(_084_),
    .B1(_119_),
    .X(_120_));
 sky130_fd_sc_hd__inv_2 _567_ (.A(_120_),
    .Y(_121_));
 sky130_fd_sc_hd__and4_1 _568_ (.A(_013_),
    .B(_051_),
    .C(_084_),
    .D(_119_),
    .X(_122_));
 sky130_fd_sc_hd__a211o_1 _569_ (.A1(_079_),
    .A2(_083_),
    .B1(_121_),
    .C1(_122_),
    .X(_123_));
 sky130_fd_sc_hd__o211ai_1 _570_ (.A1(_121_),
    .A2(_122_),
    .B1(_079_),
    .C1(_083_),
    .Y(_124_));
 sky130_fd_sc_hd__nand2_1 _571_ (.A(_123_),
    .B(_124_),
    .Y(_125_));
 sky130_fd_sc_hd__o21a_1 _572_ (.A1(_328_),
    .A2(_125_),
    .B1(_082_),
    .X(_126_));
 sky130_fd_sc_hd__or2_1 _573_ (.A(_368_),
    .B(_373_),
    .X(_127_));
 sky130_fd_sc_hd__a31o_1 _574_ (.A1(_079_),
    .A2(_083_),
    .A3(_120_),
    .B1(_122_),
    .X(_128_));
 sky130_fd_sc_hd__o21ai_2 _575_ (.A1(_085_),
    .A2(_116_),
    .B1(_117_),
    .Y(_129_));
 sky130_fd_sc_hd__nor2_1 _576_ (.A(_336_),
    .B(_058_),
    .Y(_130_));
 sky130_fd_sc_hd__o211a_1 _577_ (.A1(_336_),
    .A2(_368_),
    .B1(_027_),
    .C1(_349_),
    .X(_131_));
 sky130_fd_sc_hd__and4_1 _578_ (.A(_324_),
    .B(_059_),
    .C(_087_),
    .D(_131_),
    .X(_132_));
 sky130_fd_sc_hd__a31o_1 _579_ (.A1(_324_),
    .A2(_059_),
    .A3(_087_),
    .B1(_131_),
    .X(_133_));
 sky130_fd_sc_hd__and2b_1 _580_ (.A_N(_132_),
    .B(_133_),
    .X(_134_));
 sky130_fd_sc_hd__a21bo_1 _581_ (.A1(_062_),
    .A2(_094_),
    .B1_N(_093_),
    .X(_135_));
 sky130_fd_sc_hd__xor2_2 _582_ (.A(_134_),
    .B(_135_),
    .X(_136_));
 sky130_fd_sc_hd__xnor2_1 _583_ (.A(_099_),
    .B(_136_),
    .Y(_137_));
 sky130_fd_sc_hd__and2_1 _584_ (.A(_130_),
    .B(_137_),
    .X(_138_));
 sky130_fd_sc_hd__xnor2_1 _585_ (.A(_130_),
    .B(_137_),
    .Y(_139_));
 sky130_fd_sc_hd__nor2_2 _586_ (.A(_332_),
    .B(_068_),
    .Y(_140_));
 sky130_fd_sc_hd__nor2_1 _587_ (.A(_345_),
    .B(_034_),
    .Y(_141_));
 sky130_fd_sc_hd__o211a_1 _588_ (.A1(_261_),
    .A2(_068_),
    .B1(_104_),
    .C1(_314_),
    .X(_142_));
 sky130_fd_sc_hd__and3_1 _589_ (.A(_066_),
    .B(_141_),
    .C(_142_),
    .X(_143_));
 sky130_fd_sc_hd__a32oi_2 _590_ (.A1(_314_),
    .A2(_069_),
    .A3(_104_),
    .B1(_141_),
    .B2(_066_),
    .Y(_144_));
 sky130_fd_sc_hd__nor2_1 _591_ (.A(_143_),
    .B(_144_),
    .Y(_145_));
 sky130_fd_sc_hd__a21oi_1 _592_ (.A1(_071_),
    .A2(_109_),
    .B1(_107_),
    .Y(_146_));
 sky130_fd_sc_hd__xnor2_2 _593_ (.A(_145_),
    .B(_146_),
    .Y(_147_));
 sky130_fd_sc_hd__xor2_2 _594_ (.A(_113_),
    .B(_147_),
    .X(_148_));
 sky130_fd_sc_hd__and2_1 _595_ (.A(_140_),
    .B(_148_),
    .X(_149_));
 sky130_fd_sc_hd__xnor2_2 _596_ (.A(_140_),
    .B(_148_),
    .Y(_150_));
 sky130_fd_sc_hd__or2_1 _597_ (.A(_139_),
    .B(_150_),
    .X(_151_));
 sky130_fd_sc_hd__and2_1 _598_ (.A(_139_),
    .B(_150_),
    .X(_152_));
 sky130_fd_sc_hd__xnor2_1 _599_ (.A(_139_),
    .B(_150_),
    .Y(_153_));
 sky130_fd_sc_hd__xnor2_2 _600_ (.A(_129_),
    .B(_153_),
    .Y(_154_));
 sky130_fd_sc_hd__a311o_1 _601_ (.A1(_079_),
    .A2(_083_),
    .A3(_120_),
    .B1(_122_),
    .C1(_154_),
    .X(_155_));
 sky130_fd_sc_hd__xnor2_1 _602_ (.A(_128_),
    .B(_154_),
    .Y(_156_));
 sky130_fd_sc_hd__nor2_1 _603_ (.A(_127_),
    .B(_156_),
    .Y(_157_));
 sky130_fd_sc_hd__and2_1 _604_ (.A(_127_),
    .B(_156_),
    .X(_158_));
 sky130_fd_sc_hd__or2_1 _605_ (.A(_157_),
    .B(_158_),
    .X(_159_));
 sky130_fd_sc_hd__o21ai_1 _606_ (.A1(_328_),
    .A2(_159_),
    .B1(_126_),
    .Y(_160_));
 sky130_fd_sc_hd__and4bb_1 _607_ (.A_N(_368_),
    .B_N(_373_),
    .C(_027_),
    .D(_033_),
    .X(_161_));
 sky130_fd_sc_hd__o22a_1 _608_ (.A1(_373_),
    .A2(_028_),
    .B1(_034_),
    .B2(_368_),
    .X(_162_));
 sky130_fd_sc_hd__nor2_1 _609_ (.A(_161_),
    .B(_162_),
    .Y(_163_));
 sky130_fd_sc_hd__a21o_1 _610_ (.A1(_129_),
    .A2(_151_),
    .B1(_152_),
    .X(_164_));
 sky130_fd_sc_hd__or4_1 _611_ (.A(_336_),
    .B(_350_),
    .C(_058_),
    .D(_088_),
    .X(_165_));
 sky130_fd_sc_hd__a2bb2o_1 _612_ (.A1_N(_350_),
    .A2_N(_058_),
    .B1(_087_),
    .B2(_335_),
    .X(_166_));
 sky130_fd_sc_hd__and2_1 _613_ (.A(_165_),
    .B(_166_),
    .X(_167_));
 sky130_fd_sc_hd__or2_1 _614_ (.A(_089_),
    .B(_091_),
    .X(_168_));
 sky130_fd_sc_hd__nand2_1 _615_ (.A(_089_),
    .B(_091_),
    .Y(_169_));
 sky130_fd_sc_hd__a41o_1 _616_ (.A1(_089_),
    .A2(_090_),
    .A3(_091_),
    .A4(_092_),
    .B1(_132_),
    .X(_170_));
 sky130_fd_sc_hd__a22o_1 _617_ (.A1(_168_),
    .A2(_169_),
    .B1(_170_),
    .B2(_133_),
    .X(_171_));
 sky130_fd_sc_hd__nand3b_1 _618_ (.A_N(_099_),
    .B(_136_),
    .C(_171_),
    .Y(_172_));
 sky130_fd_sc_hd__a31o_1 _619_ (.A1(_097_),
    .A2(_098_),
    .A3(_136_),
    .B1(_171_),
    .X(_173_));
 sky130_fd_sc_hd__nand3_1 _620_ (.A(_167_),
    .B(_172_),
    .C(_173_),
    .Y(_174_));
 sky130_fd_sc_hd__a21o_1 _621_ (.A1(_172_),
    .A2(_173_),
    .B1(_167_),
    .X(_175_));
 sky130_fd_sc_hd__and3_1 _622_ (.A(_138_),
    .B(_174_),
    .C(_175_),
    .X(_176_));
 sky130_fd_sc_hd__a21oi_1 _623_ (.A1(_174_),
    .A2(_175_),
    .B1(_138_),
    .Y(_177_));
 sky130_fd_sc_hd__a2bb2oi_1 _624_ (.A1_N(_345_),
    .A2_N(_068_),
    .B1(_104_),
    .B2(_331_),
    .Y(_178_));
 sky130_fd_sc_hd__a31oi_2 _625_ (.A1(_344_),
    .A2(_104_),
    .A3(_140_),
    .B1(_178_),
    .Y(_179_));
 sky130_fd_sc_hd__xnor2_1 _626_ (.A(_101_),
    .B(_105_),
    .Y(_180_));
 sky130_fd_sc_hd__nor2_1 _627_ (.A(_107_),
    .B(_143_),
    .Y(_181_));
 sky130_fd_sc_hd__o21ai_1 _628_ (.A1(_144_),
    .A2(_181_),
    .B1(_180_),
    .Y(_182_));
 sky130_fd_sc_hd__nand3_2 _629_ (.A(_113_),
    .B(_147_),
    .C(_182_),
    .Y(_183_));
 sky130_fd_sc_hd__a21o_1 _630_ (.A1(_113_),
    .A2(_147_),
    .B1(_182_),
    .X(_184_));
 sky130_fd_sc_hd__nand3_1 _631_ (.A(_179_),
    .B(_183_),
    .C(_184_),
    .Y(_185_));
 sky130_fd_sc_hd__a21o_1 _632_ (.A1(_183_),
    .A2(_184_),
    .B1(_179_),
    .X(_186_));
 sky130_fd_sc_hd__nand3_1 _633_ (.A(_149_),
    .B(_185_),
    .C(_186_),
    .Y(_187_));
 sky130_fd_sc_hd__a21o_1 _634_ (.A1(_185_),
    .A2(_186_),
    .B1(_149_),
    .X(_188_));
 sky130_fd_sc_hd__or4bb_2 _635_ (.A(_176_),
    .B(_177_),
    .C_N(_187_),
    .D_N(_188_),
    .X(_189_));
 sky130_fd_sc_hd__a2bb2o_1 _636_ (.A1_N(_176_),
    .A2_N(_177_),
    .B1(_187_),
    .B2(_188_),
    .X(_190_));
 sky130_fd_sc_hd__a21o_1 _637_ (.A1(_189_),
    .A2(_190_),
    .B1(_164_),
    .X(_191_));
 sky130_fd_sc_hd__nand3_1 _638_ (.A(_164_),
    .B(_189_),
    .C(_190_),
    .Y(_192_));
 sky130_fd_sc_hd__a21o_1 _639_ (.A1(_191_),
    .A2(_192_),
    .B1(_155_),
    .X(_193_));
 sky130_fd_sc_hd__nand3_1 _640_ (.A(_155_),
    .B(_191_),
    .C(_192_),
    .Y(_194_));
 sky130_fd_sc_hd__and3_1 _641_ (.A(_163_),
    .B(_193_),
    .C(_194_),
    .X(_195_));
 sky130_fd_sc_hd__a21o_1 _642_ (.A1(_193_),
    .A2(_194_),
    .B1(_163_),
    .X(_196_));
 sky130_fd_sc_hd__and2b_1 _643_ (.A_N(_195_),
    .B(_196_),
    .X(_197_));
 sky130_fd_sc_hd__xnor2_2 _644_ (.A(_157_),
    .B(_197_),
    .Y(_198_));
 sky130_fd_sc_hd__o21ba_1 _645_ (.A1(_328_),
    .A2(_198_),
    .B1_N(_160_),
    .X(_199_));
 sky130_fd_sc_hd__o21a_1 _646_ (.A1(_157_),
    .A2(_195_),
    .B1(_196_),
    .X(_200_));
 sky130_fd_sc_hd__o21a_1 _647_ (.A1(_089_),
    .A2(_091_),
    .B1(_172_),
    .X(_201_));
 sky130_fd_sc_hd__o211a_1 _648_ (.A1(_336_),
    .A2(_058_),
    .B1(_087_),
    .C1(_349_),
    .X(_202_));
 sky130_fd_sc_hd__xnor2_2 _649_ (.A(_201_),
    .B(_202_),
    .Y(_203_));
 sky130_fd_sc_hd__a21bo_1 _650_ (.A1(_138_),
    .A2(_175_),
    .B1_N(_174_),
    .X(_204_));
 sky130_fd_sc_hd__xnor2_2 _651_ (.A(_203_),
    .B(_204_),
    .Y(_205_));
 sky130_fd_sc_hd__o21ai_2 _652_ (.A1(_101_),
    .A2(_105_),
    .B1(_183_),
    .Y(_206_));
 sky130_fd_sc_hd__o211a_1 _653_ (.A1(_332_),
    .A2(_068_),
    .B1(_104_),
    .C1(_344_),
    .X(_207_));
 sky130_fd_sc_hd__xnor2_2 _654_ (.A(_206_),
    .B(_207_),
    .Y(_208_));
 sky130_fd_sc_hd__a21bo_1 _655_ (.A1(_149_),
    .A2(_186_),
    .B1_N(_185_),
    .X(_209_));
 sky130_fd_sc_hd__and2b_1 _656_ (.A_N(_208_),
    .B(_209_),
    .X(_210_));
 sky130_fd_sc_hd__xor2_2 _657_ (.A(_208_),
    .B(_209_),
    .X(_211_));
 sky130_fd_sc_hd__nor2_1 _658_ (.A(_205_),
    .B(_211_),
    .Y(_212_));
 sky130_fd_sc_hd__xor2_2 _659_ (.A(_205_),
    .B(_211_),
    .X(_213_));
 sky130_fd_sc_hd__a21boi_2 _660_ (.A1(_164_),
    .A2(_189_),
    .B1_N(_190_),
    .Y(_214_));
 sky130_fd_sc_hd__xor2_1 _661_ (.A(_213_),
    .B(_214_),
    .X(_215_));
 sky130_fd_sc_hd__nand2b_1 _662_ (.A_N(_193_),
    .B(_215_),
    .Y(_216_));
 sky130_fd_sc_hd__xnor2_1 _663_ (.A(_193_),
    .B(_215_),
    .Y(_217_));
 sky130_fd_sc_hd__nor2_1 _664_ (.A(_373_),
    .B(_058_),
    .Y(_218_));
 sky130_fd_sc_hd__nor2_1 _665_ (.A(_368_),
    .B(_068_),
    .Y(_219_));
 sky130_fd_sc_hd__nor2_1 _666_ (.A(_028_),
    .B(_034_),
    .Y(_220_));
 sky130_fd_sc_hd__a211o_1 _667_ (.A1(_127_),
    .A2(_220_),
    .B1(_219_),
    .C1(_218_),
    .X(_221_));
 sky130_fd_sc_hd__nand2_1 _668_ (.A(_218_),
    .B(_219_),
    .Y(_222_));
 sky130_fd_sc_hd__o211a_1 _669_ (.A1(_218_),
    .A2(_219_),
    .B1(_220_),
    .C1(_127_),
    .X(_223_));
 sky130_fd_sc_hd__inv_2 _670_ (.A(_223_),
    .Y(_224_));
 sky130_fd_sc_hd__and3_1 _671_ (.A(_221_),
    .B(_222_),
    .C(_224_),
    .X(_225_));
 sky130_fd_sc_hd__and2_1 _672_ (.A(_217_),
    .B(_225_),
    .X(_226_));
 sky130_fd_sc_hd__or2_1 _673_ (.A(_217_),
    .B(_225_),
    .X(_227_));
 sky130_fd_sc_hd__and2b_1 _674_ (.A_N(_226_),
    .B(_227_),
    .X(_228_));
 sky130_fd_sc_hd__xnor2_2 _675_ (.A(_200_),
    .B(_228_),
    .Y(_229_));
 sky130_fd_sc_hd__o21ai_2 _676_ (.A1(_328_),
    .A2(_229_),
    .B1(_199_),
    .Y(_230_));
 sky130_fd_sc_hd__o21a_1 _677_ (.A1(_200_),
    .A2(_226_),
    .B1(_227_),
    .X(_231_));
 sky130_fd_sc_hd__o41a_1 _678_ (.A1(_350_),
    .A2(_088_),
    .A3(_130_),
    .A4(_201_),
    .B1(_165_),
    .X(_232_));
 sky130_fd_sc_hd__a21boi_2 _679_ (.A1(_203_),
    .A2(_204_),
    .B1_N(_232_),
    .Y(_233_));
 sky130_fd_sc_hd__o211a_1 _680_ (.A1(_140_),
    .A2(_206_),
    .B1(_344_),
    .C1(_104_),
    .X(_234_));
 sky130_fd_sc_hd__nor2_2 _681_ (.A(_210_),
    .B(_234_),
    .Y(_235_));
 sky130_fd_sc_hd__nor2_1 _682_ (.A(_233_),
    .B(_235_),
    .Y(_236_));
 sky130_fd_sc_hd__xor2_2 _683_ (.A(_233_),
    .B(_235_),
    .X(_237_));
 sky130_fd_sc_hd__a21oi_2 _684_ (.A1(_213_),
    .A2(_214_),
    .B1(_212_),
    .Y(_238_));
 sky130_fd_sc_hd__and2b_1 _685_ (.A_N(_238_),
    .B(_237_),
    .X(_239_));
 sky130_fd_sc_hd__xor2_2 _686_ (.A(_237_),
    .B(_238_),
    .X(_240_));
 sky130_fd_sc_hd__nor2_1 _687_ (.A(_216_),
    .B(_240_),
    .Y(_241_));
 sky130_fd_sc_hd__xor2_2 _688_ (.A(_216_),
    .B(_240_),
    .X(_242_));
 sky130_fd_sc_hd__or4_1 _689_ (.A(_373_),
    .B(_034_),
    .C(_058_),
    .D(_088_),
    .X(_243_));
 sky130_fd_sc_hd__o22ai_1 _690_ (.A1(_034_),
    .A2(_058_),
    .B1(_088_),
    .B2(_373_),
    .Y(_244_));
 sky130_fd_sc_hd__and2_1 _691_ (.A(_243_),
    .B(_244_),
    .X(_245_));
 sky130_fd_sc_hd__or4b_1 _692_ (.A(_368_),
    .B(_028_),
    .C(_068_),
    .D_N(_104_),
    .X(_246_));
 sky130_fd_sc_hd__a2bb2o_1 _693_ (.A1_N(_028_),
    .A2_N(_068_),
    .B1(_104_),
    .B2(_369_),
    .X(_247_));
 sky130_fd_sc_hd__and2_1 _694_ (.A(_246_),
    .B(_247_),
    .X(_248_));
 sky130_fd_sc_hd__nand2_1 _695_ (.A(_245_),
    .B(_248_),
    .Y(_249_));
 sky130_fd_sc_hd__nor2_1 _696_ (.A(_245_),
    .B(_248_),
    .Y(_251_));
 sky130_fd_sc_hd__or2_1 _697_ (.A(_245_),
    .B(_248_),
    .X(_252_));
 sky130_fd_sc_hd__and2_1 _698_ (.A(_249_),
    .B(_252_),
    .X(_253_));
 sky130_fd_sc_hd__xnor2_1 _699_ (.A(_222_),
    .B(_253_),
    .Y(_254_));
 sky130_fd_sc_hd__o21ai_1 _700_ (.A1(_161_),
    .A2(_223_),
    .B1(_254_),
    .Y(_255_));
 sky130_fd_sc_hd__or3_1 _701_ (.A(_161_),
    .B(_223_),
    .C(_254_),
    .X(_256_));
 sky130_fd_sc_hd__and2_1 _702_ (.A(_255_),
    .B(_256_),
    .X(_257_));
 sky130_fd_sc_hd__and2_1 _703_ (.A(_242_),
    .B(_257_),
    .X(_258_));
 sky130_fd_sc_hd__or2_1 _704_ (.A(_242_),
    .B(_257_),
    .X(_259_));
 sky130_fd_sc_hd__xor2_1 _705_ (.A(_242_),
    .B(_257_),
    .X(_260_));
 sky130_fd_sc_hd__xnor2_1 _706_ (.A(_231_),
    .B(_260_),
    .Y(_262_));
 sky130_fd_sc_hd__nor2_1 _707_ (.A(_328_),
    .B(_262_),
    .Y(_263_));
 sky130_fd_sc_hd__nor2_2 _708_ (.A(_058_),
    .B(_068_),
    .Y(_264_));
 sky130_fd_sc_hd__or3_1 _709_ (.A(_034_),
    .B(_088_),
    .C(_218_),
    .X(_265_));
 sky130_fd_sc_hd__or3b_1 _710_ (.A(_028_),
    .B(_219_),
    .C_N(_104_),
    .X(_266_));
 sky130_fd_sc_hd__or2_1 _711_ (.A(_265_),
    .B(_266_),
    .X(_267_));
 sky130_fd_sc_hd__and2_1 _712_ (.A(_265_),
    .B(_266_),
    .X(_268_));
 sky130_fd_sc_hd__nand2_1 _713_ (.A(_265_),
    .B(_266_),
    .Y(_269_));
 sky130_fd_sc_hd__nand2_1 _714_ (.A(_267_),
    .B(_269_),
    .Y(_270_));
 sky130_fd_sc_hd__o21a_1 _715_ (.A1(_222_),
    .A2(_251_),
    .B1(_249_),
    .X(_271_));
 sky130_fd_sc_hd__xnor2_1 _716_ (.A(_270_),
    .B(_271_),
    .Y(_273_));
 sky130_fd_sc_hd__nor2_1 _717_ (.A(_255_),
    .B(_273_),
    .Y(_274_));
 sky130_fd_sc_hd__and2_1 _718_ (.A(_255_),
    .B(_273_),
    .X(_275_));
 sky130_fd_sc_hd__nor2_1 _719_ (.A(_274_),
    .B(_275_),
    .Y(_276_));
 sky130_fd_sc_hd__xor2_1 _720_ (.A(_264_),
    .B(_276_),
    .X(_277_));
 sky130_fd_sc_hd__o31a_1 _721_ (.A1(_236_),
    .A2(_239_),
    .A3(_241_),
    .B1(_277_),
    .X(_278_));
 sky130_fd_sc_hd__nor4_1 _722_ (.A(_236_),
    .B(_239_),
    .C(_241_),
    .D(_277_),
    .Y(_279_));
 sky130_fd_sc_hd__or2_1 _723_ (.A(_278_),
    .B(_279_),
    .X(_280_));
 sky130_fd_sc_hd__a21o_1 _724_ (.A1(_231_),
    .A2(_259_),
    .B1(_258_),
    .X(_281_));
 sky130_fd_sc_hd__xnor2_1 _725_ (.A(_280_),
    .B(_281_),
    .Y(_282_));
 sky130_fd_sc_hd__a211o_1 _726_ (.A1(_327_),
    .A2(_282_),
    .B1(_263_),
    .C1(_230_),
    .X(_283_));
 sky130_fd_sc_hd__nand3_1 _727_ (.A(_087_),
    .B(_104_),
    .C(_264_),
    .Y(_284_));
 sky130_fd_sc_hd__nand2b_1 _728_ (.A_N(_058_),
    .B(_104_),
    .Y(_285_));
 sky130_fd_sc_hd__o21ai_1 _729_ (.A1(_068_),
    .A2(_088_),
    .B1(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__nor2_1 _730_ (.A(_243_),
    .B(_246_),
    .Y(_287_));
 sky130_fd_sc_hd__and2_1 _731_ (.A(_243_),
    .B(_246_),
    .X(_288_));
 sky130_fd_sc_hd__nor2_1 _732_ (.A(_287_),
    .B(_288_),
    .Y(_289_));
 sky130_fd_sc_hd__a21oi_1 _733_ (.A1(_249_),
    .A2(_267_),
    .B1(_268_),
    .Y(_290_));
 sky130_fd_sc_hd__o21a_1 _734_ (.A1(_289_),
    .A2(_290_),
    .B1(_274_),
    .X(_291_));
 sky130_fd_sc_hd__nor3_1 _735_ (.A(_274_),
    .B(_289_),
    .C(_290_),
    .Y(_292_));
 sky130_fd_sc_hd__nor2_1 _736_ (.A(_291_),
    .B(_292_),
    .Y(_294_));
 sky130_fd_sc_hd__and3_1 _737_ (.A(_284_),
    .B(_286_),
    .C(_294_),
    .X(_295_));
 sky130_fd_sc_hd__a21oi_1 _738_ (.A1(_284_),
    .A2(_286_),
    .B1(_294_),
    .Y(_296_));
 sky130_fd_sc_hd__nor2_1 _739_ (.A(_295_),
    .B(_296_),
    .Y(_297_));
 sky130_fd_sc_hd__and3_1 _740_ (.A(_264_),
    .B(_276_),
    .C(_297_),
    .X(_298_));
 sky130_fd_sc_hd__a21oi_1 _741_ (.A1(_264_),
    .A2(_276_),
    .B1(_297_),
    .Y(_299_));
 sky130_fd_sc_hd__nor2_1 _742_ (.A(_298_),
    .B(_299_),
    .Y(_300_));
 sky130_fd_sc_hd__a211o_1 _743_ (.A1(_231_),
    .A2(_259_),
    .B1(_278_),
    .C1(_258_),
    .X(_301_));
 sky130_fd_sc_hd__nand2b_1 _744_ (.A_N(_279_),
    .B(_301_),
    .Y(_302_));
 sky130_fd_sc_hd__and3b_1 _745_ (.A_N(_279_),
    .B(_300_),
    .C(_301_),
    .X(_303_));
 sky130_fd_sc_hd__xnor2_2 _746_ (.A(_300_),
    .B(_302_),
    .Y(_305_));
 sky130_fd_sc_hd__nor2_1 _747_ (.A(_287_),
    .B(_291_),
    .Y(_306_));
 sky130_fd_sc_hd__o211a_1 _748_ (.A1(_058_),
    .A2(_068_),
    .B1(_087_),
    .C1(_104_),
    .X(_307_));
 sky130_fd_sc_hd__xnor2_1 _749_ (.A(_306_),
    .B(_307_),
    .Y(_308_));
 sky130_fd_sc_hd__o21a_1 _750_ (.A1(_295_),
    .A2(_298_),
    .B1(_308_),
    .X(_309_));
 sky130_fd_sc_hd__nor3_1 _751_ (.A(_295_),
    .B(_298_),
    .C(_308_),
    .Y(_310_));
 sky130_fd_sc_hd__nor2_1 _752_ (.A(_309_),
    .B(_310_),
    .Y(_311_));
 sky130_fd_sc_hd__o311a_1 _753_ (.A1(_264_),
    .A2(_287_),
    .A3(_291_),
    .B1(_104_),
    .C1(_087_),
    .X(_312_));
 sky130_fd_sc_hd__a211o_1 _754_ (.A1(_303_),
    .A2(_311_),
    .B1(_312_),
    .C1(_309_),
    .X(_313_));
 sky130_fd_sc_hd__a211o_1 _755_ (.A1(_327_),
    .A2(_305_),
    .B1(_313_),
    .C1(_283_),
    .X(\FP15.d ));
 sky130_fd_sc_hd__xor2_1 _756_ (.A(_303_),
    .B(_311_),
    .X(_315_));
 sky130_fd_sc_hd__a211o_1 _757_ (.A1(_327_),
    .A2(_305_),
    .B1(_315_),
    .C1(_283_),
    .X(\FP14.d ));
 sky130_fd_sc_hd__xor2_1 _758_ (.A(_283_),
    .B(_305_),
    .X(\FP13.d ));
 sky130_fd_sc_hd__or3_1 _759_ (.A(_230_),
    .B(_263_),
    .C(_282_),
    .X(_316_));
 sky130_fd_sc_hd__o21ai_1 _760_ (.A1(_230_),
    .A2(_263_),
    .B1(_282_),
    .Y(_317_));
 sky130_fd_sc_hd__and2_1 _761_ (.A(_316_),
    .B(_317_),
    .X(\FP12.d ));
 sky130_fd_sc_hd__xnor2_1 _762_ (.A(_230_),
    .B(_262_),
    .Y(\FP11.d ));
 sky130_fd_sc_hd__xor2_1 _763_ (.A(_199_),
    .B(_229_),
    .X(\FP10.d ));
 sky130_fd_sc_hd__xnor2_1 _764_ (.A(_160_),
    .B(_198_),
    .Y(\FP9.d ));
 sky130_fd_sc_hd__xor2_1 _765_ (.A(_126_),
    .B(_159_),
    .X(\FP8.d ));
 sky130_fd_sc_hd__xor2_1 _766_ (.A(_082_),
    .B(_125_),
    .X(\FP7.d ));
 sky130_fd_sc_hd__xnor2_1 _767_ (.A(_048_),
    .B(_081_),
    .Y(\FP6.d ));
 sky130_fd_sc_hd__xor2_1 _768_ (.A(_012_),
    .B(_047_),
    .X(\FP5.d ));
 sky130_fd_sc_hd__xor2_1 _769_ (.A(_365_),
    .B(_011_),
    .X(\FP4.d ));
 sky130_fd_sc_hd__xnor2_1 _770_ (.A(_342_),
    .B(_364_),
    .Y(\FP3.d ));
 sky130_fd_sc_hd__nor2_1 _771_ (.A(_341_),
    .B(_355_),
    .Y(_319_));
 sky130_fd_sc_hd__xnor2_1 _772_ (.A(_329_),
    .B(_319_),
    .Y(\FP2.d ));
 sky130_fd_sc_hd__nand2_1 _773_ (.A(\FP0.d ),
    .B(_327_),
    .Y(_320_));
 sky130_fd_sc_hd__nor2_1 _774_ (.A(_326_),
    .B(_359_),
    .Y(_321_));
 sky130_fd_sc_hd__xnor2_1 _775_ (.A(_320_),
    .B(_321_),
    .Y(\FP1.d ));
 sky130_fd_sc_hd__dfrtp_1 _776_ (.CLK(net38),
    .D(\FP0.d ),
    .RESET_B(net36),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _777_ (.CLK(net38),
    .D(\FP1.d ),
    .RESET_B(net36),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _778_ (.CLK(net38),
    .D(\FP2.d ),
    .RESET_B(net36),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _779_ (.CLK(net39),
    .D(\FP3.d ),
    .RESET_B(net37),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _780_ (.CLK(net39),
    .D(\FP4.d ),
    .RESET_B(net37),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _781_ (.CLK(net39),
    .D(\FP5.d ),
    .RESET_B(net37),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _782_ (.CLK(net39),
    .D(\FP6.d ),
    .RESET_B(net37),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _783_ (.CLK(net39),
    .D(\FP7.d ),
    .RESET_B(net37),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _784_ (.CLK(net39),
    .D(\FP8.d ),
    .RESET_B(net37),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _785_ (.CLK(net39),
    .D(\FP9.d ),
    .RESET_B(net37),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _786_ (.CLK(net39),
    .D(\FP10.d ),
    .RESET_B(net37),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _787_ (.CLK(net39),
    .D(\FP11.d ),
    .RESET_B(net37),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _788_ (.CLK(net39),
    .D(\FP12.d ),
    .RESET_B(net37),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _789_ (.CLK(net39),
    .D(\FP13.d ),
    .RESET_B(net37),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _790_ (.CLK(net39),
    .D(\FP14.d ),
    .RESET_B(net37),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _791_ (.CLK(net39),
    .D(\FP15.d ),
    .RESET_B(net37),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_4 _792_ (.CLK(net38),
    .D(net1),
    .RESET_B(net36),
    .Q(\FA0.q ));
 sky130_fd_sc_hd__dfrtp_4 _793_ (.CLK(net38),
    .D(net2),
    .RESET_B(net36),
    .Q(\FA1.q ));
 sky130_fd_sc_hd__dfrtp_4 _794_ (.CLK(net38),
    .D(net3),
    .RESET_B(net36),
    .Q(\FA2.q ));
 sky130_fd_sc_hd__dfrtp_4 _795_ (.CLK(net38),
    .D(net4),
    .RESET_B(net36),
    .Q(\FA3.q ));
 sky130_fd_sc_hd__dfrtp_4 _796_ (.CLK(net38),
    .D(net5),
    .RESET_B(net36),
    .Q(\FA4.q ));
 sky130_fd_sc_hd__dfrtp_4 _797_ (.CLK(net38),
    .D(net6),
    .RESET_B(net36),
    .Q(\FA5.q ));
 sky130_fd_sc_hd__dfrtp_2 _798_ (.CLK(net38),
    .D(net7),
    .RESET_B(net36),
    .Q(\FA6.q ));
 sky130_fd_sc_hd__dfrtp_2 _799_ (.CLK(net38),
    .D(net8),
    .RESET_B(net36),
    .Q(\FA7.q ));
 sky130_fd_sc_hd__dfrtp_4 _800_ (.CLK(net38),
    .D(net9),
    .RESET_B(net36),
    .Q(\FB0.q ));
 sky130_fd_sc_hd__dfrtp_4 _801_ (.CLK(net38),
    .D(net10),
    .RESET_B(net36),
    .Q(\FB1.q ));
 sky130_fd_sc_hd__dfrtp_4 _802_ (.CLK(net38),
    .D(net11),
    .RESET_B(net36),
    .Q(\FB2.q ));
 sky130_fd_sc_hd__dfrtp_4 _803_ (.CLK(net38),
    .D(net12),
    .RESET_B(net36),
    .Q(\FB3.q ));
 sky130_fd_sc_hd__dfrtp_4 _804_ (.CLK(net38),
    .D(net13),
    .RESET_B(net36),
    .Q(\FB4.q ));
 sky130_fd_sc_hd__dfrtp_4 _805_ (.CLK(net38),
    .D(net14),
    .RESET_B(net36),
    .Q(\FB5.q ));
 sky130_fd_sc_hd__dfrtp_4 _806_ (.CLK(net38),
    .D(net15),
    .RESET_B(net36),
    .Q(\FB6.q ));
 sky130_fd_sc_hd__dfrtp_4 _807_ (.CLK(net38),
    .D(net16),
    .RESET_B(net36),
    .Q(\FB7.q ));
 sky130_fd_sc_hd__dfrtp_4 _808_ (.CLK(net38),
    .D(net18),
    .RESET_B(net36),
    .Q(\FC.q ));
 sky130_fd_sc_hd__buf_6 fanout36 (.A(net19),
    .X(net36));
 sky130_fd_sc_hd__buf_4 fanout37 (.A(net19),
    .X(net37));
 sky130_fd_sc_hd__buf_4 fanout38 (.A(net17),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net17),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(clk),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(control),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(rst),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(p[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(p[10]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(p[11]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(p[12]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(p[13]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(p[14]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(p[15]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(p[1]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(p[2]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(p[3]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(p[4]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(p[5]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(p[6]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(p[7]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(p[8]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(p[9]));
endmodule

