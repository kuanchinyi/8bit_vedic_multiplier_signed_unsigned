// This is the unpowered netlist.
module vmsu_8bit_top (clk,
    control,
    rst,
    a,
    b,
    p);
 input clk;
 input control;
 input rst;
 input [7:0] a;
 input [7:0] b;
 output [15:0] p;

 wire \FA0.q ;
 wire \FA1.q ;
 wire \FA2.q ;
 wire \FA3.q ;
 wire \FA4.q ;
 wire \FA5.q ;
 wire \FA6.q ;
 wire \FA7.q ;
 wire \FB0.q ;
 wire \FB1.q ;
 wire \FB2.q ;
 wire \FB3.q ;
 wire \FB4.q ;
 wire \FB5.q ;
 wire \FB6.q ;
 wire \FB7.q ;
 wire \FC.q ;
 wire \FP0.d ;
 wire \FP1.d ;
 wire \FP10.d ;
 wire \FP11.d ;
 wire \FP12.d ;
 wire \FP13.d ;
 wire \FP14.d ;
 wire \FP15.d ;
 wire \FP2.d ;
 wire \FP3.d ;
 wire \FP4.d ;
 wire \FP5.d ;
 wire \FP6.d ;
 wire \FP7.d ;
 wire \FP8.d ;
 wire \FP9.d ;
 wire \M0.FAM0.d ;
 wire \M0.FAM0.q ;
 wire \M0.FAM1.d ;
 wire \M0.FAM1.q ;
 wire \M0.FAM2.d ;
 wire \M0.FAM2.q ;
 wire \M0.FAM3.d ;
 wire \M0.FAM3.q ;
 wire \M0.FAM4.d ;
 wire \M0.FAM4.q ;
 wire \M0.FAM5.d ;
 wire \M0.FAM5.q ;
 wire \M0.FAM6.d ;
 wire \M0.FAM6.q ;
 wire \M0.FAM7.d ;
 wire \M0.FAM7.q ;
 wire \M0.FBM0.d ;
 wire \M0.FBM0.q ;
 wire \M0.FBM1.d ;
 wire \M0.FBM1.q ;
 wire \M0.FBM2.d ;
 wire \M0.FBM2.q ;
 wire \M0.FBM3.d ;
 wire \M0.FBM3.q ;
 wire \M0.FBM4.d ;
 wire \M0.FBM4.q ;
 wire \M0.FBM5.d ;
 wire \M0.FBM5.q ;
 wire \M0.FBM6.d ;
 wire \M0.FBM6.q ;
 wire \M0.FBM7.d ;
 wire \M0.FBM7.q ;
 wire \M0.FCM1.d ;
 wire \M0.FCM1.q ;
 wire \M0.FCM2.d ;
 wire \M0.FCM2.q ;
 wire \M0.FCM3.q ;
 wire \M0.FCM4.q ;
 wire \M0.FPM0.d ;
 wire \M0.FPM0.q ;
 wire \M0.FPM1.d ;
 wire \M0.FPM1.q ;
 wire \M0.FPM10.d ;
 wire \M0.FPM10.q ;
 wire \M0.FPM11.d ;
 wire \M0.FPM11.q ;
 wire \M0.FPM12.d ;
 wire \M0.FPM12.q ;
 wire \M0.FPM13.d ;
 wire \M0.FPM13.q ;
 wire \M0.FPM14.d ;
 wire \M0.FPM14.q ;
 wire \M0.FPM15.d ;
 wire \M0.FPM15.q ;
 wire \M0.FPM2.d ;
 wire \M0.FPM2.q ;
 wire \M0.FPM3.d ;
 wire \M0.FPM3.q ;
 wire \M0.FPM4.d ;
 wire \M0.FPM4.q ;
 wire \M0.FPM5.d ;
 wire \M0.FPM5.q ;
 wire \M0.FPM6.d ;
 wire \M0.FPM6.q ;
 wire \M0.FPM7.d ;
 wire \M0.FPM7.q ;
 wire \M0.FPM8.d ;
 wire \M0.FPM8.q ;
 wire \M0.FPM9.d ;
 wire \M0.FPM9.q ;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net6;
 wire net7;
 wire net8;
 wire net9;

 sky130_fd_sc_hd__diode_2 ANTENNA__0648__B1 (.DIODE(_0100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0650__A (.DIODE(_0100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0652__B1 (.DIODE(_0100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0654__B1 (.DIODE(_0100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0656__B (.DIODE(_0100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0663__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__B (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__C (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0668__D (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__C (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0669__D (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__C (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0670__D (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0672__B (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0673__B (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0674__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__A1 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0675__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0678__B (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0679__B (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0681__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0682__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0683__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0684__B (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0692__B (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0693__B (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0698__A2 (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0700__A2 (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0701__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0702__B (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0713__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0716__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0719__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__A (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0721__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0724__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0726__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__A (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0729__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0730__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0732__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0733__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0737__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__A (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0739__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__C (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0740__D (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__C (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0745__D (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0746__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0749__A (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0750__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0751__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0752__A1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__A1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__A2 (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0756__B1 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__A1 (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0757__A2 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__A_N (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__C (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0772__D (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A1 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__A2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0773__B1_N (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0774__B1_N (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0775__C (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__A1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0776__B1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0777__B1 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A1 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__A2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0778__B1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0779__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0780__A1 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0781__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0782__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0786__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0787__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0789__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0810__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0814__A (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0815__B (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0816__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__A1 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0818__A2 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0821__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0822__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0823__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A1 (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0824__A3 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__A (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0825__B_N (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0826__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0827__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0828__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__A2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0829__B1 (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__A_N (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__C (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0831__D (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0833__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__A2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0834__B1 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__C (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0836__D (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0837__B_N (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A1 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__A2 (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0838__B1_N (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0839__C (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__A1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0840__C1 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A1 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__A2 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0850__B1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0851__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0852__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__A_N (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__C (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0853__D (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A1 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__A2 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0854__B1_N (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0855__B1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0856__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A1 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0857__A2 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0859__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0860__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0863__B1 (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0864__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0868__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0869__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0871__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0872__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0877__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0878__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0897__B (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0898__B (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0899__C1 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0900__A1 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0910__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0914__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0915__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__B (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__C (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0917__D (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0918__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0919__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0921__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0922__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0923__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__A (.DIODE(_0121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0938__B (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0939__B (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0952__B (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0953__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__0970__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0971__A (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0974__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0978__B_N (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0979__B (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0980__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0994__A1 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0995__B (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0996__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0997__A (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A1_N (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__0998__A2_N (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1000__A1 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A1 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A2 (.DIODE(_0124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A3 (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1008__A4 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1009__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__A (.DIODE(_0117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1013__B (.DIODE(_0172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__A1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1031__B1 (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1032__A1 (.DIODE(_0119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1033__A (.DIODE(\M0.FBM7.q ));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__A1 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1035__B1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1036__B1 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1107__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__A1 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1108__S (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1109__A (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1111__B2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__A (.DIODE(_0175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1113__B (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__A (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1114__B (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__A (.DIODE(_0171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1117__C (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A1 (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__A2 (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1119__B2 (.DIODE(_0177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1120__A (.DIODE(_0169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1121__A3 (.DIODE(_0180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1122__A1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1134__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1135__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1136__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1137__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1138__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1139__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1140__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1141__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1142__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1143__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1144__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1145__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1146__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1147__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1148__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1149__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1150__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1151__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1152__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1153__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1154__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1155__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1156__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1157__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1158__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1159__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1160__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1161__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1162__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1163__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1164__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1165__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1166__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1167__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1168__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1169__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1170__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1171__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1172__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1173__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1174__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1175__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1176__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1177__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1178__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1179__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1180__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1181__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1182__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1183__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1184__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1185__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1186__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1187__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1188__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1189__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1190__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1191__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1192__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1193__A (.DIODE(_0577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1194__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1195__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1196__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1197__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1198__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1199__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1200__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1201__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1202__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1203__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1204__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1205__A (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__1206__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1207__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1208__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1209__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1210__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1211__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1212__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1213__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1214__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1215__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1216__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1217__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1218__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1219__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1220__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1221__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1222__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1223__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1224__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1225__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1226__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1227__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1228__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1229__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1230__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1231__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1232__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1233__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1234__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1235__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1236__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1237__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1238__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1239__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1240__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1241__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1242__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1243__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1244__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1245__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1246__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1247__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1248__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1249__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1250__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1251__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1252__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1253__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1254__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1255__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1256__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1257__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1258__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1259__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1260__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1261__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1262__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1263__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1264__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1265__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1266__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1267__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1268__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1269__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1270__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1271__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1272__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1273__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__1274__CLK (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap49_A (.DIODE(_0100_));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_226 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_6 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_18 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_340 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_344 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__and2_1 _0578_ (.A(\FC.q ),
    .B(\FB7.q ),
    .X(_0069_));
 sky130_fd_sc_hd__clkbuf_2 _0579_ (.A(_0069_),
    .X(\M0.FCM2.d ));
 sky130_fd_sc_hd__or4_1 _0580_ (.A(\FB0.q ),
    .B(\FB1.q ),
    .C(\FB2.q ),
    .D(\FB3.q ),
    .X(_0070_));
 sky130_fd_sc_hd__or3_1 _0581_ (.A(\FB4.q ),
    .B(\FB5.q ),
    .C(_0070_),
    .X(_0071_));
 sky130_fd_sc_hd__o21ai_1 _0582_ (.A1(\FB6.q ),
    .A2(_0071_),
    .B1(\FC.q ),
    .Y(_0072_));
 sky130_fd_sc_hd__and2_1 _0583_ (.A(\FB7.q ),
    .B(_0072_),
    .X(_0073_));
 sky130_fd_sc_hd__clkbuf_1 _0584_ (.A(_0073_),
    .X(\M0.FBM7.d ));
 sky130_fd_sc_hd__and2_1 _0585_ (.A(\M0.FCM2.d ),
    .B(_0071_),
    .X(_0074_));
 sky130_fd_sc_hd__xor2_1 _0586_ (.A(\FB6.q ),
    .B(_0074_),
    .X(\M0.FBM6.d ));
 sky130_fd_sc_hd__o21ai_1 _0587_ (.A1(\FB4.q ),
    .A2(_0070_),
    .B1(\M0.FCM2.d ),
    .Y(_0075_));
 sky130_fd_sc_hd__xnor2_1 _0588_ (.A(\FB5.q ),
    .B(_0075_),
    .Y(\M0.FBM5.d ));
 sky130_fd_sc_hd__nand2_1 _0589_ (.A(\M0.FCM2.d ),
    .B(_0070_),
    .Y(_0076_));
 sky130_fd_sc_hd__xnor2_1 _0590_ (.A(\FB4.q ),
    .B(_0076_),
    .Y(\M0.FBM4.d ));
 sky130_fd_sc_hd__o31a_1 _0591_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .A3(\FB2.q ),
    .B1(\M0.FCM2.d ),
    .X(_0077_));
 sky130_fd_sc_hd__xor2_1 _0592_ (.A(\FB3.q ),
    .B(_0077_),
    .X(\M0.FBM3.d ));
 sky130_fd_sc_hd__o21a_1 _0593_ (.A1(\FB0.q ),
    .A2(\FB1.q ),
    .B1(\M0.FCM2.d ),
    .X(_0078_));
 sky130_fd_sc_hd__xor2_1 _0594_ (.A(\FB2.q ),
    .B(_0078_),
    .X(\M0.FBM2.d ));
 sky130_fd_sc_hd__and3_1 _0595_ (.A(\FC.q ),
    .B(\FB7.q ),
    .C(\FB0.q ),
    .X(_0079_));
 sky130_fd_sc_hd__xor2_1 _0596_ (.A(\FB1.q ),
    .B(_0079_),
    .X(\M0.FBM1.d ));
 sky130_fd_sc_hd__clkbuf_1 _0597_ (.A(\FB0.q ),
    .X(_0080_));
 sky130_fd_sc_hd__clkbuf_1 _0598_ (.A(_0080_),
    .X(\M0.FBM0.d ));
 sky130_fd_sc_hd__and2_1 _0599_ (.A(\FC.q ),
    .B(\FA7.q ),
    .X(_0081_));
 sky130_fd_sc_hd__clkbuf_2 _0600_ (.A(_0081_),
    .X(\M0.FCM1.d ));
 sky130_fd_sc_hd__or4_2 _0601_ (.A(\FA0.q ),
    .B(\FA1.q ),
    .C(\FA2.q ),
    .D(\FA3.q ),
    .X(_0082_));
 sky130_fd_sc_hd__or3_1 _0602_ (.A(\FA4.q ),
    .B(\FA5.q ),
    .C(_0082_),
    .X(_0083_));
 sky130_fd_sc_hd__o21ai_1 _0603_ (.A1(\FA6.q ),
    .A2(_0083_),
    .B1(\FC.q ),
    .Y(_0084_));
 sky130_fd_sc_hd__and2_1 _0604_ (.A(\FA7.q ),
    .B(_0084_),
    .X(_0085_));
 sky130_fd_sc_hd__clkbuf_1 _0605_ (.A(_0085_),
    .X(\M0.FAM7.d ));
 sky130_fd_sc_hd__and2_1 _0606_ (.A(\M0.FCM1.d ),
    .B(_0083_),
    .X(_0086_));
 sky130_fd_sc_hd__xor2_1 _0607_ (.A(\FA6.q ),
    .B(_0086_),
    .X(\M0.FAM6.d ));
 sky130_fd_sc_hd__o21ai_1 _0608_ (.A1(\FA4.q ),
    .A2(_0082_),
    .B1(\M0.FCM1.d ),
    .Y(_0087_));
 sky130_fd_sc_hd__xnor2_1 _0609_ (.A(\FA5.q ),
    .B(_0087_),
    .Y(\M0.FAM5.d ));
 sky130_fd_sc_hd__nand2_1 _0610_ (.A(\M0.FCM1.d ),
    .B(_0082_),
    .Y(_0088_));
 sky130_fd_sc_hd__xnor2_1 _0611_ (.A(\FA4.q ),
    .B(_0088_),
    .Y(\M0.FAM4.d ));
 sky130_fd_sc_hd__o31a_1 _0612_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .A3(\FA2.q ),
    .B1(\M0.FCM1.d ),
    .X(_0089_));
 sky130_fd_sc_hd__xor2_1 _0613_ (.A(\FA3.q ),
    .B(_0089_),
    .X(\M0.FAM3.d ));
 sky130_fd_sc_hd__o21a_1 _0614_ (.A1(\FA0.q ),
    .A2(\FA1.q ),
    .B1(\M0.FCM1.d ),
    .X(_0090_));
 sky130_fd_sc_hd__xor2_1 _0615_ (.A(\FA2.q ),
    .B(_0090_),
    .X(\M0.FAM2.d ));
 sky130_fd_sc_hd__and3_1 _0616_ (.A(\FC.q ),
    .B(\FA7.q ),
    .C(\FA0.q ),
    .X(_0091_));
 sky130_fd_sc_hd__xor2_1 _0617_ (.A(\FA1.q ),
    .B(_0091_),
    .X(\M0.FAM1.d ));
 sky130_fd_sc_hd__clkbuf_1 _0618_ (.A(\FA0.q ),
    .X(_0092_));
 sky130_fd_sc_hd__clkbuf_1 _0619_ (.A(_0092_),
    .X(\M0.FAM0.d ));
 sky130_fd_sc_hd__or4_1 _0620_ (.A(\M0.FPM0.q ),
    .B(\M0.FPM1.q ),
    .C(\M0.FPM2.q ),
    .D(\M0.FPM3.q ),
    .X(_0093_));
 sky130_fd_sc_hd__or3_1 _0621_ (.A(\M0.FPM4.q ),
    .B(\M0.FPM5.q ),
    .C(_0093_),
    .X(_0094_));
 sky130_fd_sc_hd__or2_1 _0622_ (.A(\M0.FPM6.q ),
    .B(_0094_),
    .X(_0095_));
 sky130_fd_sc_hd__or3_1 _0623_ (.A(\M0.FPM7.q ),
    .B(\M0.FPM8.q ),
    .C(_0095_),
    .X(_0096_));
 sky130_fd_sc_hd__or2_1 _0624_ (.A(\M0.FPM9.q ),
    .B(_0096_),
    .X(_0097_));
 sky130_fd_sc_hd__or3_1 _0625_ (.A(\M0.FPM10.q ),
    .B(\M0.FPM11.q ),
    .C(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__or2_1 _0626_ (.A(\M0.FPM12.q ),
    .B(_0098_),
    .X(_0099_));
 sky130_fd_sc_hd__xor2_4 _0627_ (.A(\M0.FCM3.q ),
    .B(\M0.FCM4.q ),
    .X(_0100_));
 sky130_fd_sc_hd__o31a_1 _0628_ (.A1(\M0.FPM14.q ),
    .A2(\M0.FPM13.q ),
    .A3(_0099_),
    .B1(net49),
    .X(_0101_));
 sky130_fd_sc_hd__xor2_1 _0629_ (.A(\M0.FPM15.q ),
    .B(_0101_),
    .X(\FP15.d ));
 sky130_fd_sc_hd__o21ai_1 _0630_ (.A1(\M0.FPM13.q ),
    .A2(_0099_),
    .B1(net49),
    .Y(_0102_));
 sky130_fd_sc_hd__xnor2_1 _0631_ (.A(\M0.FPM14.q ),
    .B(_0102_),
    .Y(\FP14.d ));
 sky130_fd_sc_hd__nand2_1 _0632_ (.A(net49),
    .B(_0099_),
    .Y(_0103_));
 sky130_fd_sc_hd__xnor2_1 _0633_ (.A(\M0.FPM13.q ),
    .B(_0103_),
    .Y(\FP13.d ));
 sky130_fd_sc_hd__nand2_1 _0634_ (.A(net49),
    .B(_0098_),
    .Y(_0104_));
 sky130_fd_sc_hd__xnor2_1 _0635_ (.A(\M0.FPM12.q ),
    .B(_0104_),
    .Y(\FP12.d ));
 sky130_fd_sc_hd__o21ai_1 _0636_ (.A1(\M0.FPM10.q ),
    .A2(_0097_),
    .B1(net49),
    .Y(_0105_));
 sky130_fd_sc_hd__xnor2_1 _0637_ (.A(\M0.FPM11.q ),
    .B(_0105_),
    .Y(\FP11.d ));
 sky130_fd_sc_hd__nand2_1 _0638_ (.A(net49),
    .B(_0097_),
    .Y(_0106_));
 sky130_fd_sc_hd__xnor2_1 _0639_ (.A(\M0.FPM10.q ),
    .B(_0106_),
    .Y(\FP10.d ));
 sky130_fd_sc_hd__nand2_1 _0640_ (.A(net49),
    .B(_0096_),
    .Y(_0107_));
 sky130_fd_sc_hd__xnor2_1 _0641_ (.A(\M0.FPM9.q ),
    .B(_0107_),
    .Y(\FP9.d ));
 sky130_fd_sc_hd__o21ai_1 _0642_ (.A1(\M0.FPM7.q ),
    .A2(_0095_),
    .B1(net49),
    .Y(_0108_));
 sky130_fd_sc_hd__xnor2_1 _0643_ (.A(\M0.FPM8.q ),
    .B(_0108_),
    .Y(\FP8.d ));
 sky130_fd_sc_hd__nand2_1 _0644_ (.A(net49),
    .B(_0095_),
    .Y(_0109_));
 sky130_fd_sc_hd__xnor2_1 _0645_ (.A(\M0.FPM7.q ),
    .B(_0109_),
    .Y(\FP7.d ));
 sky130_fd_sc_hd__nand2_1 _0646_ (.A(net49),
    .B(_0094_),
    .Y(_0110_));
 sky130_fd_sc_hd__xnor2_1 _0647_ (.A(\M0.FPM6.q ),
    .B(_0110_),
    .Y(\FP6.d ));
 sky130_fd_sc_hd__o21ai_1 _0648_ (.A1(\M0.FPM4.q ),
    .A2(_0093_),
    .B1(_0100_),
    .Y(_0111_));
 sky130_fd_sc_hd__xnor2_1 _0649_ (.A(\M0.FPM5.q ),
    .B(_0111_),
    .Y(\FP5.d ));
 sky130_fd_sc_hd__nand2_1 _0650_ (.A(_0100_),
    .B(_0093_),
    .Y(_0112_));
 sky130_fd_sc_hd__xnor2_1 _0651_ (.A(\M0.FPM4.q ),
    .B(_0112_),
    .Y(\FP4.d ));
 sky130_fd_sc_hd__o31a_1 _0652_ (.A1(\M0.FPM0.q ),
    .A2(\M0.FPM1.q ),
    .A3(\M0.FPM2.q ),
    .B1(_0100_),
    .X(_0113_));
 sky130_fd_sc_hd__xor2_1 _0653_ (.A(\M0.FPM3.q ),
    .B(_0113_),
    .X(\FP3.d ));
 sky130_fd_sc_hd__o21ai_1 _0654_ (.A1(\M0.FPM0.q ),
    .A2(\M0.FPM1.q ),
    .B1(_0100_),
    .Y(_0114_));
 sky130_fd_sc_hd__xnor2_1 _0655_ (.A(\M0.FPM2.q ),
    .B(_0114_),
    .Y(\FP2.d ));
 sky130_fd_sc_hd__nand2_1 _0656_ (.A(\M0.FPM0.q ),
    .B(_0100_),
    .Y(_0115_));
 sky130_fd_sc_hd__xnor2_1 _0657_ (.A(\M0.FPM1.q ),
    .B(_0115_),
    .Y(\FP1.d ));
 sky130_fd_sc_hd__clkbuf_1 _0658_ (.A(\M0.FPM0.q ),
    .X(_0116_));
 sky130_fd_sc_hd__clkbuf_1 _0659_ (.A(_0116_),
    .X(\FP0.d ));
 sky130_fd_sc_hd__buf_4 _0660_ (.A(\M0.FAM7.q ),
    .X(_0117_));
 sky130_fd_sc_hd__clkbuf_8 _0661_ (.A(\M0.FAM6.q ),
    .X(_0118_));
 sky130_fd_sc_hd__buf_6 _0662_ (.A(\M0.FBM6.q ),
    .X(_0119_));
 sky130_fd_sc_hd__and2_1 _0663_ (.A(_0118_),
    .B(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_4 _0664_ (.A(\M0.FAM5.q ),
    .X(_0121_));
 sky130_fd_sc_hd__buf_8 _0665_ (.A(\M0.FAM4.q ),
    .X(_0122_));
 sky130_fd_sc_hd__clkbuf_8 _0666_ (.A(\M0.FBM5.q ),
    .X(_0123_));
 sky130_fd_sc_hd__buf_6 _0667_ (.A(\M0.FBM4.q ),
    .X(_0124_));
 sky130_fd_sc_hd__and4_1 _0668_ (.A(_0121_),
    .B(_0122_),
    .C(_0123_),
    .D(_0124_),
    .X(_0125_));
 sky130_fd_sc_hd__and4_1 _0669_ (.A(\M0.FBM7.q ),
    .B(_0119_),
    .C(_0121_),
    .D(_0122_),
    .X(_0126_));
 sky130_fd_sc_hd__and4_1 _0670_ (.A(_0117_),
    .B(_0118_),
    .C(_0123_),
    .D(_0124_),
    .X(_0127_));
 sky130_fd_sc_hd__xnor2_1 _0671_ (.A(_0126_),
    .B(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__nand2_1 _0672_ (.A(_0121_),
    .B(_0123_),
    .Y(_0129_));
 sky130_fd_sc_hd__nand2_1 _0673_ (.A(_0119_),
    .B(_0122_),
    .Y(_0130_));
 sky130_fd_sc_hd__nand2_1 _0674_ (.A(_0118_),
    .B(_0124_),
    .Y(_0131_));
 sky130_fd_sc_hd__o22a_1 _0675_ (.A1(_0124_),
    .A2(_0130_),
    .B1(_0131_),
    .B2(_0122_),
    .X(_0132_));
 sky130_fd_sc_hd__nor2_1 _0676_ (.A(_0129_),
    .B(_0132_),
    .Y(_0133_));
 sky130_fd_sc_hd__nor2_1 _0677_ (.A(_0125_),
    .B(_0133_),
    .Y(_0134_));
 sky130_fd_sc_hd__nand2_1 _0678_ (.A(\M0.FBM7.q ),
    .B(_0122_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _0679_ (.A(_0119_),
    .B(_0121_),
    .Y(_0136_));
 sky130_fd_sc_hd__xor2_1 _0680_ (.A(_0135_),
    .B(_0136_),
    .X(_0137_));
 sky130_fd_sc_hd__nand2_2 _0681_ (.A(_0122_),
    .B(_0124_),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _0682_ (.A(_0118_),
    .B(_0119_),
    .Y(_0139_));
 sky130_fd_sc_hd__nand2_1 _0683_ (.A(_0117_),
    .B(_0124_),
    .Y(_0140_));
 sky130_fd_sc_hd__nand2_1 _0684_ (.A(_0118_),
    .B(_0123_),
    .Y(_0141_));
 sky130_fd_sc_hd__xnor2_1 _0685_ (.A(_0140_),
    .B(_0141_),
    .Y(_0142_));
 sky130_fd_sc_hd__nor3_1 _0686_ (.A(_0138_),
    .B(_0139_),
    .C(_0142_),
    .Y(_0143_));
 sky130_fd_sc_hd__o21ai_1 _0687_ (.A1(_0138_),
    .A2(_0139_),
    .B1(_0142_),
    .Y(_0144_));
 sky130_fd_sc_hd__and2b_1 _0688_ (.A_N(_0143_),
    .B(_0144_),
    .X(_0145_));
 sky130_fd_sc_hd__xnor2_1 _0689_ (.A(_0137_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__nor2_2 _0690_ (.A(_0134_),
    .B(_0146_),
    .Y(_0147_));
 sky130_fd_sc_hd__o21a_1 _0691_ (.A1(_0137_),
    .A2(_0143_),
    .B1(_0144_),
    .X(_0148_));
 sky130_fd_sc_hd__and3_1 _0692_ (.A(_0117_),
    .B(_0123_),
    .C(_0131_),
    .X(_0149_));
 sky130_fd_sc_hd__and3_1 _0693_ (.A(\M0.FBM7.q ),
    .B(_0121_),
    .C(_0130_),
    .X(_0150_));
 sky130_fd_sc_hd__xnor2_1 _0694_ (.A(_0149_),
    .B(_0150_),
    .Y(_0151_));
 sky130_fd_sc_hd__xnor2_2 _0695_ (.A(_0148_),
    .B(_0151_),
    .Y(_0152_));
 sky130_fd_sc_hd__and3b_1 _0696_ (.A_N(_0128_),
    .B(_0147_),
    .C(_0152_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_1 _0697_ (.A(_0125_),
    .B(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__a31o_1 _0698_ (.A1(_0117_),
    .A2(\M0.FBM7.q ),
    .A3(_0120_),
    .B1(_0154_),
    .X(_0155_));
 sky130_fd_sc_hd__o21ba_1 _0699_ (.A1(_0125_),
    .A2(_0139_),
    .B1_N(_0154_),
    .X(_0156_));
 sky130_fd_sc_hd__a32o_1 _0700_ (.A1(_0117_),
    .A2(\M0.FBM7.q ),
    .A3(_0156_),
    .B1(_0153_),
    .B2(_0133_),
    .X(_0157_));
 sky130_fd_sc_hd__nand2_1 _0701_ (.A(_0117_),
    .B(_0119_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(\M0.FBM7.q ),
    .B(_0118_),
    .Y(_0159_));
 sky130_fd_sc_hd__xnor2_1 _0703_ (.A(_0158_),
    .B(_0159_),
    .Y(_0160_));
 sky130_fd_sc_hd__or2_1 _0704_ (.A(_0147_),
    .B(_0150_),
    .X(_0161_));
 sky130_fd_sc_hd__a21o_1 _0705_ (.A1(_0147_),
    .A2(_0150_),
    .B1(_0149_),
    .X(_0162_));
 sky130_fd_sc_hd__a21o_1 _0706_ (.A1(_0161_),
    .A2(_0162_),
    .B1(_0148_),
    .X(_0163_));
 sky130_fd_sc_hd__o21ai_1 _0707_ (.A1(_0149_),
    .A2(_0161_),
    .B1(_0163_),
    .Y(_0164_));
 sky130_fd_sc_hd__a21o_1 _0708_ (.A1(_0128_),
    .A2(_0164_),
    .B1(_0153_),
    .X(_0165_));
 sky130_fd_sc_hd__nor2_1 _0709_ (.A(_0160_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__nand2_1 _0710_ (.A(_0157_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__buf_6 _0711_ (.A(\M0.FAM3.q ),
    .X(_0168_));
 sky130_fd_sc_hd__buf_8 _0712_ (.A(\M0.FBM2.q ),
    .X(_0169_));
 sky130_fd_sc_hd__nand2_2 _0713_ (.A(_0168_),
    .B(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__buf_8 _0714_ (.A(\M0.FAM2.q ),
    .X(_0171_));
 sky130_fd_sc_hd__buf_4 _0715_ (.A(\M0.FBM3.q ),
    .X(_0172_));
 sky130_fd_sc_hd__nand2_2 _0716_ (.A(_0171_),
    .B(_0172_),
    .Y(_0173_));
 sky130_fd_sc_hd__xnor2_4 _0717_ (.A(_0170_),
    .B(_0173_),
    .Y(_0174_));
 sky130_fd_sc_hd__buf_6 _0718_ (.A(\M0.FAM1.q ),
    .X(_0175_));
 sky130_fd_sc_hd__nand2_2 _0719_ (.A(_0175_),
    .B(_0169_),
    .Y(_0176_));
 sky130_fd_sc_hd__buf_6 _0720_ (.A(\M0.FAM0.q ),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_2 _0721_ (.A(_0177_),
    .B(_0172_),
    .Y(_0178_));
 sky130_fd_sc_hd__xor2_4 _0722_ (.A(_0176_),
    .B(_0178_),
    .X(_0179_));
 sky130_fd_sc_hd__buf_8 _0723_ (.A(\M0.FBM0.q ),
    .X(_0180_));
 sky130_fd_sc_hd__nand2_2 _0724_ (.A(_0168_),
    .B(_0180_),
    .Y(_0181_));
 sky130_fd_sc_hd__clkbuf_8 _0725_ (.A(\M0.FBM1.q ),
    .X(_0182_));
 sky130_fd_sc_hd__nand2_2 _0726_ (.A(_0171_),
    .B(_0182_),
    .Y(_0183_));
 sky130_fd_sc_hd__xor2_4 _0727_ (.A(_0181_),
    .B(_0183_),
    .X(_0184_));
 sky130_fd_sc_hd__nand2_2 _0728_ (.A(_0179_),
    .B(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__and2_2 _0729_ (.A(_0177_),
    .B(_0169_),
    .X(_0186_));
 sky130_fd_sc_hd__nand2_2 _0730_ (.A(_0175_),
    .B(_0172_),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _0731_ (.A(_0186_),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__nand2_2 _0732_ (.A(_0168_),
    .B(_0182_),
    .Y(_0189_));
 sky130_fd_sc_hd__and2_1 _0733_ (.A(_0171_),
    .B(_0180_),
    .X(_0190_));
 sky130_fd_sc_hd__buf_2 _0734_ (.A(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_1 _0735_ (.A(_0189_),
    .B(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__xnor2_1 _0736_ (.A(_0188_),
    .B(_0192_),
    .Y(_0193_));
 sky130_fd_sc_hd__nand2_1 _0737_ (.A(_0171_),
    .B(_0180_),
    .Y(_0194_));
 sky130_fd_sc_hd__or4b_1 _0738_ (.A(_0184_),
    .B(_0186_),
    .C(_0194_),
    .D_N(_0187_),
    .X(_0195_));
 sky130_fd_sc_hd__nand2_4 _0739_ (.A(_0177_),
    .B(_0169_),
    .Y(_0196_));
 sky130_fd_sc_hd__and4_1 _0740_ (.A(_0168_),
    .B(_0175_),
    .C(_0172_),
    .D(_0182_),
    .X(_0197_));
 sky130_fd_sc_hd__and3_1 _0741_ (.A(_0196_),
    .B(_0194_),
    .C(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__o211a_1 _0742_ (.A1(_0186_),
    .A2(_0187_),
    .B1(_0194_),
    .C1(_0189_),
    .X(_0199_));
 sky130_fd_sc_hd__o2bb2ai_1 _0743_ (.A1_N(_0179_),
    .A2_N(_0184_),
    .B1(_0198_),
    .B2(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__o211a_2 _0744_ (.A1(_0185_),
    .A2(_0193_),
    .B1(_0195_),
    .C1(_0200_),
    .X(_0201_));
 sky130_fd_sc_hd__and4_1 _0745_ (.A(_0171_),
    .B(_0177_),
    .C(_0169_),
    .D(_0180_),
    .X(_0202_));
 sky130_fd_sc_hd__and2_1 _0746_ (.A(_0175_),
    .B(_0182_),
    .X(_0203_));
 sky130_fd_sc_hd__and2_1 _0747_ (.A(_0202_),
    .B(_0203_),
    .X(_0204_));
 sky130_fd_sc_hd__xnor2_1 _0748_ (.A(_0196_),
    .B(_0191_),
    .Y(_0205_));
 sky130_fd_sc_hd__inv_2 _0749_ (.A(_0180_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand2_1 _0750_ (.A(_0175_),
    .B(_0182_),
    .Y(_0207_));
 sky130_fd_sc_hd__nor2_1 _0751_ (.A(_0171_),
    .B(_0177_),
    .Y(_0208_));
 sky130_fd_sc_hd__a2111o_1 _0752_ (.A1(_0206_),
    .A2(_0196_),
    .B1(_0202_),
    .C1(_0207_),
    .D1(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__a21oi_1 _0753_ (.A1(_0197_),
    .A2(_0205_),
    .B1(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__xor2_4 _0754_ (.A(_0179_),
    .B(_0184_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_2 _0755_ (.A0(_0204_),
    .A1(_0210_),
    .S(_0211_),
    .X(_0212_));
 sky130_fd_sc_hd__a21o_1 _0756_ (.A1(_0177_),
    .A2(_0172_),
    .B1(_0175_),
    .X(_0213_));
 sky130_fd_sc_hd__o221a_1 _0757_ (.A1(_0172_),
    .A2(_0169_),
    .B1(_0176_),
    .B2(_0178_),
    .C1(_0213_),
    .X(_0214_));
 sky130_fd_sc_hd__a211o_2 _0758_ (.A1(_0184_),
    .A2(_0186_),
    .B1(_0194_),
    .C1(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__and2_1 _0759_ (.A(_0189_),
    .B(_0187_),
    .X(_0216_));
 sky130_fd_sc_hd__a31oi_4 _0760_ (.A1(_0185_),
    .A2(_0196_),
    .A3(_0189_),
    .B1(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__a21o_1 _0761_ (.A1(_0179_),
    .A2(_0184_),
    .B1(_0188_),
    .X(_0218_));
 sky130_fd_sc_hd__a21oi_1 _0762_ (.A1(_0191_),
    .A2(_0187_),
    .B1(_0189_),
    .Y(_0219_));
 sky130_fd_sc_hd__o41ai_1 _0763_ (.A1(_0179_),
    .A2(_0184_),
    .A3(_0187_),
    .A4(_0202_),
    .B1(_0219_),
    .Y(_0220_));
 sky130_fd_sc_hd__and3_1 _0764_ (.A(_0179_),
    .B(_0184_),
    .C(_0196_),
    .X(_0221_));
 sky130_fd_sc_hd__a211o_2 _0765_ (.A1(_0194_),
    .A2(_0218_),
    .B1(net48),
    .C1(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__a32oi_4 _0766_ (.A1(_0201_),
    .A2(_0212_),
    .A3(_0215_),
    .B1(_0217_),
    .B2(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__xnor2_1 _0767_ (.A(_0174_),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__inv_2 _0768_ (.A(_0209_),
    .Y(_0225_));
 sky130_fd_sc_hd__mux2_1 _0769_ (.A0(_0204_),
    .A1(_0225_),
    .S(_0211_),
    .X(_0226_));
 sky130_fd_sc_hd__a21oi_4 _0770_ (.A1(_0201_),
    .A2(_0215_),
    .B1(_0226_),
    .Y(_0227_));
 sky130_fd_sc_hd__and3_2 _0771_ (.A(_0201_),
    .B(_0215_),
    .C(_0226_),
    .X(_0228_));
 sky130_fd_sc_hd__and4b_1 _0772_ (.A_N(_0182_),
    .B(_0180_),
    .C(_0124_),
    .D(_0177_),
    .X(_0229_));
 sky130_fd_sc_hd__a21boi_1 _0773_ (.A1(_0124_),
    .A2(_0177_),
    .B1_N(_0182_),
    .Y(_0230_));
 sky130_fd_sc_hd__o21ba_1 _0774_ (.A1(_0229_),
    .A2(_0230_),
    .B1_N(_0121_),
    .X(_0231_));
 sky130_fd_sc_hd__and3_1 _0775_ (.A(_0121_),
    .B(_0124_),
    .C(_0177_),
    .X(_0232_));
 sky130_fd_sc_hd__o21a_1 _0776_ (.A1(_0206_),
    .A2(_0232_),
    .B1(_0182_),
    .X(_0233_));
 sky130_fd_sc_hd__o21ai_1 _0777_ (.A1(_0231_),
    .A2(_0233_),
    .B1(_0122_),
    .Y(_0234_));
 sky130_fd_sc_hd__a21o_1 _0778_ (.A1(_0124_),
    .A2(_0177_),
    .B1(_0182_),
    .X(_0235_));
 sky130_fd_sc_hd__nand2_1 _0779_ (.A(_0121_),
    .B(_0180_),
    .Y(_0236_));
 sky130_fd_sc_hd__a21o_1 _0780_ (.A1(_0122_),
    .A2(_0235_),
    .B1(_0236_),
    .X(_0237_));
 sky130_fd_sc_hd__nand2_1 _0781_ (.A(_0123_),
    .B(_0177_),
    .Y(_0238_));
 sky130_fd_sc_hd__nand2_1 _0782_ (.A(_0124_),
    .B(_0175_),
    .Y(_0239_));
 sky130_fd_sc_hd__xor2_2 _0783_ (.A(_0238_),
    .B(_0239_),
    .X(_0240_));
 sky130_fd_sc_hd__a21o_1 _0784_ (.A1(_0234_),
    .A2(_0237_),
    .B1(_0240_),
    .X(_0241_));
 sky130_fd_sc_hd__nand3_1 _0785_ (.A(_0240_),
    .B(_0234_),
    .C(_0237_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _0786_ (.A(_0124_),
    .B(_0177_),
    .Y(_0243_));
 sky130_fd_sc_hd__nand2_1 _0787_ (.A(_0122_),
    .B(_0180_),
    .Y(_0244_));
 sky130_fd_sc_hd__xnor2_2 _0788_ (.A(_0243_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_2 _0789_ (.A(_0171_),
    .B(_0169_),
    .Y(_0246_));
 sky130_fd_sc_hd__nand2_1 _0790_ (.A(_0245_),
    .B(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__a21bo_1 _0791_ (.A1(_0241_),
    .A2(_0242_),
    .B1_N(_0247_),
    .X(_0248_));
 sky130_fd_sc_hd__or2_1 _0792_ (.A(_0245_),
    .B(_0246_),
    .X(_0249_));
 sky130_fd_sc_hd__a21o_1 _0793_ (.A1(_0241_),
    .A2(_0242_),
    .B1(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__o31a_1 _0794_ (.A1(_0227_),
    .A2(_0228_),
    .A3(_0248_),
    .B1(_0250_),
    .X(_0251_));
 sky130_fd_sc_hd__nand3_1 _0795_ (.A(_0174_),
    .B(_0222_),
    .C(_0217_),
    .Y(_0252_));
 sky130_fd_sc_hd__a21o_1 _0796_ (.A1(_0222_),
    .A2(_0217_),
    .B1(_0174_),
    .X(_0253_));
 sky130_fd_sc_hd__a2111oi_1 _0797_ (.A1(_0252_),
    .A2(_0253_),
    .B1(_0227_),
    .C1(_0228_),
    .D1(_0246_),
    .Y(_0254_));
 sky130_fd_sc_hd__and2_1 _0798_ (.A(_0241_),
    .B(_0242_),
    .X(_0255_));
 sky130_fd_sc_hd__o311a_1 _0799_ (.A1(_0227_),
    .A2(_0228_),
    .A3(_0245_),
    .B1(_0249_),
    .C1(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__a211o_1 _0800_ (.A1(_0224_),
    .A2(_0251_),
    .B1(net36),
    .C1(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__a2111o_1 _0801_ (.A1(_0252_),
    .A2(_0253_),
    .B1(_0227_),
    .C1(_0228_),
    .D1(_0246_),
    .X(_0258_));
 sky130_fd_sc_hd__nor2_1 _0802_ (.A(_0221_),
    .B(net57),
    .Y(_0259_));
 sky130_fd_sc_hd__a311o_1 _0803_ (.A1(_0185_),
    .A2(_0196_),
    .A3(_0189_),
    .B1(_0216_),
    .C1(_0174_),
    .X(_0260_));
 sky130_fd_sc_hd__or3b_1 _0804_ (.A(_0174_),
    .B(_0191_),
    .C_N(_0218_),
    .X(_0261_));
 sky130_fd_sc_hd__a31o_1 _0805_ (.A1(_0185_),
    .A2(_0196_),
    .A3(_0189_),
    .B1(_0216_),
    .X(_0262_));
 sky130_fd_sc_hd__o21a_1 _0806_ (.A1(_0186_),
    .A2(_0191_),
    .B1(_0197_),
    .X(_0263_));
 sky130_fd_sc_hd__a22oi_2 _0807_ (.A1(_0202_),
    .A2(_0197_),
    .B1(_0211_),
    .B2(_0263_),
    .Y(_0264_));
 sky130_fd_sc_hd__o221a_1 _0808_ (.A1(_0259_),
    .A2(_0260_),
    .B1(_0261_),
    .B2(_0262_),
    .C1(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__nand4b_2 _0809_ (.A_N(_0174_),
    .B(_0201_),
    .C(_0212_),
    .D(_0215_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _0810_ (.A(_0168_),
    .B(_0172_),
    .Y(_0267_));
 sky130_fd_sc_hd__or2b_1 _0811_ (.A(_0267_),
    .B_N(_0246_),
    .X(_0268_));
 sky130_fd_sc_hd__and3_1 _0812_ (.A(_0265_),
    .B(_0266_),
    .C(_0268_),
    .X(_0269_));
 sky130_fd_sc_hd__a21oi_1 _0813_ (.A1(_0265_),
    .A2(_0266_),
    .B1(_0268_),
    .Y(_0270_));
 sky130_fd_sc_hd__inv_2 _0814_ (.A(_0177_),
    .Y(_0271_));
 sky130_fd_sc_hd__nor2_1 _0815_ (.A(_0271_),
    .B(_0206_),
    .Y(\M0.FPM0.d ));
 sky130_fd_sc_hd__nand2_1 _0816_ (.A(_0122_),
    .B(_0182_),
    .Y(_0272_));
 sky130_fd_sc_hd__xor2_1 _0817_ (.A(_0236_),
    .B(_0272_),
    .X(_0273_));
 sky130_fd_sc_hd__a32o_1 _0818_ (.A1(_0122_),
    .A2(_0124_),
    .A3(\M0.FPM0.d ),
    .B1(_0240_),
    .B2(_0273_),
    .X(_0274_));
 sky130_fd_sc_hd__or2_1 _0819_ (.A(_0240_),
    .B(_0273_),
    .X(_0275_));
 sky130_fd_sc_hd__nand2_2 _0820_ (.A(_0274_),
    .B(_0275_),
    .Y(_0276_));
 sky130_fd_sc_hd__inv_2 _0821_ (.A(_0122_),
    .Y(_0277_));
 sky130_fd_sc_hd__and2_1 _0822_ (.A(_0122_),
    .B(_0169_),
    .X(_0278_));
 sky130_fd_sc_hd__inv_2 _0823_ (.A(_0118_),
    .Y(_0279_));
 sky130_fd_sc_hd__a311o_1 _0824_ (.A1(_0121_),
    .A2(_0277_),
    .A3(_0182_),
    .B1(_0278_),
    .C1(_0279_),
    .X(_0280_));
 sky130_fd_sc_hd__or2b_1 _0825_ (.A(_0169_),
    .B_N(_0122_),
    .X(_0281_));
 sky130_fd_sc_hd__a21oi_1 _0826_ (.A1(_0279_),
    .A2(_0281_),
    .B1(_0206_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _0827_ (.A(_0121_),
    .B(_0182_),
    .Y(_0283_));
 sky130_fd_sc_hd__nand2_1 _0828_ (.A(_0122_),
    .B(_0169_),
    .Y(_0284_));
 sky130_fd_sc_hd__o21ai_1 _0829_ (.A1(_0118_),
    .A2(_0122_),
    .B1(_0180_),
    .Y(_0285_));
 sky130_fd_sc_hd__and3_1 _0830_ (.A(_0283_),
    .B(_0284_),
    .C(_0285_),
    .X(_0286_));
 sky130_fd_sc_hd__and4bb_1 _0831_ (.A_N(_0180_),
    .B_N(_0283_),
    .C(_0122_),
    .D(_0169_),
    .X(_0287_));
 sky130_fd_sc_hd__a211o_2 _0832_ (.A1(_0280_),
    .A2(_0282_),
    .B1(_0286_),
    .C1(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _0833_ (.A(_0123_),
    .B(_0175_),
    .Y(_0289_));
 sky130_fd_sc_hd__a21oi_1 _0834_ (.A1(_0119_),
    .A2(_0177_),
    .B1(_0124_),
    .Y(_0290_));
 sky130_fd_sc_hd__or2_1 _0835_ (.A(_0208_),
    .B(_0290_),
    .X(_0291_));
 sky130_fd_sc_hd__and4_1 _0836_ (.A(_0123_),
    .B(_0124_),
    .C(_0171_),
    .D(_0175_),
    .X(_0292_));
 sky130_fd_sc_hd__nor2b_1 _0837_ (.A(_0171_),
    .B_N(_0124_),
    .Y(_0293_));
 sky130_fd_sc_hd__a21bo_1 _0838_ (.A1(_0124_),
    .A2(_0171_),
    .B1_N(_0119_),
    .X(_0294_));
 sky130_fd_sc_hd__and3b_1 _0839_ (.A_N(\M0.FBM4.q ),
    .B(_0175_),
    .C(_0123_),
    .X(_0295_));
 sky130_fd_sc_hd__o221a_1 _0840_ (.A1(_0119_),
    .A2(_0293_),
    .B1(_0294_),
    .B2(_0295_),
    .C1(_0177_),
    .X(_0296_));
 sky130_fd_sc_hd__a221o_2 _0841_ (.A1(_0289_),
    .A2(_0291_),
    .B1(_0292_),
    .B2(_0271_),
    .C1(_0296_),
    .X(_0297_));
 sky130_fd_sc_hd__xnor2_2 _0842_ (.A(_0288_),
    .B(_0297_),
    .Y(_0298_));
 sky130_fd_sc_hd__xnor2_2 _0843_ (.A(_0276_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__a211o_1 _0844_ (.A1(_0258_),
    .A2(_0269_),
    .B1(_0270_),
    .C1(_0299_),
    .X(_0300_));
 sky130_fd_sc_hd__o2111a_1 _0845_ (.A1(_0174_),
    .A2(_0223_),
    .B1(_0299_),
    .C1(_0264_),
    .D1(_0268_),
    .X(_0301_));
 sky130_fd_sc_hd__xor2_1 _0846_ (.A(_0276_),
    .B(_0298_),
    .X(_0302_));
 sky130_fd_sc_hd__a211o_1 _0847_ (.A1(_0265_),
    .A2(_0266_),
    .B1(_0268_),
    .C1(_0302_),
    .X(_0303_));
 sky130_fd_sc_hd__a21bo_1 _0848_ (.A1(_0258_),
    .A2(_0301_),
    .B1_N(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__a21o_2 _0849_ (.A1(_0257_),
    .A2(_0300_),
    .B1(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__a21o_1 _0850_ (.A1(_0122_),
    .A2(_0169_),
    .B1(_0182_),
    .X(_0306_));
 sky130_fd_sc_hd__nand2_2 _0851_ (.A(_0117_),
    .B(_0180_),
    .Y(_0307_));
 sky130_fd_sc_hd__a21oi_2 _0852_ (.A1(_0118_),
    .A2(_0306_),
    .B1(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand4b_2 _0853_ (.A_N(_0182_),
    .B(_0180_),
    .C(_0122_),
    .D(_0169_),
    .Y(_0309_));
 sky130_fd_sc_hd__a21bo_1 _0854_ (.A1(_0122_),
    .A2(_0169_),
    .B1_N(_0182_),
    .X(_0310_));
 sky130_fd_sc_hd__a21oi_2 _0855_ (.A1(_0309_),
    .A2(_0310_),
    .B1(_0117_),
    .Y(_0311_));
 sky130_fd_sc_hd__and2_1 _0856_ (.A(_0117_),
    .B(_0182_),
    .X(_0312_));
 sky130_fd_sc_hd__a22o_1 _0857_ (.A1(_0182_),
    .A2(_0206_),
    .B1(_0278_),
    .B2(_0312_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _0858_ (.A(_0279_),
    .B(_0307_),
    .Y(_0314_));
 sky130_fd_sc_hd__nand2_4 _0859_ (.A(_0121_),
    .B(_0169_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_2 _0860_ (.A(_0122_),
    .B(_0172_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_4 _0861_ (.A(_0315_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__o311ai_4 _0862_ (.A1(_0308_),
    .A2(_0311_),
    .A3(_0313_),
    .B1(_0314_),
    .C1(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__a211oi_1 _0863_ (.A1(_0309_),
    .A2(_0310_),
    .B1(_0117_),
    .C1(_0279_),
    .Y(_0319_));
 sky130_fd_sc_hd__a2111o_1 _0864_ (.A1(_0118_),
    .A2(_0313_),
    .B1(_0319_),
    .C1(_0317_),
    .D1(_0308_),
    .X(_0320_));
 sky130_fd_sc_hd__a21o_1 _0865_ (.A1(_0284_),
    .A2(_0285_),
    .B1(_0283_),
    .X(_0321_));
 sky130_fd_sc_hd__a21o_2 _0866_ (.A1(_0318_),
    .A2(_0320_),
    .B1(_0321_),
    .X(_0322_));
 sky130_fd_sc_hd__nand3_2 _0867_ (.A(_0321_),
    .B(_0318_),
    .C(_0320_),
    .Y(_0323_));
 sky130_fd_sc_hd__nand2_2 _0868_ (.A(_0123_),
    .B(_0171_),
    .Y(_0324_));
 sky130_fd_sc_hd__nand2_2 _0869_ (.A(_0124_),
    .B(_0168_),
    .Y(_0325_));
 sky130_fd_sc_hd__xor2_2 _0870_ (.A(_0324_),
    .B(_0325_),
    .X(_0326_));
 sky130_fd_sc_hd__nand2_1 _0871_ (.A(_0119_),
    .B(_0177_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_2 _0872_ (.A(\M0.FBM4.q ),
    .B(_0171_),
    .Y(_0328_));
 sky130_fd_sc_hd__nor2_2 _0873_ (.A(_0327_),
    .B(_0328_),
    .Y(_0329_));
 sky130_fd_sc_hd__xnor2_2 _0874_ (.A(_0326_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__or3_1 _0875_ (.A(_0289_),
    .B(_0208_),
    .C(_0290_),
    .X(_0331_));
 sky130_fd_sc_hd__buf_2 _0876_ (.A(_0331_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_2 _0877_ (.A(\M0.FBM7.q ),
    .B(_0177_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_2 _0878_ (.A(_0119_),
    .B(_0175_),
    .Y(_0334_));
 sky130_fd_sc_hd__xor2_2 _0879_ (.A(_0333_),
    .B(_0334_),
    .X(_0335_));
 sky130_fd_sc_hd__xnor2_2 _0880_ (.A(_0332_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__xnor2_4 _0881_ (.A(_0330_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__a21o_1 _0882_ (.A1(_0322_),
    .A2(_0323_),
    .B1(_0337_),
    .X(_0338_));
 sky130_fd_sc_hd__nand3_1 _0883_ (.A(_0322_),
    .B(_0323_),
    .C(_0337_),
    .Y(_0339_));
 sky130_fd_sc_hd__nand2_1 _0884_ (.A(_0288_),
    .B(_0297_),
    .Y(_0340_));
 sky130_fd_sc_hd__a2bb2o_1 _0885_ (.A1_N(_0288_),
    .A2_N(_0297_),
    .B1(_0274_),
    .B2(_0275_),
    .X(_0341_));
 sky130_fd_sc_hd__and2_1 _0886_ (.A(_0340_),
    .B(_0341_),
    .X(_0342_));
 sky130_fd_sc_hd__a21oi_1 _0887_ (.A1(_0338_),
    .A2(_0339_),
    .B1(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__and3_1 _0888_ (.A(_0338_),
    .B(_0342_),
    .C(_0339_),
    .X(_0344_));
 sky130_fd_sc_hd__and3_1 _0889_ (.A(_0246_),
    .B(_0265_),
    .C(_0266_),
    .X(_0345_));
 sky130_fd_sc_hd__or4_4 _0890_ (.A(_0343_),
    .B(_0344_),
    .C(_0267_),
    .D(_0345_),
    .X(_0346_));
 sky130_fd_sc_hd__a21oi_1 _0891_ (.A1(_0322_),
    .A2(_0323_),
    .B1(_0337_),
    .Y(_0347_));
 sky130_fd_sc_hd__a32oi_4 _0892_ (.A1(_0322_),
    .A2(_0323_),
    .A3(_0337_),
    .B1(_0340_),
    .B2(_0341_),
    .Y(_0348_));
 sky130_fd_sc_hd__xnor2_2 _0893_ (.A(_0324_),
    .B(_0325_),
    .Y(_0349_));
 sky130_fd_sc_hd__o21ba_1 _0894_ (.A1(_0332_),
    .A2(_0349_),
    .B1_N(_0329_),
    .X(_0350_));
 sky130_fd_sc_hd__and2_1 _0895_ (.A(_0332_),
    .B(_0349_),
    .X(_0351_));
 sky130_fd_sc_hd__xnor2_2 _0896_ (.A(_0333_),
    .B(_0334_),
    .Y(_0352_));
 sky130_fd_sc_hd__and2_2 _0897_ (.A(_0119_),
    .B(_0177_),
    .X(_0353_));
 sky130_fd_sc_hd__nand2_2 _0898_ (.A(\M0.FBM7.q ),
    .B(_0175_),
    .Y(_0354_));
 sky130_fd_sc_hd__o2111ai_4 _0899_ (.A1(_0353_),
    .A2(_0354_),
    .B1(_0328_),
    .C1(_0123_),
    .D1(_0168_),
    .Y(_0355_));
 sky130_fd_sc_hd__a311o_1 _0900_ (.A1(_0123_),
    .A2(_0168_),
    .A3(_0328_),
    .B1(_0354_),
    .C1(_0353_),
    .X(_0356_));
 sky130_fd_sc_hd__and2_1 _0901_ (.A(_0355_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__o211ai_2 _0902_ (.A1(_0350_),
    .A2(_0351_),
    .B1(_0352_),
    .C1(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__a211o_1 _0903_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0332_),
    .C1(_0352_),
    .X(_0359_));
 sky130_fd_sc_hd__nand4_1 _0904_ (.A(_0332_),
    .B(_0349_),
    .C(_0355_),
    .D(_0356_),
    .Y(_0360_));
 sky130_fd_sc_hd__a21o_1 _0905_ (.A1(_0359_),
    .A2(_0360_),
    .B1(_0329_),
    .X(_0361_));
 sky130_fd_sc_hd__a21o_1 _0906_ (.A1(_0355_),
    .A2(_0356_),
    .B1(_0332_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _0907_ (.A(_0353_),
    .B(_0292_),
    .Y(_0363_));
 sky130_fd_sc_hd__a31o_1 _0908_ (.A1(_0355_),
    .A2(_0356_),
    .A3(_0363_),
    .B1(_0352_),
    .X(_0364_));
 sky130_fd_sc_hd__a21o_1 _0909_ (.A1(_0362_),
    .A2(_0364_),
    .B1(_0349_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _0910_ (.A(_0119_),
    .B(_0171_),
    .Y(_0366_));
 sky130_fd_sc_hd__a31o_1 _0911_ (.A1(_0358_),
    .A2(_0361_),
    .A3(_0365_),
    .B1(_0366_),
    .X(_0367_));
 sky130_fd_sc_hd__nand4_2 _0912_ (.A(_0366_),
    .B(_0358_),
    .C(_0361_),
    .D(_0365_),
    .Y(_0368_));
 sky130_fd_sc_hd__o211a_1 _0913_ (.A1(_0347_),
    .A2(_0348_),
    .B1(_0367_),
    .C1(_0368_),
    .X(_0369_));
 sky130_fd_sc_hd__nand2_1 _0914_ (.A(_0118_),
    .B(_0169_),
    .Y(_0370_));
 sky130_fd_sc_hd__nand2_2 _0915_ (.A(_0118_),
    .B(_0182_),
    .Y(_0371_));
 sky130_fd_sc_hd__xor2_4 _0916_ (.A(_0307_),
    .B(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__and4_2 _0917_ (.A(_0118_),
    .B(_0122_),
    .C(_0169_),
    .D(_0180_),
    .X(_0373_));
 sky130_fd_sc_hd__nand2_1 _0918_ (.A(_0121_),
    .B(_0172_),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_1 _0919_ (.A(_0118_),
    .B(_0180_),
    .Y(_0375_));
 sky130_fd_sc_hd__o211a_1 _0920_ (.A1(_0278_),
    .A2(_0374_),
    .B1(_0312_),
    .C1(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__and2_1 _0921_ (.A(_0118_),
    .B(_0180_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _0922_ (.A(_0117_),
    .B(_0182_),
    .Y(_0378_));
 sky130_fd_sc_hd__and2_1 _0923_ (.A(_0121_),
    .B(_0172_),
    .X(_0379_));
 sky130_fd_sc_hd__o211a_1 _0924_ (.A1(_0377_),
    .A2(_0378_),
    .B1(_0379_),
    .C1(_0284_),
    .X(_0380_));
 sky130_fd_sc_hd__a211o_1 _0925_ (.A1(_0372_),
    .A2(_0373_),
    .B1(_0376_),
    .C1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__xor2_2 _0926_ (.A(_0315_),
    .B(_0316_),
    .X(_0382_));
 sky130_fd_sc_hd__a211o_1 _0927_ (.A1(_0284_),
    .A2(_0379_),
    .B1(_0378_),
    .C1(_0377_),
    .X(_0383_));
 sky130_fd_sc_hd__a211o_1 _0928_ (.A1(_0375_),
    .A2(_0312_),
    .B1(_0374_),
    .C1(_0278_),
    .X(_0384_));
 sky130_fd_sc_hd__o2111a_1 _0929_ (.A1(_0372_),
    .A2(_0373_),
    .B1(_0382_),
    .C1(_0383_),
    .D1(_0384_),
    .X(_0385_));
 sky130_fd_sc_hd__a211oi_1 _0930_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0372_),
    .C1(_0373_),
    .Y(_0386_));
 sky130_fd_sc_hd__a211o_1 _0931_ (.A1(_0317_),
    .A2(_0381_),
    .B1(_0385_),
    .C1(_0386_),
    .X(_0387_));
 sky130_fd_sc_hd__xnor2_1 _0932_ (.A(_0370_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__xnor2_1 _0933_ (.A(_0322_),
    .B(_0388_),
    .Y(_0389_));
 sky130_fd_sc_hd__a211oi_2 _0934_ (.A1(_0367_),
    .A2(_0368_),
    .B1(_0347_),
    .C1(_0348_),
    .Y(_0390_));
 sky130_fd_sc_hd__or3_1 _0935_ (.A(_0369_),
    .B(_0389_),
    .C(_0390_),
    .X(_0391_));
 sky130_fd_sc_hd__o21ai_1 _0936_ (.A1(_0369_),
    .A2(_0390_),
    .B1(_0389_),
    .Y(_0392_));
 sky130_fd_sc_hd__and2_2 _0937_ (.A(_0391_),
    .B(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _0938_ (.A(_0121_),
    .B(_0124_),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2_1 _0939_ (.A(_0122_),
    .B(_0123_),
    .Y(_0395_));
 sky130_fd_sc_hd__xnor2_2 _0940_ (.A(_0394_),
    .B(_0395_),
    .Y(_0396_));
 sky130_fd_sc_hd__o22a_2 _0941_ (.A1(_0343_),
    .A2(_0344_),
    .B1(_0267_),
    .B2(_0345_),
    .X(_0397_));
 sky130_fd_sc_hd__a2111o_1 _0942_ (.A1(_0305_),
    .A2(_0346_),
    .B1(_0393_),
    .C1(_0396_),
    .D1(_0397_),
    .X(_0398_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(_0138_),
    .B(_0396_),
    .X(_0399_));
 sky130_fd_sc_hd__a211o_1 _0944_ (.A1(_0305_),
    .A2(_0346_),
    .B1(_0399_),
    .C1(_0397_),
    .X(_0400_));
 sky130_fd_sc_hd__o21bai_2 _0945_ (.A1(_0389_),
    .A2(_0390_),
    .B1_N(_0369_),
    .Y(_0401_));
 sky130_fd_sc_hd__o311a_1 _0946_ (.A1(_0308_),
    .A2(_0311_),
    .A3(_0313_),
    .B1(_0314_),
    .C1(_0317_),
    .X(_0402_));
 sky130_fd_sc_hd__nor3_1 _0947_ (.A(_0317_),
    .B(_0372_),
    .C(_0373_),
    .Y(_0403_));
 sky130_fd_sc_hd__a21oi_1 _0948_ (.A1(_0383_),
    .A2(_0384_),
    .B1(_0321_),
    .Y(_0404_));
 sky130_fd_sc_hd__o21ai_1 _0949_ (.A1(_0402_),
    .A2(_0403_),
    .B1(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__a21oi_1 _0950_ (.A1(_0318_),
    .A2(_0320_),
    .B1(_0321_),
    .Y(_0406_));
 sky130_fd_sc_hd__o2bb2a_1 _0951_ (.A1_N(_0370_),
    .A2_N(_0405_),
    .B1(_0387_),
    .B2(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__nand2_1 _0952_ (.A(_0117_),
    .B(_0169_),
    .Y(_0408_));
 sky130_fd_sc_hd__nand2_1 _0953_ (.A(_0118_),
    .B(_0172_),
    .Y(_0409_));
 sky130_fd_sc_hd__xor2_2 _0954_ (.A(_0408_),
    .B(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__inv_2 _0955_ (.A(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__a211o_1 _0956_ (.A1(_0382_),
    .A2(_0372_),
    .B1(_0312_),
    .C1(_0278_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _0957_ (.A(_0377_),
    .B(_0378_),
    .Y(_0413_));
 sky130_fd_sc_hd__or3b_1 _0958_ (.A(_0378_),
    .B(_0374_),
    .C_N(_0373_),
    .X(_0414_));
 sky130_fd_sc_hd__a21o_1 _0959_ (.A1(_0377_),
    .A2(_0312_),
    .B1(_0379_),
    .X(_0415_));
 sky130_fd_sc_hd__a32o_1 _0960_ (.A1(_0382_),
    .A2(_0413_),
    .A3(_0372_),
    .B1(_0414_),
    .B2(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__and2_1 _0961_ (.A(_0412_),
    .B(_0416_),
    .X(_0417_));
 sky130_fd_sc_hd__clkbuf_2 _0962_ (.A(_0417_),
    .X(_0418_));
 sky130_fd_sc_hd__xnor2_1 _0963_ (.A(_0411_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__xnor2_1 _0964_ (.A(_0407_),
    .B(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__or3_1 _0965_ (.A(_0349_),
    .B(_0352_),
    .C(_0357_),
    .X(_0421_));
 sky130_fd_sc_hd__or4bb_1 _0966_ (.A(_0326_),
    .B(_0329_),
    .C_N(_0357_),
    .D_N(_0332_),
    .X(_0422_));
 sky130_fd_sc_hd__nor2_1 _0967_ (.A(_0326_),
    .B(_0335_),
    .Y(_0423_));
 sky130_fd_sc_hd__o21ai_1 _0968_ (.A1(_0362_),
    .A2(_0423_),
    .B1(_0366_),
    .Y(_0424_));
 sky130_fd_sc_hd__and4_1 _0969_ (.A(_0358_),
    .B(_0421_),
    .C(_0422_),
    .D(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__nand2_1 _0970_ (.A(\M0.FBM7.q ),
    .B(_0171_),
    .Y(_0426_));
 sky130_fd_sc_hd__nand2_1 _0971_ (.A(_0119_),
    .B(_0168_),
    .Y(_0427_));
 sky130_fd_sc_hd__xor2_1 _0972_ (.A(_0426_),
    .B(_0427_),
    .X(_0428_));
 sky130_fd_sc_hd__nand2_1 _0973_ (.A(_0328_),
    .B(_0354_),
    .Y(_0429_));
 sky130_fd_sc_hd__nand2_1 _0974_ (.A(_0123_),
    .B(_0168_),
    .Y(_0430_));
 sky130_fd_sc_hd__or4_1 _0975_ (.A(_0327_),
    .B(_0328_),
    .C(_0354_),
    .D(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__o21ai_1 _0976_ (.A1(_0327_),
    .A2(_0354_),
    .B1(_0430_),
    .Y(_0432_));
 sky130_fd_sc_hd__inv_2 _0977_ (.A(_0168_),
    .Y(_0433_));
 sky130_fd_sc_hd__or2b_1 _0978_ (.A(_0123_),
    .B_N(_0124_),
    .X(_0434_));
 sky130_fd_sc_hd__xnor2_1 _0979_ (.A(_0124_),
    .B(_0171_),
    .Y(_0435_));
 sky130_fd_sc_hd__inv_2 _0980_ (.A(_0123_),
    .Y(_0436_));
 sky130_fd_sc_hd__o32a_1 _0981_ (.A1(_0353_),
    .A2(_0354_),
    .A3(_0434_),
    .B1(_0435_),
    .B2(_0436_),
    .X(_0437_));
 sky130_fd_sc_hd__or4_1 _0982_ (.A(_0168_),
    .B(_0353_),
    .C(_0324_),
    .D(_0354_),
    .X(_0438_));
 sky130_fd_sc_hd__o21ai_1 _0983_ (.A1(_0433_),
    .A2(_0437_),
    .B1(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__a32o_1 _0984_ (.A1(_0429_),
    .A2(_0431_),
    .A3(_0432_),
    .B1(_0439_),
    .B2(_0335_),
    .X(_0440_));
 sky130_fd_sc_hd__xor2_1 _0985_ (.A(_0428_),
    .B(_0440_),
    .X(_0441_));
 sky130_fd_sc_hd__xnor2_1 _0986_ (.A(_0425_),
    .B(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__xnor2_1 _0987_ (.A(_0420_),
    .B(_0442_),
    .Y(_0443_));
 sky130_fd_sc_hd__xnor2_2 _0988_ (.A(_0401_),
    .B(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__o21a_1 _0989_ (.A1(_0393_),
    .A2(_0399_),
    .B1(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__a31o_1 _0990_ (.A1(_0397_),
    .A2(_0391_),
    .A3(_0392_),
    .B1(_0138_),
    .X(_0446_));
 sky130_fd_sc_hd__a31o_1 _0991_ (.A1(_0305_),
    .A2(_0346_),
    .A3(_0393_),
    .B1(_0446_),
    .X(_0447_));
 sky130_fd_sc_hd__a32o_1 _0992_ (.A1(_0398_),
    .A2(_0400_),
    .A3(_0445_),
    .B1(_0447_),
    .B2(_0396_),
    .X(_0448_));
 sky130_fd_sc_hd__a2111o_2 _0993_ (.A1(_0305_),
    .A2(_0346_),
    .B1(_0393_),
    .C1(_0397_),
    .D1(_0444_),
    .X(_0449_));
 sky130_fd_sc_hd__o21ai_1 _0994_ (.A1(_0122_),
    .A2(_0129_),
    .B1(_0130_),
    .Y(_0450_));
 sky130_fd_sc_hd__nor2_1 _0995_ (.A(_0118_),
    .B(_0119_),
    .Y(_0451_));
 sky130_fd_sc_hd__a22o_1 _0996_ (.A1(_0118_),
    .A2(_0450_),
    .B1(_0451_),
    .B2(_0122_),
    .X(_0452_));
 sky130_fd_sc_hd__nor2_1 _0997_ (.A(_0124_),
    .B(_0130_),
    .Y(_0453_));
 sky130_fd_sc_hd__a2bb2o_1 _0998_ (.A1_N(_0119_),
    .A2_N(_0124_),
    .B1(_0131_),
    .B2(_0277_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(_0453_),
    .A1(_0454_),
    .S(_0129_),
    .X(_0455_));
 sky130_fd_sc_hd__a21oi_2 _1000_ (.A1(_0124_),
    .A2(_0452_),
    .B1(_0455_),
    .Y(_0456_));
 sky130_fd_sc_hd__inv_2 _1001_ (.A(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__a21o_1 _1002_ (.A1(_0448_),
    .A2(_0449_),
    .B1(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__and2_1 _1003_ (.A(_0134_),
    .B(_0146_),
    .X(_0459_));
 sky130_fd_sc_hd__or2_1 _1004_ (.A(_0420_),
    .B(_0442_),
    .X(_0460_));
 sky130_fd_sc_hd__and2_1 _1005_ (.A(_0420_),
    .B(_0442_),
    .X(_0461_));
 sky130_fd_sc_hd__a21o_2 _1006_ (.A1(_0401_),
    .A2(_0460_),
    .B1(_0461_),
    .X(_0462_));
 sky130_fd_sc_hd__and2_1 _1007_ (.A(_0428_),
    .B(_0440_),
    .X(_0463_));
 sky130_fd_sc_hd__a41o_1 _1008_ (.A1(_0123_),
    .A2(_0124_),
    .A3(_0175_),
    .A4(_0177_),
    .B1(_0366_),
    .X(_0464_));
 sky130_fd_sc_hd__nand3_1 _1009_ (.A(\M0.FBM7.q ),
    .B(_0168_),
    .C(_0464_),
    .Y(_0465_));
 sky130_fd_sc_hd__or2_1 _1010_ (.A(_0428_),
    .B(_0440_),
    .X(_0466_));
 sky130_fd_sc_hd__o211a_1 _1011_ (.A1(_0425_),
    .A2(_0463_),
    .B1(_0465_),
    .C1(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__o21ba_2 _1012_ (.A1(_0463_),
    .A2(_0465_),
    .B1_N(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__nand2_1 _1013_ (.A(_0117_),
    .B(_0172_),
    .Y(_0469_));
 sky130_fd_sc_hd__or2b_1 _1014_ (.A(_0469_),
    .B_N(_0370_),
    .X(_0470_));
 sky130_fd_sc_hd__nand2_1 _1015_ (.A(_0414_),
    .B(_0470_),
    .Y(_0471_));
 sky130_fd_sc_hd__a211o_1 _1016_ (.A1(_0410_),
    .A2(_0418_),
    .B1(_0406_),
    .C1(_0387_),
    .X(_0472_));
 sky130_fd_sc_hd__o21a_1 _1017_ (.A1(_0410_),
    .A2(_0418_),
    .B1(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__nand2_1 _1018_ (.A(_0402_),
    .B(_0404_),
    .Y(_0474_));
 sky130_fd_sc_hd__and4b_1 _1019_ (.A_N(_0321_),
    .B(_0382_),
    .C(_0372_),
    .D(_0373_),
    .X(_0475_));
 sky130_fd_sc_hd__a21oi_1 _1020_ (.A1(_0403_),
    .A2(_0404_),
    .B1(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__and3_1 _1021_ (.A(_0469_),
    .B(_0474_),
    .C(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__a31oi_1 _1022_ (.A1(_0411_),
    .A2(_0474_),
    .A3(_0476_),
    .B1(_0469_),
    .Y(_0478_));
 sky130_fd_sc_hd__mux2_1 _1023_ (.A0(_0477_),
    .A1(_0478_),
    .S(_0418_),
    .X(_0479_));
 sky130_fd_sc_hd__a2bb2o_2 _1024_ (.A1_N(_0471_),
    .A2_N(_0473_),
    .B1(_0479_),
    .B2(_0370_),
    .X(_0480_));
 sky130_fd_sc_hd__xor2_1 _1025_ (.A(_0468_),
    .B(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__xnor2_2 _1026_ (.A(_0462_),
    .B(_0481_),
    .Y(_0482_));
 sky130_fd_sc_hd__o21ba_1 _1027_ (.A1(_0147_),
    .A2(_0459_),
    .B1_N(_0482_),
    .X(_0483_));
 sky130_fd_sc_hd__or2_1 _1028_ (.A(_0147_),
    .B(_0459_),
    .X(_0484_));
 sky130_fd_sc_hd__and3_1 _1029_ (.A(_0457_),
    .B(_0448_),
    .C(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__and2_1 _1030_ (.A(_0468_),
    .B(_0480_),
    .X(_0486_));
 sky130_fd_sc_hd__o21a_1 _1031_ (.A1(_0119_),
    .A2(_0440_),
    .B1(_0171_),
    .X(_0487_));
 sky130_fd_sc_hd__a21o_1 _1032_ (.A1(_0119_),
    .A2(_0440_),
    .B1(_0487_),
    .X(_0488_));
 sky130_fd_sc_hd__and3_2 _1033_ (.A(\M0.FBM7.q ),
    .B(_0168_),
    .C(_0488_),
    .X(_0489_));
 sky130_fd_sc_hd__nand2_1 _1034_ (.A(_0474_),
    .B(_0476_),
    .Y(_0490_));
 sky130_fd_sc_hd__o31a_1 _1035_ (.A1(_0169_),
    .A2(_0418_),
    .A3(_0490_),
    .B1(_0118_),
    .X(_0491_));
 sky130_fd_sc_hd__o21a_1 _1036_ (.A1(_0418_),
    .A2(_0490_),
    .B1(_0169_),
    .X(_0492_));
 sky130_fd_sc_hd__o21ba_1 _1037_ (.A1(_0491_),
    .A2(_0492_),
    .B1_N(_0469_),
    .X(_0493_));
 sky130_fd_sc_hd__xnor2_2 _1038_ (.A(_0489_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__a211oi_1 _1039_ (.A1(_0468_),
    .A2(_0480_),
    .B1(_0494_),
    .C1(_0462_),
    .Y(_0495_));
 sky130_fd_sc_hd__o211a_1 _1040_ (.A1(_0468_),
    .A2(_0480_),
    .B1(_0494_),
    .C1(_0462_),
    .X(_0496_));
 sky130_fd_sc_hd__nor3_1 _1041_ (.A(_0468_),
    .B(_0480_),
    .C(_0494_),
    .Y(_0497_));
 sky130_fd_sc_hd__a2111o_1 _1042_ (.A1(_0486_),
    .A2(_0494_),
    .B1(_0495_),
    .C1(_0496_),
    .D1(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__nor3b_1 _1043_ (.A(_0449_),
    .B(_0498_),
    .C_N(_0482_),
    .Y(_0499_));
 sky130_fd_sc_hd__a211oi_2 _1044_ (.A1(_0458_),
    .A2(_0483_),
    .B1(_0485_),
    .C1(_0499_),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _1045_ (.A(_0456_),
    .B(_0482_),
    .Y(_0501_));
 sky130_fd_sc_hd__nor2_1 _1046_ (.A(_0456_),
    .B(_0482_),
    .Y(_0502_));
 sky130_fd_sc_hd__a31o_1 _1047_ (.A1(_0448_),
    .A2(_0449_),
    .A3(_0501_),
    .B1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__o21ai_1 _1048_ (.A1(_0484_),
    .A2(_0503_),
    .B1(_0498_),
    .Y(_0504_));
 sky130_fd_sc_hd__nand2_1 _1049_ (.A(_0500_),
    .B(_0504_),
    .Y(_0505_));
 sky130_fd_sc_hd__xor2_2 _1050_ (.A(_0147_),
    .B(_0152_),
    .X(_0506_));
 sky130_fd_sc_hd__nand2_1 _1051_ (.A(_0120_),
    .B(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__or2_1 _1052_ (.A(_0120_),
    .B(_0506_),
    .X(_0508_));
 sky130_fd_sc_hd__and2_1 _1053_ (.A(_0507_),
    .B(_0508_),
    .X(_0509_));
 sky130_fd_sc_hd__nand2b_1 _1054_ (.A_N(_0449_),
    .B(_0482_),
    .Y(_0510_));
 sky130_fd_sc_hd__nand2_1 _1055_ (.A(_0489_),
    .B(_0493_),
    .Y(_0511_));
 sky130_fd_sc_hd__nor2_1 _1056_ (.A(_0489_),
    .B(_0493_),
    .Y(_0512_));
 sky130_fd_sc_hd__o211a_1 _1057_ (.A1(_0468_),
    .A2(_0480_),
    .B1(_0511_),
    .C1(_0462_),
    .X(_0513_));
 sky130_fd_sc_hd__a211o_1 _1058_ (.A1(_0486_),
    .A2(_0511_),
    .B1(_0512_),
    .C1(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__o211a_1 _1059_ (.A1(_0462_),
    .A2(_0480_),
    .B1(_0512_),
    .C1(_0468_),
    .X(_0515_));
 sky130_fd_sc_hd__a31o_1 _1060_ (.A1(_0462_),
    .A2(_0480_),
    .A3(_0512_),
    .B1(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__a21oi_4 _1061_ (.A1(_0510_),
    .A2(_0514_),
    .B1(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_1 _1062_ (.A(_0509_),
    .B(_0517_),
    .Y(_0518_));
 sky130_fd_sc_hd__nand2_1 _1063_ (.A(_0507_),
    .B(_0157_),
    .Y(_0519_));
 sky130_fd_sc_hd__and2_1 _1064_ (.A(_0160_),
    .B(_0165_),
    .X(_0520_));
 sky130_fd_sc_hd__a21oi_1 _1065_ (.A1(_0157_),
    .A2(_0520_),
    .B1(_0166_),
    .Y(_0521_));
 sky130_fd_sc_hd__o22a_1 _1066_ (.A1(_0519_),
    .A2(_0520_),
    .B1(_0521_),
    .B2(_0507_),
    .X(_0522_));
 sky130_fd_sc_hd__nor2_1 _1067_ (.A(_0509_),
    .B(_0517_),
    .Y(_0523_));
 sky130_fd_sc_hd__a211o_1 _1068_ (.A1(_0505_),
    .A2(_0518_),
    .B1(_0522_),
    .C1(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__nand3b_1 _1069_ (.A_N(_0155_),
    .B(_0167_),
    .C(_0524_),
    .Y(\M0.FPM15.d ));
 sky130_fd_sc_hd__a21oi_1 _1070_ (.A1(_0505_),
    .A2(_0518_),
    .B1(_0523_),
    .Y(_0525_));
 sky130_fd_sc_hd__or2_1 _1071_ (.A(_0506_),
    .B(_0517_),
    .X(_0526_));
 sky130_fd_sc_hd__a22o_1 _1072_ (.A1(_0500_),
    .A2(_0504_),
    .B1(_0508_),
    .B2(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a311o_1 _1073_ (.A1(_0500_),
    .A2(_0504_),
    .A3(_0506_),
    .B1(_0517_),
    .C1(_0120_),
    .X(_0528_));
 sky130_fd_sc_hd__xor2_2 _1074_ (.A(_0158_),
    .B(_0159_),
    .X(_0529_));
 sky130_fd_sc_hd__a211o_1 _1075_ (.A1(_0527_),
    .A2(_0528_),
    .B1(_0529_),
    .C1(_0157_),
    .X(_0530_));
 sky130_fd_sc_hd__a21oi_1 _1076_ (.A1(_0529_),
    .A2(_0526_),
    .B1(_0120_),
    .Y(_0531_));
 sky130_fd_sc_hd__a21oi_1 _1077_ (.A1(_0506_),
    .A2(_0517_),
    .B1(_0529_),
    .Y(_0532_));
 sky130_fd_sc_hd__and3_1 _1078_ (.A(_0508_),
    .B(_0517_),
    .C(_0529_),
    .X(_0533_));
 sky130_fd_sc_hd__or2_1 _1079_ (.A(_0507_),
    .B(_0160_),
    .X(_0534_));
 sky130_fd_sc_hd__and4bb_1 _1080_ (.A_N(_0533_),
    .B_N(_0157_),
    .C(_0165_),
    .D(_0534_),
    .X(_0535_));
 sky130_fd_sc_hd__o31ai_1 _1081_ (.A1(_0505_),
    .A2(_0531_),
    .A3(_0532_),
    .B1(_0535_),
    .Y(_0536_));
 sky130_fd_sc_hd__o2111a_1 _1082_ (.A1(_0525_),
    .A2(_0167_),
    .B1(_0530_),
    .C1(_0536_),
    .D1(_0524_),
    .X(\M0.FPM14.d ));
 sky130_fd_sc_hd__nand2_1 _1083_ (.A(_0507_),
    .B(_0160_),
    .Y(_0537_));
 sky130_fd_sc_hd__nand2_1 _1084_ (.A(_0534_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__xnor2_1 _1085_ (.A(_0165_),
    .B(_0538_),
    .Y(_0539_));
 sky130_fd_sc_hd__xnor2_1 _1086_ (.A(_0525_),
    .B(_0539_),
    .Y(\M0.FPM13.d ));
 sky130_fd_sc_hd__xor2_1 _1087_ (.A(_0509_),
    .B(_0517_),
    .X(_0540_));
 sky130_fd_sc_hd__xnor2_1 _1088_ (.A(_0505_),
    .B(_0540_),
    .Y(\M0.FPM12.d ));
 sky130_fd_sc_hd__xor2_1 _1089_ (.A(_0484_),
    .B(_0498_),
    .X(_0541_));
 sky130_fd_sc_hd__xnor2_1 _1090_ (.A(_0503_),
    .B(_0541_),
    .Y(\M0.FPM11.d ));
 sky130_fd_sc_hd__nand2_1 _1091_ (.A(_0448_),
    .B(_0449_),
    .Y(_0542_));
 sky130_fd_sc_hd__or2_1 _1092_ (.A(_0456_),
    .B(_0482_),
    .X(_0543_));
 sky130_fd_sc_hd__nand2_1 _1093_ (.A(_0501_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__xnor2_1 _1094_ (.A(_0542_),
    .B(_0544_),
    .Y(\M0.FPM10.d ));
 sky130_fd_sc_hd__a21oi_1 _1095_ (.A1(_0305_),
    .A2(_0346_),
    .B1(_0397_),
    .Y(_0545_));
 sky130_fd_sc_hd__or2b_1 _1096_ (.A(_0393_),
    .B_N(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__xor2_1 _1097_ (.A(_0444_),
    .B(_0396_),
    .X(_0547_));
 sky130_fd_sc_hd__a21oi_1 _1098_ (.A1(_0546_),
    .A2(_0447_),
    .B1(_0547_),
    .Y(_0548_));
 sky130_fd_sc_hd__and3_1 _1099_ (.A(_0546_),
    .B(_0447_),
    .C(_0547_),
    .X(_0549_));
 sky130_fd_sc_hd__or2_1 _1100_ (.A(_0548_),
    .B(_0549_),
    .X(_0550_));
 sky130_fd_sc_hd__clkbuf_1 _1101_ (.A(_0550_),
    .X(\M0.FPM9.d ));
 sky130_fd_sc_hd__nor2_1 _1102_ (.A(_0227_),
    .B(_0228_),
    .Y(_0551_));
 sky130_fd_sc_hd__nand2_1 _1103_ (.A(_0247_),
    .B(_0249_),
    .Y(_0552_));
 sky130_fd_sc_hd__xnor2_1 _1104_ (.A(_0551_),
    .B(_0552_),
    .Y(\M0.FPM4.d ));
 sky130_fd_sc_hd__xnor2_1 _1105_ (.A(_0138_),
    .B(_0393_),
    .Y(_0553_));
 sky130_fd_sc_hd__xnor2_1 _1106_ (.A(_0545_),
    .B(_0553_),
    .Y(\M0.FPM8.d ));
 sky130_fd_sc_hd__inv_2 _1107_ (.A(_0171_),
    .Y(_0554_));
 sky130_fd_sc_hd__mux2_1 _1108_ (.A0(_0554_),
    .A1(_0169_),
    .S(_0206_),
    .X(_0555_));
 sky130_fd_sc_hd__and3_1 _1109_ (.A(_0169_),
    .B(_0191_),
    .C(_0207_),
    .X(_0556_));
 sky130_fd_sc_hd__a21o_1 _1110_ (.A1(_0203_),
    .A2(_0555_),
    .B1(_0556_),
    .X(_0557_));
 sky130_fd_sc_hd__a32o_1 _1111_ (.A1(_0196_),
    .A2(_0191_),
    .A3(_0203_),
    .B1(_0557_),
    .B2(_0177_),
    .X(_0558_));
 sky130_fd_sc_hd__xor2_1 _1112_ (.A(_0211_),
    .B(_0558_),
    .X(\M0.FPM3.d ));
 sky130_fd_sc_hd__nand2_1 _1113_ (.A(_0175_),
    .B(_0180_),
    .Y(_0559_));
 sky130_fd_sc_hd__nand2_1 _1114_ (.A(_0177_),
    .B(_0182_),
    .Y(_0560_));
 sky130_fd_sc_hd__xor2_1 _1115_ (.A(_0559_),
    .B(_0560_),
    .X(\M0.FPM1.d ));
 sky130_fd_sc_hd__a21oi_1 _1116_ (.A1(_0271_),
    .A2(_0203_),
    .B1(_0186_),
    .Y(_0561_));
 sky130_fd_sc_hd__or3_1 _1117_ (.A(_0171_),
    .B(_0271_),
    .C(_0169_),
    .X(_0562_));
 sky130_fd_sc_hd__o21a_1 _1118_ (.A1(_0554_),
    .A2(_0561_),
    .B1(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__o221a_1 _1119_ (.A1(_0169_),
    .A2(_0180_),
    .B1(_0191_),
    .B2(_0177_),
    .C1(_0207_),
    .X(_0564_));
 sky130_fd_sc_hd__inv_2 _1120_ (.A(_0169_),
    .Y(_0565_));
 sky130_fd_sc_hd__o31a_1 _1121_ (.A1(_0271_),
    .A2(_0565_),
    .A3(_0180_),
    .B1(_0203_),
    .X(_0566_));
 sky130_fd_sc_hd__o22a_1 _1122_ (.A1(_0206_),
    .A2(_0563_),
    .B1(_0564_),
    .B2(_0566_),
    .X(\M0.FPM2.d ));
 sky130_fd_sc_hd__and2b_1 _1123_ (.A_N(_0397_),
    .B(_0346_),
    .X(_0567_));
 sky130_fd_sc_hd__xnor2_1 _1124_ (.A(_0305_),
    .B(_0567_),
    .Y(\M0.FPM7.d ));
 sky130_fd_sc_hd__a21o_1 _1125_ (.A1(_0258_),
    .A2(_0269_),
    .B1(_0270_),
    .X(_0568_));
 sky130_fd_sc_hd__xnor2_1 _1126_ (.A(_0299_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__xor2_1 _1127_ (.A(_0257_),
    .B(_0569_),
    .X(\M0.FPM6.d ));
 sky130_fd_sc_hd__or2_1 _1128_ (.A(_0227_),
    .B(_0228_),
    .X(_0570_));
 sky130_fd_sc_hd__a21o_1 _1129_ (.A1(_0570_),
    .A2(_0245_),
    .B1(_0246_),
    .X(_0571_));
 sky130_fd_sc_hd__o21ai_1 _1130_ (.A1(_0570_),
    .A2(_0245_),
    .B1(_0571_),
    .Y(_0572_));
 sky130_fd_sc_hd__xnor2_1 _1131_ (.A(_0224_),
    .B(_0255_),
    .Y(_0573_));
 sky130_fd_sc_hd__xnor2_1 _1132_ (.A(_0572_),
    .B(_0573_),
    .Y(\M0.FPM5.d ));
 sky130_fd_sc_hd__buf_8 _1133_ (.A(net19),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_16 _1134_ (.A(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__inv_2 _1135_ (.A(_0575_),
    .Y(_0000_));
 sky130_fd_sc_hd__inv_2 _1136_ (.A(_0575_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _1137_ (.A(_0575_),
    .Y(_0002_));
 sky130_fd_sc_hd__inv_2 _1138_ (.A(_0575_),
    .Y(_0003_));
 sky130_fd_sc_hd__inv_2 _1139_ (.A(_0575_),
    .Y(_0004_));
 sky130_fd_sc_hd__inv_2 _1140_ (.A(_0575_),
    .Y(_0005_));
 sky130_fd_sc_hd__inv_2 _1141_ (.A(_0575_),
    .Y(_0006_));
 sky130_fd_sc_hd__inv_2 _1142_ (.A(_0575_),
    .Y(_0007_));
 sky130_fd_sc_hd__inv_2 _1143_ (.A(_0575_),
    .Y(_0008_));
 sky130_fd_sc_hd__inv_2 _1144_ (.A(_0575_),
    .Y(_0009_));
 sky130_fd_sc_hd__inv_2 _1145_ (.A(_0575_),
    .Y(_0010_));
 sky130_fd_sc_hd__inv_2 _1146_ (.A(_0575_),
    .Y(_0011_));
 sky130_fd_sc_hd__inv_2 _1147_ (.A(_0575_),
    .Y(_0012_));
 sky130_fd_sc_hd__inv_2 _1148_ (.A(_0575_),
    .Y(_0013_));
 sky130_fd_sc_hd__inv_2 _1149_ (.A(_0575_),
    .Y(_0014_));
 sky130_fd_sc_hd__inv_2 _1150_ (.A(_0575_),
    .Y(_0015_));
 sky130_fd_sc_hd__inv_2 _1151_ (.A(_0575_),
    .Y(_0016_));
 sky130_fd_sc_hd__inv_2 _1152_ (.A(_0575_),
    .Y(_0017_));
 sky130_fd_sc_hd__inv_2 _1153_ (.A(_0575_),
    .Y(_0018_));
 sky130_fd_sc_hd__clkbuf_16 _1154_ (.A(_0574_),
    .X(_0576_));
 sky130_fd_sc_hd__inv_2 _1155_ (.A(_0576_),
    .Y(_0019_));
 sky130_fd_sc_hd__inv_2 _1156_ (.A(_0576_),
    .Y(_0020_));
 sky130_fd_sc_hd__inv_2 _1157_ (.A(_0576_),
    .Y(_0021_));
 sky130_fd_sc_hd__inv_2 _1158_ (.A(_0576_),
    .Y(_0022_));
 sky130_fd_sc_hd__inv_2 _1159_ (.A(_0576_),
    .Y(_0023_));
 sky130_fd_sc_hd__inv_2 _1160_ (.A(_0576_),
    .Y(_0024_));
 sky130_fd_sc_hd__inv_2 _1161_ (.A(_0576_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _1162_ (.A(_0576_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _1163_ (.A(_0576_),
    .Y(_0027_));
 sky130_fd_sc_hd__inv_2 _1164_ (.A(_0576_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _1165_ (.A(_0576_),
    .Y(_0029_));
 sky130_fd_sc_hd__inv_2 _1166_ (.A(_0576_),
    .Y(_0030_));
 sky130_fd_sc_hd__inv_2 _1167_ (.A(_0576_),
    .Y(_0031_));
 sky130_fd_sc_hd__inv_2 _1168_ (.A(_0576_),
    .Y(_0032_));
 sky130_fd_sc_hd__inv_2 _1169_ (.A(_0576_),
    .Y(_0033_));
 sky130_fd_sc_hd__inv_2 _1170_ (.A(_0576_),
    .Y(_0034_));
 sky130_fd_sc_hd__inv_2 _1171_ (.A(_0576_),
    .Y(_0035_));
 sky130_fd_sc_hd__inv_2 _1172_ (.A(_0576_),
    .Y(_0036_));
 sky130_fd_sc_hd__inv_2 _1173_ (.A(_0576_),
    .Y(_0037_));
 sky130_fd_sc_hd__clkbuf_16 _1174_ (.A(_0574_),
    .X(_0577_));
 sky130_fd_sc_hd__inv_2 _1175_ (.A(_0577_),
    .Y(_0038_));
 sky130_fd_sc_hd__inv_2 _1176_ (.A(_0577_),
    .Y(_0039_));
 sky130_fd_sc_hd__inv_2 _1177_ (.A(_0577_),
    .Y(_0040_));
 sky130_fd_sc_hd__inv_2 _1178_ (.A(_0577_),
    .Y(_0041_));
 sky130_fd_sc_hd__inv_2 _1179_ (.A(_0577_),
    .Y(_0042_));
 sky130_fd_sc_hd__inv_2 _1180_ (.A(_0577_),
    .Y(_0043_));
 sky130_fd_sc_hd__inv_2 _1181_ (.A(_0577_),
    .Y(_0044_));
 sky130_fd_sc_hd__inv_2 _1182_ (.A(_0577_),
    .Y(_0045_));
 sky130_fd_sc_hd__inv_2 _1183_ (.A(_0577_),
    .Y(_0046_));
 sky130_fd_sc_hd__inv_2 _1184_ (.A(_0577_),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _1185_ (.A(_0577_),
    .Y(_0048_));
 sky130_fd_sc_hd__inv_2 _1186_ (.A(_0577_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _1187_ (.A(_0577_),
    .Y(_0050_));
 sky130_fd_sc_hd__inv_2 _1188_ (.A(_0577_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _1189_ (.A(_0577_),
    .Y(_0052_));
 sky130_fd_sc_hd__inv_2 _1190_ (.A(_0577_),
    .Y(_0053_));
 sky130_fd_sc_hd__inv_2 _1191_ (.A(_0577_),
    .Y(_0054_));
 sky130_fd_sc_hd__inv_2 _1192_ (.A(_0577_),
    .Y(_0055_));
 sky130_fd_sc_hd__inv_2 _1193_ (.A(_0577_),
    .Y(_0056_));
 sky130_fd_sc_hd__inv_2 _1194_ (.A(_0574_),
    .Y(_0057_));
 sky130_fd_sc_hd__inv_2 _1195_ (.A(_0574_),
    .Y(_0058_));
 sky130_fd_sc_hd__inv_2 _1196_ (.A(_0574_),
    .Y(_0059_));
 sky130_fd_sc_hd__inv_2 _1197_ (.A(_0574_),
    .Y(_0060_));
 sky130_fd_sc_hd__inv_2 _1198_ (.A(_0574_),
    .Y(_0061_));
 sky130_fd_sc_hd__inv_2 _1199_ (.A(_0574_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _1200_ (.A(_0574_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _1201_ (.A(_0574_),
    .Y(_0064_));
 sky130_fd_sc_hd__inv_2 _1202_ (.A(_0574_),
    .Y(_0065_));
 sky130_fd_sc_hd__inv_2 _1203_ (.A(_0574_),
    .Y(_0066_));
 sky130_fd_sc_hd__inv_2 _1204_ (.A(_0574_),
    .Y(_0067_));
 sky130_fd_sc_hd__inv_2 _1205_ (.A(_0574_),
    .Y(_0068_));
 sky130_fd_sc_hd__dfrtp_2 _1206_ (.CLK(net17),
    .D(\M0.FCM2.q ),
    .RESET_B(_0000_),
    .Q(\M0.FCM4.q ));
 sky130_fd_sc_hd__dfrtp_2 _1207_ (.CLK(net17),
    .D(\M0.FCM1.q ),
    .RESET_B(_0001_),
    .Q(\M0.FCM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1208_ (.CLK(net17),
    .D(\M0.FPM15.d ),
    .RESET_B(_0002_),
    .Q(\M0.FPM15.q ));
 sky130_fd_sc_hd__dfrtp_1 _1209_ (.CLK(net17),
    .D(\M0.FPM14.d ),
    .RESET_B(_0003_),
    .Q(\M0.FPM14.q ));
 sky130_fd_sc_hd__dfrtp_1 _1210_ (.CLK(net17),
    .D(\M0.FPM13.d ),
    .RESET_B(_0004_),
    .Q(\M0.FPM13.q ));
 sky130_fd_sc_hd__dfrtp_1 _1211_ (.CLK(net17),
    .D(\M0.FPM12.d ),
    .RESET_B(_0005_),
    .Q(\M0.FPM12.q ));
 sky130_fd_sc_hd__dfrtp_1 _1212_ (.CLK(net17),
    .D(\M0.FPM11.d ),
    .RESET_B(_0006_),
    .Q(\M0.FPM11.q ));
 sky130_fd_sc_hd__dfrtp_1 _1213_ (.CLK(net17),
    .D(\M0.FPM10.d ),
    .RESET_B(_0007_),
    .Q(\M0.FPM10.q ));
 sky130_fd_sc_hd__dfrtp_1 _1214_ (.CLK(net17),
    .D(\M0.FPM9.d ),
    .RESET_B(_0008_),
    .Q(\M0.FPM9.q ));
 sky130_fd_sc_hd__dfrtp_1 _1215_ (.CLK(net17),
    .D(\M0.FPM8.d ),
    .RESET_B(_0009_),
    .Q(\M0.FPM8.q ));
 sky130_fd_sc_hd__dfrtp_1 _1216_ (.CLK(net17),
    .D(\M0.FPM7.d ),
    .RESET_B(_0010_),
    .Q(\M0.FPM7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1217_ (.CLK(net17),
    .D(\M0.FPM6.d ),
    .RESET_B(_0011_),
    .Q(\M0.FPM6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1218_ (.CLK(net17),
    .D(\M0.FPM5.d ),
    .RESET_B(_0012_),
    .Q(\M0.FPM5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1219_ (.CLK(net17),
    .D(\M0.FPM4.d ),
    .RESET_B(_0013_),
    .Q(\M0.FPM4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1220_ (.CLK(net17),
    .D(\M0.FPM3.d ),
    .RESET_B(_0014_),
    .Q(\M0.FPM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1221_ (.CLK(net17),
    .D(\M0.FPM2.d ),
    .RESET_B(_0015_),
    .Q(\M0.FPM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1222_ (.CLK(net17),
    .D(\M0.FPM1.d ),
    .RESET_B(_0016_),
    .Q(\M0.FPM1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1223_ (.CLK(net17),
    .D(\M0.FPM0.d ),
    .RESET_B(_0017_),
    .Q(\M0.FPM0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1224_ (.CLK(net17),
    .D(\M0.FCM2.d ),
    .RESET_B(_0018_),
    .Q(\M0.FCM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1225_ (.CLK(net17),
    .D(\M0.FCM1.d ),
    .RESET_B(_0019_),
    .Q(\M0.FCM1.q ));
 sky130_fd_sc_hd__dfrtp_4 _1226_ (.CLK(net17),
    .D(\M0.FBM7.d ),
    .RESET_B(_0020_),
    .Q(\M0.FBM7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1227_ (.CLK(net17),
    .D(\M0.FBM6.d ),
    .RESET_B(_0021_),
    .Q(\M0.FBM6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1228_ (.CLK(net17),
    .D(\M0.FBM5.d ),
    .RESET_B(_0022_),
    .Q(\M0.FBM5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1229_ (.CLK(net17),
    .D(\M0.FBM4.d ),
    .RESET_B(_0023_),
    .Q(\M0.FBM4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1230_ (.CLK(net17),
    .D(\M0.FBM3.d ),
    .RESET_B(_0024_),
    .Q(\M0.FBM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1231_ (.CLK(net17),
    .D(\M0.FBM2.d ),
    .RESET_B(_0025_),
    .Q(\M0.FBM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1232_ (.CLK(net17),
    .D(\M0.FBM1.d ),
    .RESET_B(_0026_),
    .Q(\M0.FBM1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1233_ (.CLK(net17),
    .D(\M0.FBM0.d ),
    .RESET_B(_0027_),
    .Q(\M0.FBM0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1234_ (.CLK(net17),
    .D(\M0.FAM7.d ),
    .RESET_B(_0028_),
    .Q(\M0.FAM7.q ));
 sky130_fd_sc_hd__dfrtp_1 _1235_ (.CLK(net17),
    .D(\M0.FAM6.d ),
    .RESET_B(_0029_),
    .Q(\M0.FAM6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1236_ (.CLK(net17),
    .D(\M0.FAM5.d ),
    .RESET_B(_0030_),
    .Q(\M0.FAM5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1237_ (.CLK(net17),
    .D(\M0.FAM4.d ),
    .RESET_B(_0031_),
    .Q(\M0.FAM4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1238_ (.CLK(net17),
    .D(\M0.FAM3.d ),
    .RESET_B(_0032_),
    .Q(\M0.FAM3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1239_ (.CLK(net17),
    .D(\M0.FAM2.d ),
    .RESET_B(_0033_),
    .Q(\M0.FAM2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1240_ (.CLK(net17),
    .D(\M0.FAM1.d ),
    .RESET_B(_0034_),
    .Q(\M0.FAM1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1241_ (.CLK(net17),
    .D(\M0.FAM0.d ),
    .RESET_B(_0035_),
    .Q(\M0.FAM0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1242_ (.CLK(net17),
    .D(\FP0.d ),
    .RESET_B(_0036_),
    .Q(net20));
 sky130_fd_sc_hd__dfrtp_1 _1243_ (.CLK(net17),
    .D(\FP1.d ),
    .RESET_B(_0037_),
    .Q(net27));
 sky130_fd_sc_hd__dfrtp_1 _1244_ (.CLK(net17),
    .D(\FP2.d ),
    .RESET_B(_0038_),
    .Q(net28));
 sky130_fd_sc_hd__dfrtp_1 _1245_ (.CLK(net17),
    .D(\FP3.d ),
    .RESET_B(_0039_),
    .Q(net29));
 sky130_fd_sc_hd__dfrtp_1 _1246_ (.CLK(net17),
    .D(\FP4.d ),
    .RESET_B(_0040_),
    .Q(net30));
 sky130_fd_sc_hd__dfrtp_1 _1247_ (.CLK(net17),
    .D(\FP5.d ),
    .RESET_B(_0041_),
    .Q(net31));
 sky130_fd_sc_hd__dfrtp_1 _1248_ (.CLK(net17),
    .D(\FP6.d ),
    .RESET_B(_0042_),
    .Q(net32));
 sky130_fd_sc_hd__dfrtp_1 _1249_ (.CLK(net17),
    .D(\FP7.d ),
    .RESET_B(_0043_),
    .Q(net33));
 sky130_fd_sc_hd__dfrtp_1 _1250_ (.CLK(net17),
    .D(\FP8.d ),
    .RESET_B(_0044_),
    .Q(net34));
 sky130_fd_sc_hd__dfrtp_1 _1251_ (.CLK(net17),
    .D(\FP9.d ),
    .RESET_B(_0045_),
    .Q(net35));
 sky130_fd_sc_hd__dfrtp_1 _1252_ (.CLK(net17),
    .D(\FP10.d ),
    .RESET_B(_0046_),
    .Q(net21));
 sky130_fd_sc_hd__dfrtp_1 _1253_ (.CLK(net17),
    .D(\FP11.d ),
    .RESET_B(_0047_),
    .Q(net22));
 sky130_fd_sc_hd__dfrtp_1 _1254_ (.CLK(net17),
    .D(\FP12.d ),
    .RESET_B(_0048_),
    .Q(net23));
 sky130_fd_sc_hd__dfrtp_1 _1255_ (.CLK(net17),
    .D(\FP13.d ),
    .RESET_B(_0049_),
    .Q(net24));
 sky130_fd_sc_hd__dfrtp_1 _1256_ (.CLK(net17),
    .D(\FP14.d ),
    .RESET_B(_0050_),
    .Q(net25));
 sky130_fd_sc_hd__dfrtp_1 _1257_ (.CLK(net17),
    .D(\FP15.d ),
    .RESET_B(_0051_),
    .Q(net26));
 sky130_fd_sc_hd__dfrtp_1 _1258_ (.CLK(net17),
    .D(net1),
    .RESET_B(_0052_),
    .Q(\FA0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1259_ (.CLK(net17),
    .D(net2),
    .RESET_B(_0053_),
    .Q(\FA1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1260_ (.CLK(net17),
    .D(net3),
    .RESET_B(_0054_),
    .Q(\FA2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1261_ (.CLK(net17),
    .D(net4),
    .RESET_B(_0055_),
    .Q(\FA3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1262_ (.CLK(net17),
    .D(net5),
    .RESET_B(_0056_),
    .Q(\FA4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1263_ (.CLK(net17),
    .D(net6),
    .RESET_B(_0057_),
    .Q(\FA5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1264_ (.CLK(net17),
    .D(net7),
    .RESET_B(_0058_),
    .Q(\FA6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1265_ (.CLK(net17),
    .D(net8),
    .RESET_B(_0059_),
    .Q(\FA7.q ));
 sky130_fd_sc_hd__dfrtp_2 _1266_ (.CLK(net17),
    .D(net9),
    .RESET_B(_0060_),
    .Q(\FB0.q ));
 sky130_fd_sc_hd__dfrtp_1 _1267_ (.CLK(net17),
    .D(net10),
    .RESET_B(_0061_),
    .Q(\FB1.q ));
 sky130_fd_sc_hd__dfrtp_1 _1268_ (.CLK(net17),
    .D(net11),
    .RESET_B(_0062_),
    .Q(\FB2.q ));
 sky130_fd_sc_hd__dfrtp_1 _1269_ (.CLK(net17),
    .D(net12),
    .RESET_B(_0063_),
    .Q(\FB3.q ));
 sky130_fd_sc_hd__dfrtp_1 _1270_ (.CLK(net17),
    .D(net13),
    .RESET_B(_0064_),
    .Q(\FB4.q ));
 sky130_fd_sc_hd__dfrtp_1 _1271_ (.CLK(net17),
    .D(net14),
    .RESET_B(_0065_),
    .Q(\FB5.q ));
 sky130_fd_sc_hd__dfrtp_1 _1272_ (.CLK(net17),
    .D(net15),
    .RESET_B(_0066_),
    .Q(\FB6.q ));
 sky130_fd_sc_hd__dfrtp_1 _1273_ (.CLK(net17),
    .D(net16),
    .RESET_B(_0067_),
    .Q(\FB7.q ));
 sky130_fd_sc_hd__dfrtp_2 _1274_ (.CLK(net17),
    .D(net18),
    .RESET_B(_0068_),
    .Q(\FC.q ));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(a[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(b[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(b[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(b[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(b[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(b[5]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(b[6]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(b[7]),
    .X(net16));
 sky130_fd_sc_hd__buf_12 input17 (.A(clk),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(control),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(rst),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(a[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(a[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(a[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(a[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(a[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(a[6]),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(a[7]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(b[0]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 max_cap48 (.A(net58),
    .X(net48));
 sky130_fd_sc_hd__buf_2 max_cap49 (.A(_0100_),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 max_cap8 (.A(net58),
    .X(net57));
 sky130_fd_sc_hd__buf_12 output20 (.A(net20),
    .X(p[0]));
 sky130_fd_sc_hd__buf_12 output21 (.A(net21),
    .X(p[10]));
 sky130_fd_sc_hd__buf_12 output22 (.A(net22),
    .X(p[11]));
 sky130_fd_sc_hd__buf_12 output23 (.A(net23),
    .X(p[12]));
 sky130_fd_sc_hd__buf_12 output24 (.A(net24),
    .X(p[13]));
 sky130_fd_sc_hd__buf_12 output25 (.A(net25),
    .X(p[14]));
 sky130_fd_sc_hd__buf_12 output26 (.A(net26),
    .X(p[15]));
 sky130_fd_sc_hd__buf_12 output27 (.A(net27),
    .X(p[1]));
 sky130_fd_sc_hd__buf_12 output28 (.A(net28),
    .X(p[2]));
 sky130_fd_sc_hd__buf_12 output29 (.A(net29),
    .X(p[3]));
 sky130_fd_sc_hd__buf_12 output30 (.A(net30),
    .X(p[4]));
 sky130_fd_sc_hd__buf_12 output31 (.A(net31),
    .X(p[5]));
 sky130_fd_sc_hd__buf_12 output32 (.A(net32),
    .X(p[6]));
 sky130_fd_sc_hd__buf_12 output33 (.A(net33),
    .X(p[7]));
 sky130_fd_sc_hd__buf_12 output34 (.A(net34),
    .X(p[8]));
 sky130_fd_sc_hd__buf_12 output35 (.A(net35),
    .X(p[9]));
 sky130_fd_sc_hd__clkbuf_1 wire1 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 wire2 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 wire3 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 wire36 (.A(net37),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 wire37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 wire38 (.A(net39),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 wire39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 wire4 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 wire40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 wire41 (.A(net42),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 wire42 (.A(net43),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 wire43 (.A(net44),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 wire44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 wire45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 wire46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 wire47 (.A(net50),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 wire5 (.A(net55),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 wire6 (.A(net56),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 wire7 (.A(_0254_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 wire9 (.A(_0220_),
    .X(net58));
endmodule

